magic
tech sky130B
magscale 1 2
timestamp 1661721387
<< obsli1 >>
rect 0 0 584000 704000
<< metal1 >>
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 206278 702448 206284 702500
rect 206336 702488 206342 702500
rect 559650 702488 559656 702500
rect 206336 702460 559656 702488
rect 206336 702448 206342 702460
rect 559650 702448 559656 702460
rect 559708 702448 559714 702500
rect 300118 700408 300124 700460
rect 300176 700448 300182 700460
rect 310514 700448 310520 700460
rect 300176 700420 310520 700448
rect 300176 700408 300182 700420
rect 310514 700408 310520 700420
rect 310572 700408 310578 700460
rect 149698 700340 149704 700392
rect 149756 700380 149762 700392
rect 170306 700380 170312 700392
rect 149756 700352 170312 700380
rect 149756 700340 149762 700352
rect 170306 700340 170312 700352
rect 170364 700340 170370 700392
rect 218974 700340 218980 700392
rect 219032 700380 219038 700392
rect 309134 700380 309140 700392
rect 219032 700352 309140 700380
rect 219032 700340 219038 700352
rect 309134 700340 309140 700352
rect 309192 700340 309198 700392
rect 354582 700340 354588 700392
rect 354640 700380 354646 700392
rect 364978 700380 364984 700392
rect 354640 700352 364984 700380
rect 354640 700340 354646 700352
rect 364978 700340 364984 700352
rect 365036 700340 365042 700392
rect 383562 700340 383568 700392
rect 383620 700380 383626 700392
rect 478506 700380 478512 700392
rect 383620 700352 478512 700380
rect 383620 700340 383626 700352
rect 478506 700340 478512 700352
rect 478564 700340 478570 700392
rect 559650 700340 559656 700392
rect 559708 700380 559714 700392
rect 582374 700380 582380 700392
rect 559708 700352 582380 700380
rect 559708 700340 559714 700352
rect 582374 700340 582380 700352
rect 582432 700340 582438 700392
rect 72970 700272 72976 700324
rect 73028 700312 73034 700324
rect 94498 700312 94504 700324
rect 73028 700284 94504 700312
rect 73028 700272 73034 700284
rect 94498 700272 94504 700284
rect 94556 700272 94562 700324
rect 105446 700272 105452 700324
rect 105504 700312 105510 700324
rect 193214 700312 193220 700324
rect 105504 700284 193220 700312
rect 105504 700272 105510 700284
rect 193214 700272 193220 700284
rect 193272 700272 193278 700324
rect 235166 700272 235172 700324
rect 235224 700312 235230 700324
rect 299474 700312 299480 700324
rect 235224 700284 299480 700312
rect 235224 700272 235230 700284
rect 299474 700272 299480 700284
rect 299532 700272 299538 700324
rect 302050 700272 302056 700324
rect 302108 700312 302114 700324
rect 429838 700312 429844 700324
rect 302108 700284 429844 700312
rect 302108 700272 302114 700284
rect 429838 700272 429844 700284
rect 429896 700272 429902 700324
rect 527174 700272 527180 700324
rect 527232 700312 527238 700324
rect 565814 700312 565820 700324
rect 527232 700284 565820 700312
rect 527232 700272 527238 700284
rect 565814 700272 565820 700284
rect 565872 700272 565878 700324
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 25498 699700 25504 699712
rect 24360 699672 25504 699700
rect 24360 699660 24366 699672
rect 25498 699660 25504 699672
rect 25556 699660 25562 699712
rect 307662 698912 307668 698964
rect 307720 698952 307726 698964
rect 397454 698952 397460 698964
rect 307720 698924 397460 698952
rect 307720 698912 307726 698924
rect 397454 698912 397460 698924
rect 397512 698912 397518 698964
rect 179046 697552 179052 697604
rect 179104 697592 179110 697604
rect 267642 697592 267648 697604
rect 179104 697564 267648 697592
rect 179104 697552 179110 697564
rect 267642 697552 267648 697564
rect 267700 697552 267706 697604
rect 212442 696192 212448 696244
rect 212500 696232 212506 696244
rect 348786 696232 348792 696244
rect 212500 696204 348792 696232
rect 212500 696192 212506 696204
rect 348786 696192 348792 696204
rect 348844 696192 348850 696244
rect 3418 684156 3424 684208
rect 3476 684196 3482 684208
rect 8938 684196 8944 684208
rect 3476 684168 8944 684196
rect 3476 684156 3482 684168
rect 8938 684156 8944 684168
rect 8996 684156 9002 684208
rect 567838 683136 567844 683188
rect 567896 683176 567902 683188
rect 580166 683176 580172 683188
rect 567896 683148 580172 683176
rect 567896 683136 567902 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 66898 670732 66904 670744
rect 3568 670704 66904 670732
rect 3568 670692 3574 670704
rect 66898 670692 66904 670704
rect 66956 670692 66962 670744
rect 6914 669944 6920 669996
rect 6972 669984 6978 669996
rect 62758 669984 62764 669996
rect 6972 669956 62764 669984
rect 6972 669944 6978 669956
rect 62758 669944 62764 669956
rect 62816 669944 62822 669996
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 32398 656928 32404 656940
rect 3476 656900 32404 656928
rect 3476 656888 3482 656900
rect 32398 656888 32404 656900
rect 32456 656888 32462 656940
rect 574738 643084 574744 643136
rect 574796 643124 574802 643136
rect 580166 643124 580172 643136
rect 574796 643096 580172 643124
rect 574796 643084 574802 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 44818 632108 44824 632120
rect 3476 632080 44824 632108
rect 3476 632068 3482 632080
rect 44818 632068 44824 632080
rect 44876 632068 44882 632120
rect 502978 630640 502984 630692
rect 503036 630680 503042 630692
rect 580166 630680 580172 630692
rect 503036 630652 580172 630680
rect 503036 630640 503042 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 22738 618304 22744 618316
rect 3200 618276 22744 618304
rect 3200 618264 3206 618276
rect 22738 618264 22744 618276
rect 22796 618264 22802 618316
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 90358 605860 90364 605872
rect 3292 605832 90364 605860
rect 3292 605820 3298 605832
rect 90358 605820 90364 605832
rect 90416 605820 90422 605872
rect 530578 590656 530584 590708
rect 530636 590696 530642 590708
rect 579798 590696 579804 590708
rect 530636 590668 579804 590696
rect 530636 590656 530642 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 391198 576852 391204 576904
rect 391256 576892 391262 576904
rect 580166 576892 580172 576904
rect 391256 576864 580172 576892
rect 391256 576852 391262 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 57238 565876 57244 565888
rect 3476 565848 57244 565876
rect 3476 565836 3482 565848
rect 57238 565836 57244 565848
rect 57296 565836 57302 565888
rect 3418 553392 3424 553444
rect 3476 553432 3482 553444
rect 36538 553432 36544 553444
rect 3476 553404 36544 553432
rect 3476 553392 3482 553404
rect 36538 553392 36544 553404
rect 36596 553392 36602 553444
rect 576118 536800 576124 536852
rect 576176 536840 576182 536852
rect 580166 536840 580172 536852
rect 576176 536812 580172 536840
rect 576176 536800 576182 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 3418 527144 3424 527196
rect 3476 527184 3482 527196
rect 39298 527184 39304 527196
rect 3476 527156 39304 527184
rect 3476 527144 3482 527156
rect 39298 527144 39304 527156
rect 39356 527144 39362 527196
rect 3418 514768 3424 514820
rect 3476 514808 3482 514820
rect 48958 514808 48964 514820
rect 3476 514780 48964 514808
rect 3476 514768 3482 514780
rect 48958 514768 48964 514780
rect 49016 514768 49022 514820
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 120718 501004 120724 501016
rect 3108 500976 120724 501004
rect 3108 500964 3114 500976
rect 120718 500964 120724 500976
rect 120776 500964 120782 501016
rect 536098 484372 536104 484424
rect 536156 484412 536162 484424
rect 580166 484412 580172 484424
rect 536156 484384 580172 484412
rect 536156 484372 536162 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 3418 474716 3424 474768
rect 3476 474756 3482 474768
rect 31018 474756 31024 474768
rect 3476 474728 31024 474756
rect 3476 474716 3482 474728
rect 31018 474716 31024 474728
rect 31076 474716 31082 474768
rect 274542 470568 274548 470620
rect 274600 470608 274606 470620
rect 580166 470608 580172 470620
rect 274600 470580 580172 470608
rect 274600 470568 274606 470580
rect 580166 470568 580172 470580
rect 580224 470568 580230 470620
rect 3234 462340 3240 462392
rect 3292 462380 3298 462392
rect 98638 462380 98644 462392
rect 3292 462352 98644 462380
rect 3292 462340 3298 462352
rect 98638 462340 98644 462352
rect 98696 462340 98702 462392
rect 573358 458804 573364 458856
rect 573416 458844 573422 458856
rect 580258 458844 580264 458856
rect 573416 458816 580264 458844
rect 573416 458804 573422 458816
rect 580258 458804 580264 458816
rect 580316 458804 580322 458856
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 53098 448576 53104 448588
rect 3200 448548 53104 448576
rect 3200 448536 3206 448548
rect 53098 448536 53104 448548
rect 53156 448536 53162 448588
rect 392578 430584 392584 430636
rect 392636 430624 392642 430636
rect 580166 430624 580172 430636
rect 392636 430596 580172 430624
rect 392636 430584 392642 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 3418 422288 3424 422340
rect 3476 422328 3482 422340
rect 13078 422328 13084 422340
rect 3476 422300 13084 422328
rect 3476 422288 3482 422300
rect 13078 422288 13084 422300
rect 13136 422288 13142 422340
rect 577498 418140 577504 418192
rect 577556 418180 577562 418192
rect 579614 418180 579620 418192
rect 577556 418152 579620 418180
rect 577556 418140 577562 418152
rect 579614 418140 579620 418152
rect 579672 418140 579678 418192
rect 3142 409844 3148 409896
rect 3200 409884 3206 409896
rect 50338 409884 50344 409896
rect 3200 409856 50344 409884
rect 3200 409844 3206 409856
rect 50338 409844 50344 409856
rect 50396 409844 50402 409896
rect 388438 404336 388444 404388
rect 388496 404376 388502 404388
rect 580166 404376 580172 404388
rect 388496 404348 580172 404376
rect 388496 404336 388502 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3418 397468 3424 397520
rect 3476 397508 3482 397520
rect 58618 397508 58624 397520
rect 3476 397480 58624 397508
rect 3476 397468 3482 397480
rect 58618 397468 58624 397480
rect 58676 397468 58682 397520
rect 48958 381488 48964 381540
rect 49016 381528 49022 381540
rect 247034 381528 247040 381540
rect 49016 381500 247040 381528
rect 49016 381488 49022 381500
rect 247034 381488 247040 381500
rect 247092 381488 247098 381540
rect 153194 380128 153200 380180
rect 153252 380168 153258 380180
rect 270494 380168 270500 380180
rect 153252 380140 270500 380168
rect 153252 380128 153258 380140
rect 270494 380128 270500 380140
rect 270552 380128 270558 380180
rect 55030 378768 55036 378820
rect 55088 378808 55094 378820
rect 138014 378808 138020 378820
rect 55088 378780 138020 378808
rect 55088 378768 55094 378780
rect 138014 378768 138020 378780
rect 138072 378808 138078 378820
rect 295334 378808 295340 378820
rect 138072 378780 295340 378808
rect 138072 378768 138078 378780
rect 295334 378768 295340 378780
rect 295392 378768 295398 378820
rect 574094 377408 574100 377460
rect 574152 377448 574158 377460
rect 580166 377448 580172 377460
rect 574152 377420 580172 377448
rect 574152 377408 574158 377420
rect 580166 377408 580172 377420
rect 580224 377408 580230 377460
rect 209038 376728 209044 376780
rect 209096 376768 209102 376780
rect 574094 376768 574100 376780
rect 209096 376740 574100 376768
rect 209096 376728 209102 376740
rect 574094 376728 574100 376740
rect 574152 376728 574158 376780
rect 195238 374620 195244 374672
rect 195296 374660 195302 374672
rect 331214 374660 331220 374672
rect 195296 374632 331220 374660
rect 195296 374620 195302 374632
rect 331214 374620 331220 374632
rect 331272 374620 331278 374672
rect 53098 372580 53104 372632
rect 53156 372620 53162 372632
rect 53742 372620 53748 372632
rect 53156 372592 53748 372620
rect 53156 372580 53162 372592
rect 53742 372580 53748 372592
rect 53800 372620 53806 372632
rect 291838 372620 291844 372632
rect 53800 372592 291844 372620
rect 53800 372580 53806 372592
rect 291838 372580 291844 372592
rect 291896 372580 291902 372632
rect 98638 371832 98644 371884
rect 98696 371872 98702 371884
rect 125594 371872 125600 371884
rect 98696 371844 125600 371872
rect 98696 371832 98702 371844
rect 125594 371832 125600 371844
rect 125652 371872 125658 371884
rect 126606 371872 126612 371884
rect 125652 371844 126612 371872
rect 125652 371832 125658 371844
rect 126606 371832 126612 371844
rect 126664 371832 126670 371884
rect 232498 371288 232504 371340
rect 232556 371328 232562 371340
rect 313918 371328 313924 371340
rect 232556 371300 313924 371328
rect 232556 371288 232562 371300
rect 313918 371288 313924 371300
rect 313976 371288 313982 371340
rect 3418 371220 3424 371272
rect 3476 371260 3482 371272
rect 111058 371260 111064 371272
rect 3476 371232 111064 371260
rect 3476 371220 3482 371232
rect 111058 371220 111064 371232
rect 111116 371220 111122 371272
rect 126606 371220 126612 371272
rect 126664 371260 126670 371272
rect 266998 371260 267004 371272
rect 126664 371232 267004 371260
rect 126664 371220 126670 371232
rect 266998 371220 267004 371232
rect 267056 371220 267062 371272
rect 8938 370472 8944 370524
rect 8996 370512 9002 370524
rect 144086 370512 144092 370524
rect 8996 370484 144092 370512
rect 8996 370472 9002 370484
rect 144086 370472 144092 370484
rect 144144 370472 144150 370524
rect 143534 369860 143540 369912
rect 143592 369900 143598 369912
rect 144086 369900 144092 369912
rect 143592 369872 144092 369900
rect 143592 369860 143598 369872
rect 144086 369860 144092 369872
rect 144144 369900 144150 369912
rect 198734 369900 198740 369912
rect 144144 369872 198740 369900
rect 144144 369860 144150 369872
rect 198734 369860 198740 369872
rect 198792 369860 198798 369912
rect 211798 369860 211804 369912
rect 211856 369900 211862 369912
rect 212442 369900 212448 369912
rect 211856 369872 212448 369900
rect 211856 369860 211862 369872
rect 212442 369860 212448 369872
rect 212500 369900 212506 369912
rect 583018 369900 583024 369912
rect 212500 369872 583024 369900
rect 212500 369860 212506 369872
rect 583018 369860 583024 369872
rect 583076 369860 583082 369912
rect 31018 369112 31024 369164
rect 31076 369152 31082 369164
rect 146938 369152 146944 369164
rect 31076 369124 146944 369152
rect 31076 369112 31082 369124
rect 146938 369112 146944 369124
rect 146996 369112 147002 369164
rect 146938 368636 146944 368688
rect 146996 368676 147002 368688
rect 202874 368676 202880 368688
rect 146996 368648 202880 368676
rect 146996 368636 147002 368648
rect 202874 368636 202880 368648
rect 202932 368636 202938 368688
rect 140038 368568 140044 368620
rect 140096 368608 140102 368620
rect 282914 368608 282920 368620
rect 140096 368580 282920 368608
rect 140096 368568 140102 368580
rect 282914 368568 282920 368580
rect 282972 368568 282978 368620
rect 170950 368500 170956 368552
rect 171008 368540 171014 368552
rect 578234 368540 578240 368552
rect 171008 368512 578240 368540
rect 171008 368500 171014 368512
rect 578234 368500 578240 368512
rect 578292 368540 578298 368552
rect 578878 368540 578884 368552
rect 578292 368512 578884 368540
rect 578292 368500 578298 368512
rect 578878 368500 578884 368512
rect 578936 368500 578942 368552
rect 39298 368432 39304 368484
rect 39356 368472 39362 368484
rect 39942 368472 39948 368484
rect 39356 368444 39948 368472
rect 39356 368432 39362 368444
rect 39942 368432 39948 368444
rect 40000 368432 40006 368484
rect 282914 367752 282920 367804
rect 282972 367792 282978 367804
rect 293954 367792 293960 367804
rect 282972 367764 293960 367792
rect 282972 367752 282978 367764
rect 293954 367752 293960 367764
rect 294012 367752 294018 367804
rect 226334 367276 226340 367328
rect 226392 367316 226398 367328
rect 340874 367316 340880 367328
rect 226392 367288 340880 367316
rect 226392 367276 226398 367288
rect 340874 367276 340880 367288
rect 340932 367276 340938 367328
rect 114554 367208 114560 367260
rect 114612 367248 114618 367260
rect 295978 367248 295984 367260
rect 114612 367220 295984 367248
rect 114612 367208 114618 367220
rect 295978 367208 295984 367220
rect 296036 367208 296042 367260
rect 39942 367140 39948 367192
rect 40000 367180 40006 367192
rect 264238 367180 264244 367192
rect 40000 367152 264244 367180
rect 40000 367140 40006 367152
rect 264238 367140 264244 367152
rect 264296 367140 264302 367192
rect 175090 367072 175096 367124
rect 175148 367112 175154 367124
rect 561950 367112 561956 367124
rect 175148 367084 561956 367112
rect 175148 367072 175154 367084
rect 561950 367072 561956 367084
rect 562008 367072 562014 367124
rect 171778 366392 171784 366444
rect 171836 366432 171842 366444
rect 201494 366432 201500 366444
rect 171836 366404 201500 366432
rect 171836 366392 171842 366404
rect 201494 366392 201500 366404
rect 201552 366392 201558 366444
rect 32398 366324 32404 366376
rect 32456 366364 32462 366376
rect 234614 366364 234620 366376
rect 32456 366336 234620 366364
rect 32456 366324 32462 366336
rect 234614 366324 234620 366336
rect 234672 366324 234678 366376
rect 189074 365780 189080 365832
rect 189132 365820 189138 365832
rect 307018 365820 307024 365832
rect 189132 365792 307024 365820
rect 189132 365780 189138 365792
rect 307018 365780 307024 365792
rect 307076 365780 307082 365832
rect 219434 365712 219440 365764
rect 219492 365752 219498 365764
rect 571426 365752 571432 365764
rect 219492 365724 571432 365752
rect 219492 365712 219498 365724
rect 571426 365712 571432 365724
rect 571484 365712 571490 365764
rect 208394 365644 208400 365696
rect 208452 365684 208458 365696
rect 209038 365684 209044 365696
rect 208452 365656 209044 365684
rect 208452 365644 208458 365656
rect 209038 365644 209044 365656
rect 209096 365644 209102 365696
rect 238754 364556 238760 364608
rect 238812 364596 238818 364608
rect 302234 364596 302240 364608
rect 238812 364568 302240 364596
rect 238812 364556 238818 364568
rect 302234 364556 302240 364568
rect 302292 364556 302298 364608
rect 162302 364488 162308 364540
rect 162360 364528 162366 364540
rect 208394 364528 208400 364540
rect 162360 364500 208400 364528
rect 162360 364488 162366 364500
rect 208394 364488 208400 364500
rect 208452 364488 208458 364540
rect 251174 364488 251180 364540
rect 251232 364528 251238 364540
rect 331214 364528 331220 364540
rect 251232 364500 331220 364528
rect 251232 364488 251238 364500
rect 331214 364488 331220 364500
rect 331272 364488 331278 364540
rect 128998 364420 129004 364472
rect 129056 364460 129062 364472
rect 282914 364460 282920 364472
rect 129056 364432 282920 364460
rect 129056 364420 129062 364432
rect 282914 364420 282920 364432
rect 282972 364420 282978 364472
rect 120718 364352 120724 364404
rect 120776 364392 120782 364404
rect 296898 364392 296904 364404
rect 120776 364364 296904 364392
rect 120776 364352 120782 364364
rect 296898 364352 296904 364364
rect 296956 364352 296962 364404
rect 570506 364352 570512 364404
rect 570564 364392 570570 364404
rect 580166 364392 580172 364404
rect 570564 364364 580172 364392
rect 570564 364352 570570 364364
rect 580166 364352 580172 364364
rect 580224 364352 580230 364404
rect 228818 363128 228824 363180
rect 228876 363168 228882 363180
rect 318058 363168 318064 363180
rect 228876 363140 318064 363168
rect 228876 363128 228882 363140
rect 318058 363128 318064 363140
rect 318116 363128 318122 363180
rect 166258 363060 166264 363112
rect 166316 363100 166322 363112
rect 287422 363100 287428 363112
rect 166316 363072 287428 363100
rect 166316 363060 166322 363072
rect 287422 363060 287428 363072
rect 287480 363060 287486 363112
rect 130378 362992 130384 363044
rect 130436 363032 130442 363044
rect 298278 363032 298284 363044
rect 130436 363004 298284 363032
rect 130436 362992 130442 363004
rect 298278 362992 298284 363004
rect 298336 362992 298342 363044
rect 178678 362924 178684 362976
rect 178736 362964 178742 362976
rect 580350 362964 580356 362976
rect 178736 362936 580356 362964
rect 178736 362924 178742 362936
rect 580350 362924 580356 362936
rect 580408 362924 580414 362976
rect 138658 361904 138664 361956
rect 138716 361944 138722 361956
rect 193214 361944 193220 361956
rect 138716 361916 193220 361944
rect 138716 361904 138722 361916
rect 193214 361904 193220 361916
rect 193272 361904 193278 361956
rect 134518 361836 134524 361888
rect 134576 361876 134582 361888
rect 231670 361876 231676 361888
rect 134576 361848 231676 361876
rect 134576 361836 134582 361848
rect 231670 361836 231676 361848
rect 231728 361876 231734 361888
rect 315298 361876 315304 361888
rect 231728 361848 315304 361876
rect 231728 361836 231734 361848
rect 315298 361836 315304 361848
rect 315356 361836 315362 361888
rect 181622 361768 181628 361820
rect 181680 361808 181686 361820
rect 319438 361808 319444 361820
rect 181680 361780 319444 361808
rect 181680 361768 181686 361780
rect 319438 361768 319444 361780
rect 319496 361768 319502 361820
rect 111150 361700 111156 361752
rect 111208 361740 111214 361752
rect 299566 361740 299572 361752
rect 111208 361712 299572 361740
rect 111208 361700 111214 361712
rect 299566 361700 299572 361712
rect 299624 361700 299630 361752
rect 179506 361632 179512 361684
rect 179564 361672 179570 361684
rect 463418 361672 463424 361684
rect 179564 361644 463424 361672
rect 179564 361632 179570 361644
rect 463418 361632 463424 361644
rect 463476 361632 463482 361684
rect 64782 361564 64788 361616
rect 64840 361604 64846 361616
rect 195238 361604 195244 361616
rect 64840 361576 195244 361604
rect 64840 361564 64846 361576
rect 195238 361564 195244 361576
rect 195296 361564 195302 361616
rect 243630 361564 243636 361616
rect 243688 361604 243694 361616
rect 563698 361604 563704 361616
rect 243688 361576 563704 361604
rect 243688 361564 243694 361576
rect 563698 361564 563704 361576
rect 563756 361564 563762 361616
rect 126238 360612 126244 360664
rect 126296 360652 126302 360664
rect 279326 360652 279332 360664
rect 126296 360624 279332 360652
rect 126296 360612 126302 360624
rect 279326 360612 279332 360624
rect 279384 360652 279390 360664
rect 280062 360652 280068 360664
rect 279384 360624 280068 360652
rect 279384 360612 279390 360624
rect 280062 360612 280068 360624
rect 280120 360612 280126 360664
rect 250530 360544 250536 360596
rect 250588 360584 250594 360596
rect 297358 360584 297364 360596
rect 250588 360556 297364 360584
rect 250588 360544 250594 360556
rect 297358 360544 297364 360556
rect 297416 360544 297422 360596
rect 176102 360476 176108 360528
rect 176160 360516 176166 360528
rect 237466 360516 237472 360528
rect 176160 360488 237472 360516
rect 176160 360476 176166 360488
rect 237466 360476 237472 360488
rect 237524 360516 237530 360528
rect 329190 360516 329196 360528
rect 237524 360488 329196 360516
rect 237524 360476 237530 360488
rect 329190 360476 329196 360488
rect 329248 360476 329254 360528
rect 176010 360408 176016 360460
rect 176068 360448 176074 360460
rect 219434 360448 219440 360460
rect 176068 360420 219440 360448
rect 176068 360408 176074 360420
rect 219434 360408 219440 360420
rect 219492 360448 219498 360460
rect 220262 360448 220268 360460
rect 219492 360420 220268 360448
rect 219492 360408 219498 360420
rect 220262 360408 220268 360420
rect 220320 360408 220326 360460
rect 233786 360408 233792 360460
rect 233844 360448 233850 360460
rect 332594 360448 332600 360460
rect 233844 360420 332600 360448
rect 233844 360408 233850 360420
rect 332594 360408 332600 360420
rect 332652 360408 332658 360460
rect 113174 360340 113180 360392
rect 113232 360380 113238 360392
rect 296806 360380 296812 360392
rect 113232 360352 296812 360380
rect 113232 360340 113238 360352
rect 296806 360340 296812 360352
rect 296864 360340 296870 360392
rect 275002 360272 275008 360324
rect 275060 360312 275066 360324
rect 538858 360312 538864 360324
rect 275060 360284 538864 360312
rect 275060 360272 275066 360284
rect 538858 360272 538864 360284
rect 538916 360272 538922 360324
rect 79318 360204 79324 360256
rect 79376 360244 79382 360256
rect 245838 360244 245844 360256
rect 79376 360216 245844 360244
rect 79376 360204 79382 360216
rect 245838 360204 245844 360216
rect 245896 360204 245902 360256
rect 280062 360204 280068 360256
rect 280120 360244 280126 360256
rect 578326 360244 578332 360256
rect 280120 360216 578332 360244
rect 280120 360204 280126 360216
rect 578326 360204 578332 360216
rect 578384 360204 578390 360256
rect 172422 359116 172428 359168
rect 172480 359156 172486 359168
rect 218330 359156 218336 359168
rect 172480 359128 218336 359156
rect 172480 359116 172486 359128
rect 218330 359116 218336 359128
rect 218388 359116 218394 359168
rect 173158 359048 173164 359100
rect 173216 359088 173222 359100
rect 296714 359088 296720 359100
rect 173216 359060 296720 359088
rect 173216 359048 173222 359060
rect 296714 359048 296720 359060
rect 296772 359048 296778 359100
rect 142798 358980 142804 359032
rect 142856 359020 142862 359032
rect 201586 359020 201592 359032
rect 142856 358992 201592 359020
rect 142856 358980 142862 358992
rect 201586 358980 201592 358992
rect 201644 358980 201650 359032
rect 234614 358980 234620 359032
rect 234672 359020 234678 359032
rect 235534 359020 235540 359032
rect 234672 358992 235540 359020
rect 234672 358980 234678 358992
rect 235534 358980 235540 358992
rect 235592 359020 235598 359032
rect 374638 359020 374644 359032
rect 235592 358992 374644 359020
rect 235592 358980 235598 358992
rect 374638 358980 374644 358992
rect 374696 358980 374702 359032
rect 109034 358912 109040 358964
rect 109092 358952 109098 358964
rect 253934 358952 253940 358964
rect 109092 358924 253940 358952
rect 109092 358912 109098 358924
rect 253934 358912 253940 358924
rect 253992 358912 253998 358964
rect 264238 358912 264244 358964
rect 264296 358952 264302 358964
rect 264882 358952 264888 358964
rect 264296 358924 264888 358952
rect 264296 358912 264302 358924
rect 264882 358912 264888 358924
rect 264940 358952 264946 358964
rect 305638 358952 305644 358964
rect 264940 358924 305644 358952
rect 264940 358912 264946 358924
rect 305638 358912 305644 358924
rect 305696 358912 305702 358964
rect 101398 358844 101404 358896
rect 101456 358884 101462 358896
rect 293126 358884 293132 358896
rect 101456 358856 293132 358884
rect 101456 358844 101462 358856
rect 293126 358844 293132 358856
rect 293184 358844 293190 358896
rect 179230 358776 179236 358828
rect 179288 358816 179294 358828
rect 421558 358816 421564 358828
rect 179288 358788 421564 358816
rect 179288 358776 179294 358788
rect 421558 358776 421564 358788
rect 421616 358776 421622 358828
rect 213914 358708 213920 358760
rect 213972 358748 213978 358760
rect 214466 358748 214472 358760
rect 213972 358720 214472 358748
rect 213972 358708 213978 358720
rect 214466 358708 214472 358720
rect 214524 358708 214530 358760
rect 282914 358708 282920 358760
rect 282972 358748 282978 358760
rect 283558 358748 283564 358760
rect 282972 358720 283564 358748
rect 282972 358708 282978 358720
rect 283558 358708 283564 358720
rect 283616 358708 283622 358760
rect 217042 358096 217048 358148
rect 217100 358136 217106 358148
rect 232498 358136 232504 358148
rect 217100 358108 232504 358136
rect 217100 358096 217106 358108
rect 232498 358096 232504 358108
rect 232556 358096 232562 358148
rect 214558 358028 214564 358080
rect 214616 358068 214622 358080
rect 275002 358068 275008 358080
rect 214616 358040 275008 358068
rect 214616 358028 214622 358040
rect 275002 358028 275008 358040
rect 275060 358068 275066 358080
rect 276934 358068 276940 358080
rect 275060 358040 276940 358068
rect 275060 358028 275066 358040
rect 276934 358028 276940 358040
rect 276992 358028 276998 358080
rect 387702 358028 387708 358080
rect 387760 358068 387766 358080
rect 570506 358068 570512 358080
rect 387760 358040 570512 358068
rect 387760 358028 387766 358040
rect 570506 358028 570512 358040
rect 570564 358028 570570 358080
rect 158622 357756 158628 357808
rect 158680 357796 158686 357808
rect 182910 357796 182916 357808
rect 158680 357768 182916 357796
rect 158680 357756 158686 357768
rect 182910 357756 182916 357768
rect 182968 357756 182974 357808
rect 275646 357756 275652 357808
rect 275704 357796 275710 357808
rect 300854 357796 300860 357808
rect 275704 357768 300860 357796
rect 275704 357756 275710 357768
rect 300854 357756 300860 357768
rect 300912 357756 300918 357808
rect 164142 357688 164148 357740
rect 164200 357728 164206 357740
rect 186774 357728 186780 357740
rect 164200 357700 186780 357728
rect 164200 357688 164206 357700
rect 186774 357688 186780 357700
rect 186832 357688 186838 357740
rect 195238 357688 195244 357740
rect 195296 357728 195302 357740
rect 200022 357728 200028 357740
rect 195296 357700 200028 357728
rect 195296 357688 195302 357700
rect 200022 357688 200028 357700
rect 200080 357688 200086 357740
rect 266998 357688 267004 357740
rect 267056 357728 267062 357740
rect 293218 357728 293224 357740
rect 267056 357700 293224 357728
rect 267056 357688 267062 357700
rect 293218 357688 293224 357700
rect 293276 357688 293282 357740
rect 179874 357620 179880 357672
rect 179932 357660 179938 357672
rect 214466 357660 214472 357672
rect 179932 357632 214472 357660
rect 179932 357620 179938 357632
rect 214466 357620 214472 357632
rect 214524 357620 214530 357672
rect 223482 357620 223488 357672
rect 223540 357660 223546 357672
rect 298094 357660 298100 357672
rect 223540 357632 298100 357660
rect 223540 357620 223546 357632
rect 298094 357620 298100 357632
rect 298152 357620 298158 357672
rect 154482 357552 154488 357604
rect 154540 357592 154546 357604
rect 184934 357592 184940 357604
rect 154540 357564 184940 357592
rect 154540 357552 154546 357564
rect 184934 357552 184940 357564
rect 184992 357552 184998 357604
rect 191742 357552 191748 357604
rect 191800 357592 191806 357604
rect 285674 357592 285680 357604
rect 191800 357564 285680 357592
rect 191800 357552 191806 357564
rect 285674 357552 285680 357564
rect 285732 357552 285738 357604
rect 287422 357552 287428 357604
rect 287480 357592 287486 357604
rect 292206 357592 292212 357604
rect 287480 357564 292212 357592
rect 287480 357552 287486 357564
rect 292206 357552 292212 357564
rect 292264 357552 292270 357604
rect 292298 357552 292304 357604
rect 292356 357592 292362 357604
rect 363598 357592 363604 357604
rect 292356 357564 363604 357592
rect 292356 357552 292362 357564
rect 363598 357552 363604 357564
rect 363656 357552 363662 357604
rect 135898 357484 135904 357536
rect 135956 357524 135962 357536
rect 256786 357524 256792 357536
rect 135956 357496 256792 357524
rect 135956 357484 135962 357496
rect 256786 357484 256792 357496
rect 256844 357484 256850 357536
rect 283558 357484 283564 357536
rect 283616 357524 283622 357536
rect 435082 357524 435088 357536
rect 283616 357496 435088 357524
rect 283616 357484 283622 357496
rect 435082 357484 435088 357496
rect 435140 357484 435146 357536
rect 80054 357416 80060 357468
rect 80112 357456 80118 357468
rect 300946 357456 300952 357468
rect 80112 357428 300952 357456
rect 80112 357416 80118 357428
rect 300946 357416 300952 357428
rect 301004 357416 301010 357468
rect 200022 357348 200028 357400
rect 200080 357388 200086 357400
rect 201494 357388 201500 357400
rect 200080 357360 201500 357388
rect 200080 357348 200086 357360
rect 201494 357348 201500 357360
rect 201552 357348 201558 357400
rect 305086 357348 305092 357400
rect 305144 357388 305150 357400
rect 305730 357388 305736 357400
rect 305144 357360 305736 357388
rect 305144 357348 305150 357360
rect 305730 357348 305736 357360
rect 305788 357348 305794 357400
rect 273530 356736 273536 356788
rect 273588 356776 273594 356788
rect 274542 356776 274548 356788
rect 273588 356748 274548 356776
rect 273588 356736 273594 356748
rect 274542 356736 274548 356748
rect 274600 356736 274606 356788
rect 40034 356668 40040 356720
rect 40092 356708 40098 356720
rect 126974 356708 126980 356720
rect 40092 356680 126980 356708
rect 40092 356668 40098 356680
rect 126974 356668 126980 356680
rect 127032 356708 127038 356720
rect 214558 356708 214564 356720
rect 127032 356680 214564 356708
rect 127032 356668 127038 356680
rect 214558 356668 214564 356680
rect 214616 356668 214622 356720
rect 285674 356668 285680 356720
rect 285732 356708 285738 356720
rect 307754 356708 307760 356720
rect 285732 356680 307760 356708
rect 285732 356668 285738 356680
rect 307754 356668 307760 356680
rect 307812 356668 307818 356720
rect 253934 356396 253940 356448
rect 253992 356436 253998 356448
rect 300118 356436 300124 356448
rect 253992 356408 300124 356436
rect 253992 356396 253998 356408
rect 300118 356396 300124 356408
rect 300176 356396 300182 356448
rect 171042 356328 171048 356380
rect 171100 356368 171106 356380
rect 197722 356368 197728 356380
rect 171100 356340 197728 356368
rect 171100 356328 171106 356340
rect 197722 356328 197728 356340
rect 197780 356328 197786 356380
rect 225414 356328 225420 356380
rect 225472 356368 225478 356380
rect 303614 356368 303620 356380
rect 225472 356340 303620 356368
rect 225472 356328 225478 356340
rect 303614 356328 303620 356340
rect 303672 356328 303678 356380
rect 175918 356260 175924 356312
rect 175976 356300 175982 356312
rect 273530 356300 273536 356312
rect 175976 356272 273536 356300
rect 175976 356260 175982 356272
rect 273530 356260 273536 356272
rect 273588 356260 273594 356312
rect 68830 356192 68836 356244
rect 68888 356232 68894 356244
rect 270494 356232 270500 356244
rect 68888 356204 270500 356232
rect 68888 356192 68894 356204
rect 270494 356192 270500 356204
rect 270552 356232 270558 356244
rect 347038 356232 347044 356244
rect 270552 356204 347044 356232
rect 270552 356192 270558 356204
rect 347038 356192 347044 356204
rect 347096 356192 347102 356244
rect 67542 356124 67548 356176
rect 67600 356164 67606 356176
rect 305086 356164 305092 356176
rect 67600 356136 305092 356164
rect 67600 356124 67606 356136
rect 305086 356124 305092 356136
rect 305144 356124 305150 356176
rect 68922 356056 68928 356108
rect 68980 356096 68986 356108
rect 262766 356096 262772 356108
rect 68980 356068 262772 356096
rect 68980 356056 68986 356068
rect 262766 356056 262772 356068
rect 262824 356096 262830 356108
rect 582834 356096 582840 356108
rect 262824 356068 582840 356096
rect 262824 356056 262830 356068
rect 582834 356056 582840 356068
rect 582892 356056 582898 356108
rect 96614 355104 96620 355156
rect 96672 355144 96678 355156
rect 294046 355144 294052 355156
rect 96672 355116 294052 355144
rect 96672 355104 96678 355116
rect 294046 355104 294052 355116
rect 294104 355104 294110 355156
rect 75914 355036 75920 355088
rect 75972 355076 75978 355088
rect 293034 355076 293040 355088
rect 75972 355048 293040 355076
rect 75972 355036 75978 355048
rect 293034 355036 293040 355048
rect 293092 355036 293098 355088
rect 126422 354968 126428 355020
rect 126480 355008 126486 355020
rect 235074 355008 235080 355020
rect 126480 354980 235080 355008
rect 126480 354968 126486 354980
rect 235074 354968 235080 354980
rect 235132 354968 235138 355020
rect 107654 354900 107660 354952
rect 107712 354940 107718 354952
rect 298186 354940 298192 354952
rect 107712 354912 298192 354940
rect 107712 354900 107718 354912
rect 298186 354900 298192 354912
rect 298244 354900 298250 354952
rect 290458 354832 290464 354884
rect 290516 354872 290522 354884
rect 309778 354872 309784 354884
rect 290516 354844 309784 354872
rect 290516 354832 290522 354844
rect 309778 354832 309784 354844
rect 309836 354832 309842 354884
rect 285950 354764 285956 354816
rect 286008 354804 286014 354816
rect 311894 354804 311900 354816
rect 286008 354776 311900 354804
rect 286008 354764 286014 354776
rect 311894 354764 311900 354776
rect 311952 354764 311958 354816
rect 72418 354696 72424 354748
rect 72476 354736 72482 354748
rect 241698 354736 241704 354748
rect 72476 354708 241704 354736
rect 72476 354696 72482 354708
rect 241698 354696 241704 354708
rect 241756 354696 241762 354748
rect 260742 354696 260748 354748
rect 260800 354736 260806 354748
rect 304994 354736 305000 354748
rect 260800 354708 305000 354736
rect 260800 354696 260806 354708
rect 304994 354696 305000 354708
rect 305052 354696 305058 354748
rect 84286 354016 84292 354068
rect 84344 354056 84350 354068
rect 179782 354056 179788 354068
rect 84344 354028 179788 354056
rect 84344 354016 84350 354028
rect 179782 354016 179788 354028
rect 179840 354016 179846 354068
rect 44818 353948 44824 354000
rect 44876 353988 44882 354000
rect 45462 353988 45468 354000
rect 44876 353960 45468 353988
rect 44876 353948 44882 353960
rect 45462 353948 45468 353960
rect 45520 353988 45526 354000
rect 176654 353988 176660 354000
rect 45520 353960 176660 353988
rect 45520 353948 45526 353960
rect 176654 353948 176660 353960
rect 176712 353948 176718 354000
rect 62022 352520 62028 352572
rect 62080 352560 62086 352572
rect 176102 352560 176108 352572
rect 62080 352532 176108 352560
rect 62080 352520 62086 352532
rect 176102 352520 176108 352532
rect 176160 352520 176166 352572
rect 296162 352520 296168 352572
rect 296220 352560 296226 352572
rect 415762 352560 415768 352572
rect 296220 352532 415768 352560
rect 296220 352520 296226 352532
rect 415762 352520 415768 352532
rect 415820 352520 415826 352572
rect 117958 351228 117964 351280
rect 118016 351268 118022 351280
rect 179874 351268 179880 351280
rect 118016 351240 179880 351268
rect 118016 351228 118022 351240
rect 179874 351228 179880 351240
rect 179932 351228 179938 351280
rect 60642 351160 60648 351212
rect 60700 351200 60706 351212
rect 176010 351200 176016 351212
rect 60700 351172 176016 351200
rect 60700 351160 60706 351172
rect 176010 351160 176016 351172
rect 176068 351160 176074 351212
rect 295334 349800 295340 349852
rect 295392 349840 295398 349852
rect 359458 349840 359464 349852
rect 295392 349812 359464 349840
rect 295392 349800 295398 349812
rect 359458 349800 359464 349812
rect 359516 349800 359522 349852
rect 389082 349800 389088 349852
rect 389140 349840 389146 349852
rect 580350 349840 580356 349852
rect 389140 349812 580356 349840
rect 389140 349800 389146 349812
rect 580350 349800 580356 349812
rect 580408 349800 580414 349852
rect 124950 347760 124956 347812
rect 125008 347800 125014 347812
rect 179506 347800 179512 347812
rect 125008 347772 179512 347800
rect 125008 347760 125014 347772
rect 179506 347760 179512 347772
rect 179564 347760 179570 347812
rect 295978 346400 295984 346452
rect 296036 346440 296042 346452
rect 351178 346440 351184 346452
rect 296036 346412 351184 346440
rect 296036 346400 296042 346412
rect 351178 346400 351184 346412
rect 351236 346400 351242 346452
rect 3510 345176 3516 345228
rect 3568 345216 3574 345228
rect 8938 345216 8944 345228
rect 3568 345188 8944 345216
rect 3568 345176 3574 345188
rect 8938 345176 8944 345188
rect 8996 345176 9002 345228
rect 157242 345040 157248 345092
rect 157300 345080 157306 345092
rect 176654 345080 176660 345092
rect 157300 345052 176660 345080
rect 157300 345040 157306 345052
rect 176654 345040 176660 345052
rect 176712 345040 176718 345092
rect 296070 342864 296076 342916
rect 296128 342904 296134 342916
rect 349798 342904 349804 342916
rect 296128 342876 349804 342904
rect 296128 342864 296134 342876
rect 349798 342864 349804 342876
rect 349856 342864 349862 342916
rect 175182 342252 175188 342304
rect 175240 342292 175246 342304
rect 176838 342292 176844 342304
rect 175240 342264 176844 342292
rect 175240 342252 175246 342264
rect 176838 342252 176844 342264
rect 176896 342252 176902 342304
rect 520918 341504 520924 341556
rect 520976 341544 520982 341556
rect 536098 341544 536104 341556
rect 520976 341516 536104 341544
rect 520976 341504 520982 341516
rect 536098 341504 536104 341516
rect 536156 341504 536162 341556
rect 160738 340892 160744 340944
rect 160796 340932 160802 340944
rect 179322 340932 179328 340944
rect 160796 340904 179328 340932
rect 160796 340892 160802 340904
rect 179322 340892 179328 340904
rect 179380 340892 179386 340944
rect 295334 339464 295340 339516
rect 295392 339504 295398 339516
rect 308398 339504 308404 339516
rect 295392 339476 308404 339504
rect 295392 339464 295398 339476
rect 308398 339464 308404 339476
rect 308456 339464 308462 339516
rect 293862 338104 293868 338156
rect 293920 338144 293926 338156
rect 360838 338144 360844 338156
rect 293920 338116 360844 338144
rect 293920 338104 293926 338116
rect 360838 338104 360844 338116
rect 360896 338104 360902 338156
rect 293218 337356 293224 337408
rect 293276 337396 293282 337408
rect 498838 337396 498844 337408
rect 293276 337368 498844 337396
rect 293276 337356 293282 337368
rect 498838 337356 498844 337368
rect 498896 337356 498902 337408
rect 295334 336676 295340 336728
rect 295392 336716 295398 336728
rect 298278 336716 298284 336728
rect 295392 336688 298284 336716
rect 295392 336676 295398 336688
rect 298278 336676 298284 336688
rect 298336 336716 298342 336728
rect 299382 336716 299388 336728
rect 298336 336688 299388 336716
rect 298336 336676 298342 336688
rect 299382 336676 299388 336688
rect 299440 336676 299446 336728
rect 299382 335996 299388 336048
rect 299440 336036 299446 336048
rect 582926 336036 582932 336048
rect 299440 336008 582932 336036
rect 299440 335996 299446 336008
rect 582926 335996 582932 336008
rect 582984 335996 582990 336048
rect 106274 333956 106280 334008
rect 106332 333996 106338 334008
rect 176838 333996 176844 334008
rect 106332 333968 176844 333996
rect 106332 333956 106338 333968
rect 176838 333956 176844 333968
rect 176896 333956 176902 334008
rect 293954 333956 293960 334008
rect 294012 333996 294018 334008
rect 531958 333996 531964 334008
rect 294012 333968 531964 333996
rect 294012 333956 294018 333968
rect 531958 333956 531964 333968
rect 532016 333956 532022 334008
rect 175090 333684 175096 333736
rect 175148 333724 175154 333736
rect 176654 333724 176660 333736
rect 175148 333696 176660 333724
rect 175148 333684 175154 333696
rect 176654 333684 176660 333696
rect 176712 333684 176718 333736
rect 104158 333208 104164 333260
rect 104216 333248 104222 333260
rect 175090 333248 175096 333260
rect 104216 333220 175096 333248
rect 104216 333208 104222 333220
rect 175090 333208 175096 333220
rect 175148 333208 175154 333260
rect 295334 331848 295340 331900
rect 295392 331888 295398 331900
rect 296898 331888 296904 331900
rect 295392 331860 296904 331888
rect 295392 331848 295398 331860
rect 296898 331848 296904 331860
rect 296956 331888 296962 331900
rect 367738 331888 367744 331900
rect 296956 331860 367744 331888
rect 296956 331848 296962 331860
rect 367738 331848 367744 331860
rect 367796 331848 367802 331900
rect 294322 329808 294328 329860
rect 294380 329848 294386 329860
rect 369118 329848 369124 329860
rect 294380 329820 369124 329848
rect 294380 329808 294386 329820
rect 369118 329808 369124 329820
rect 369176 329808 369182 329860
rect 175090 327088 175096 327140
rect 175148 327128 175154 327140
rect 176654 327128 176660 327140
rect 175148 327100 176660 327128
rect 175148 327088 175154 327100
rect 176654 327088 176660 327100
rect 176712 327088 176718 327140
rect 293034 327088 293040 327140
rect 293092 327128 293098 327140
rect 575566 327128 575572 327140
rect 293092 327100 575572 327128
rect 293092 327088 293098 327100
rect 575566 327088 575572 327100
rect 575624 327088 575630 327140
rect 151722 325660 151728 325712
rect 151780 325700 151786 325712
rect 176654 325700 176660 325712
rect 151780 325672 176660 325700
rect 151780 325660 151786 325672
rect 176654 325660 176660 325672
rect 176712 325660 176718 325712
rect 3418 324912 3424 324964
rect 3476 324952 3482 324964
rect 98638 324952 98644 324964
rect 3476 324924 98644 324952
rect 3476 324912 3482 324924
rect 98638 324912 98644 324924
rect 98696 324912 98702 324964
rect 573542 324300 573548 324352
rect 573600 324340 573606 324352
rect 580166 324340 580172 324352
rect 573600 324312 580172 324340
rect 573600 324300 573606 324312
rect 580166 324300 580172 324312
rect 580224 324300 580230 324352
rect 295334 320152 295340 320204
rect 295392 320192 295398 320204
rect 323578 320192 323584 320204
rect 295392 320164 323584 320192
rect 295392 320152 295398 320164
rect 323578 320152 323584 320164
rect 323636 320152 323642 320204
rect 3418 318792 3424 318844
rect 3476 318832 3482 318844
rect 116578 318832 116584 318844
rect 3476 318804 116584 318832
rect 3476 318792 3482 318804
rect 116578 318792 116584 318804
rect 116636 318792 116642 318844
rect 295334 318792 295340 318844
rect 295392 318832 295398 318844
rect 325050 318832 325056 318844
rect 295392 318804 325056 318832
rect 295392 318792 295398 318804
rect 325050 318792 325056 318804
rect 325108 318792 325114 318844
rect 295334 317364 295340 317416
rect 295392 317404 295398 317416
rect 299566 317404 299572 317416
rect 295392 317376 299572 317404
rect 295392 317364 295398 317376
rect 299566 317364 299572 317376
rect 299624 317404 299630 317416
rect 300762 317404 300768 317416
rect 299624 317376 300768 317404
rect 299624 317364 299630 317376
rect 300762 317364 300768 317376
rect 300820 317364 300826 317416
rect 300762 316684 300768 316736
rect 300820 316724 300826 316736
rect 337470 316724 337476 316736
rect 300820 316696 337476 316724
rect 300820 316684 300826 316696
rect 337470 316684 337476 316696
rect 337528 316684 337534 316736
rect 129274 314644 129280 314696
rect 129332 314684 129338 314696
rect 176654 314684 176660 314696
rect 129332 314656 176660 314684
rect 129332 314644 129338 314656
rect 176654 314644 176660 314656
rect 176712 314644 176718 314696
rect 295334 313896 295340 313948
rect 295392 313936 295398 313948
rect 296806 313936 296812 313948
rect 295392 313908 296812 313936
rect 295392 313896 295398 313908
rect 296806 313896 296812 313908
rect 296864 313936 296870 313948
rect 570046 313936 570052 313948
rect 296864 313908 570052 313936
rect 296864 313896 296870 313908
rect 570046 313896 570052 313908
rect 570104 313896 570110 313948
rect 160554 312536 160560 312588
rect 160612 312576 160618 312588
rect 176654 312576 176660 312588
rect 160612 312548 176660 312576
rect 160612 312536 160618 312548
rect 176654 312536 176660 312548
rect 176712 312536 176718 312588
rect 99374 311856 99380 311908
rect 99432 311896 99438 311908
rect 160554 311896 160560 311908
rect 99432 311868 160560 311896
rect 99432 311856 99438 311868
rect 160554 311856 160560 311868
rect 160612 311856 160618 311908
rect 295334 311856 295340 311908
rect 295392 311896 295398 311908
rect 471238 311896 471244 311908
rect 295392 311868 471244 311896
rect 295392 311856 295398 311868
rect 471238 311856 471244 311868
rect 471296 311856 471302 311908
rect 8938 311108 8944 311160
rect 8996 311148 9002 311160
rect 118694 311148 118700 311160
rect 8996 311120 118700 311148
rect 8996 311108 9002 311120
rect 118694 311108 118700 311120
rect 118752 311108 118758 311160
rect 122098 311108 122104 311160
rect 122156 311148 122162 311160
rect 160738 311148 160744 311160
rect 122156 311120 160744 311148
rect 122156 311108 122162 311120
rect 160738 311108 160744 311120
rect 160796 311108 160802 311160
rect 118694 310428 118700 310480
rect 118752 310468 118758 310480
rect 173158 310468 173164 310480
rect 118752 310440 173164 310468
rect 118752 310428 118758 310440
rect 173158 310428 173164 310440
rect 173216 310428 173222 310480
rect 295334 310428 295340 310480
rect 295392 310468 295398 310480
rect 300946 310468 300952 310480
rect 295392 310440 300952 310468
rect 295392 310428 295398 310440
rect 300946 310428 300952 310440
rect 301004 310468 301010 310480
rect 301314 310468 301320 310480
rect 301004 310440 301320 310468
rect 301004 310428 301010 310440
rect 301314 310428 301320 310440
rect 301372 310428 301378 310480
rect 301314 309748 301320 309800
rect 301372 309788 301378 309800
rect 468478 309788 468484 309800
rect 301372 309760 468484 309788
rect 301372 309748 301378 309760
rect 468478 309748 468484 309760
rect 468536 309748 468542 309800
rect 295334 307776 295340 307828
rect 295392 307816 295398 307828
rect 313274 307816 313280 307828
rect 295392 307788 313280 307816
rect 295392 307776 295398 307788
rect 313274 307776 313280 307788
rect 313332 307816 313338 307828
rect 570230 307816 570236 307828
rect 313332 307788 570236 307816
rect 313332 307776 313338 307788
rect 570230 307776 570236 307788
rect 570288 307776 570294 307828
rect 25498 307028 25504 307080
rect 25556 307068 25562 307080
rect 84378 307068 84384 307080
rect 25556 307040 84384 307068
rect 25556 307028 25562 307040
rect 84378 307028 84384 307040
rect 84436 307028 84442 307080
rect 91094 307028 91100 307080
rect 91152 307068 91158 307080
rect 99374 307068 99380 307080
rect 91152 307040 99380 307068
rect 91152 307028 91158 307040
rect 99374 307028 99380 307040
rect 99432 307028 99438 307080
rect 154390 307028 154396 307080
rect 154448 307068 154454 307080
rect 176470 307068 176476 307080
rect 154448 307040 176476 307068
rect 154448 307028 154454 307040
rect 176470 307028 176476 307040
rect 176528 307028 176534 307080
rect 114738 306348 114744 306400
rect 114796 306388 114802 306400
rect 154390 306388 154396 306400
rect 114796 306360 154396 306388
rect 114796 306348 114802 306360
rect 154390 306348 154396 306360
rect 154448 306348 154454 306400
rect 81434 305124 81440 305176
rect 81492 305164 81498 305176
rect 138750 305164 138756 305176
rect 81492 305136 138756 305164
rect 81492 305124 81498 305136
rect 138750 305124 138756 305136
rect 138808 305124 138814 305176
rect 88426 305056 88432 305108
rect 88484 305096 88490 305108
rect 162118 305096 162124 305108
rect 88484 305068 162124 305096
rect 88484 305056 88490 305068
rect 162118 305056 162124 305068
rect 162176 305056 162182 305108
rect 3234 304988 3240 305040
rect 3292 305028 3298 305040
rect 122190 305028 122196 305040
rect 3292 305000 122196 305028
rect 3292 304988 3298 305000
rect 122190 304988 122196 305000
rect 122248 305028 122254 305040
rect 173802 305028 173808 305040
rect 122248 305000 173808 305028
rect 122248 304988 122254 305000
rect 173802 304988 173808 305000
rect 173860 305028 173866 305040
rect 176654 305028 176660 305040
rect 173860 305000 176660 305028
rect 173860 304988 173866 305000
rect 176654 304988 176660 305000
rect 176712 304988 176718 305040
rect 295334 304988 295340 305040
rect 295392 305028 295398 305040
rect 310606 305028 310612 305040
rect 295392 305000 310612 305028
rect 295392 304988 295398 305000
rect 310606 304988 310612 305000
rect 310664 304988 310670 305040
rect 13078 304920 13084 304972
rect 13136 304960 13142 304972
rect 72234 304960 72240 304972
rect 13136 304932 72240 304960
rect 13136 304920 13142 304932
rect 72234 304920 72240 304932
rect 72292 304920 72298 304972
rect 94498 304920 94504 304972
rect 94556 304960 94562 304972
rect 114738 304960 114744 304972
rect 94556 304932 114744 304960
rect 94556 304920 94562 304932
rect 114738 304920 114744 304932
rect 114796 304920 114802 304972
rect 90358 304716 90364 304768
rect 90416 304756 90422 304768
rect 94590 304756 94596 304768
rect 90416 304728 94596 304756
rect 90416 304716 90422 304728
rect 94590 304716 94596 304728
rect 94648 304716 94654 304768
rect 388990 304240 388996 304292
rect 389048 304280 389054 304292
rect 542354 304280 542360 304292
rect 389048 304252 542360 304280
rect 389048 304240 389054 304252
rect 542354 304240 542360 304252
rect 542412 304240 542418 304292
rect 74534 303628 74540 303680
rect 74592 303668 74598 303680
rect 142890 303668 142896 303680
rect 74592 303640 142896 303668
rect 74592 303628 74598 303640
rect 142890 303628 142896 303640
rect 142948 303628 142954 303680
rect 88334 303560 88340 303612
rect 88392 303600 88398 303612
rect 103790 303600 103796 303612
rect 88392 303572 103796 303600
rect 88392 303560 88398 303572
rect 103790 303560 103796 303572
rect 103848 303600 103854 303612
rect 104158 303600 104164 303612
rect 103848 303572 104164 303600
rect 103848 303560 103854 303572
rect 104158 303560 104164 303572
rect 104216 303560 104222 303612
rect 295334 303560 295340 303612
rect 295392 303600 295398 303612
rect 298186 303600 298192 303612
rect 295392 303572 298192 303600
rect 295392 303560 295398 303572
rect 298186 303560 298192 303572
rect 298244 303600 298250 303612
rect 412634 303600 412640 303612
rect 298244 303572 412640 303600
rect 298244 303560 298250 303572
rect 412634 303560 412640 303572
rect 412692 303600 412698 303612
rect 413278 303600 413284 303612
rect 412692 303572 413284 303600
rect 412692 303560 412698 303572
rect 413278 303560 413284 303572
rect 413336 303560 413342 303612
rect 89714 302404 89720 302456
rect 89772 302444 89778 302456
rect 134702 302444 134708 302456
rect 89772 302416 134708 302444
rect 89772 302404 89778 302416
rect 134702 302404 134708 302416
rect 134760 302404 134766 302456
rect 99374 302336 99380 302388
rect 99432 302376 99438 302388
rect 148318 302376 148324 302388
rect 99432 302348 148324 302376
rect 99432 302336 99438 302348
rect 148318 302336 148324 302348
rect 148376 302336 148382 302388
rect 92842 302268 92848 302320
rect 92900 302308 92906 302320
rect 152550 302308 152556 302320
rect 92900 302280 152556 302308
rect 92900 302268 92906 302280
rect 152550 302268 152556 302280
rect 152608 302268 152614 302320
rect 98730 302200 98736 302252
rect 98788 302240 98794 302252
rect 178678 302240 178684 302252
rect 98788 302212 178684 302240
rect 98788 302200 98794 302212
rect 178678 302200 178684 302212
rect 178736 302200 178742 302252
rect 104158 301180 104164 301232
rect 104216 301220 104222 301232
rect 144178 301220 144184 301232
rect 104216 301192 144184 301220
rect 104216 301180 104222 301192
rect 144178 301180 144184 301192
rect 144236 301180 144242 301232
rect 102134 301112 102140 301164
rect 102192 301152 102198 301164
rect 149790 301152 149796 301164
rect 102192 301124 149796 301152
rect 102192 301112 102198 301124
rect 149790 301112 149796 301124
rect 149848 301112 149854 301164
rect 76098 301044 76104 301096
rect 76156 301084 76162 301096
rect 130562 301084 130568 301096
rect 76156 301056 130568 301084
rect 76156 301044 76162 301056
rect 130562 301044 130568 301056
rect 130620 301044 130626 301096
rect 85574 300976 85580 301028
rect 85632 301016 85638 301028
rect 153838 301016 153844 301028
rect 85632 300988 153844 301016
rect 85632 300976 85638 300988
rect 153838 300976 153844 300988
rect 153896 300976 153902 301028
rect 85666 300908 85672 300960
rect 85724 300948 85730 300960
rect 155218 300948 155224 300960
rect 85724 300920 155224 300948
rect 85724 300908 85730 300920
rect 155218 300908 155224 300920
rect 155276 300908 155282 300960
rect 160002 300908 160008 300960
rect 160060 300948 160066 300960
rect 176654 300948 176660 300960
rect 160060 300920 176660 300948
rect 160060 300908 160066 300920
rect 176654 300908 176660 300920
rect 176712 300908 176718 300960
rect 75362 300840 75368 300892
rect 75420 300880 75426 300892
rect 165062 300880 165068 300892
rect 75420 300852 165068 300880
rect 75420 300840 75426 300852
rect 165062 300840 165068 300852
rect 165120 300840 165126 300892
rect 293218 300840 293224 300892
rect 293276 300880 293282 300892
rect 300210 300880 300216 300892
rect 293276 300852 300216 300880
rect 293276 300840 293282 300852
rect 300210 300840 300216 300852
rect 300268 300840 300274 300892
rect 97994 300772 98000 300824
rect 98052 300812 98058 300824
rect 98638 300812 98644 300824
rect 98052 300784 98644 300812
rect 98052 300772 98058 300784
rect 98638 300772 98644 300784
rect 98696 300772 98702 300824
rect 53742 300092 53748 300144
rect 53800 300132 53806 300144
rect 70946 300132 70952 300144
rect 53800 300104 70952 300132
rect 53800 300092 53806 300104
rect 70946 300092 70952 300104
rect 71004 300092 71010 300144
rect 296070 300092 296076 300144
rect 296128 300132 296134 300144
rect 305086 300132 305092 300144
rect 296128 300104 305092 300132
rect 296128 300092 296134 300104
rect 305086 300092 305092 300104
rect 305144 300092 305150 300144
rect 88334 299752 88340 299804
rect 88392 299792 88398 299804
rect 123478 299792 123484 299804
rect 88392 299764 123484 299792
rect 88392 299752 88398 299764
rect 123478 299752 123484 299764
rect 123536 299752 123542 299804
rect 98546 299684 98552 299736
rect 98604 299724 98610 299736
rect 136082 299724 136088 299736
rect 98604 299696 136088 299724
rect 98604 299684 98610 299696
rect 136082 299684 136088 299696
rect 136140 299684 136146 299736
rect 97994 299616 98000 299668
rect 98052 299656 98058 299668
rect 148410 299656 148416 299668
rect 98052 299628 148416 299656
rect 98052 299616 98058 299628
rect 148410 299616 148416 299628
rect 148468 299616 148474 299668
rect 84378 299548 84384 299600
rect 84436 299588 84442 299600
rect 144362 299588 144368 299600
rect 84436 299560 144368 299588
rect 84436 299548 84442 299560
rect 144362 299548 144368 299560
rect 144420 299548 144426 299600
rect 22830 299480 22836 299532
rect 22888 299520 22894 299532
rect 117958 299520 117964 299532
rect 22888 299492 117964 299520
rect 22888 299480 22894 299492
rect 117958 299480 117964 299492
rect 118016 299480 118022 299532
rect 111058 298732 111064 298784
rect 111116 298772 111122 298784
rect 124214 298772 124220 298784
rect 111116 298744 124220 298772
rect 111116 298732 111122 298744
rect 124214 298732 124220 298744
rect 124272 298732 124278 298784
rect 102870 298392 102876 298444
rect 102928 298432 102934 298444
rect 124858 298432 124864 298444
rect 102928 298404 124864 298432
rect 102928 298392 102934 298404
rect 124858 298392 124864 298404
rect 124916 298392 124922 298444
rect 90634 298324 90640 298376
rect 90692 298364 90698 298376
rect 137278 298364 137284 298376
rect 90692 298336 137284 298364
rect 90692 298324 90698 298336
rect 137278 298324 137284 298336
rect 137336 298324 137342 298376
rect 116578 298256 116584 298308
rect 116636 298296 116642 298308
rect 169110 298296 169116 298308
rect 116636 298268 169116 298296
rect 116636 298256 116642 298268
rect 169110 298256 169116 298268
rect 169168 298256 169174 298308
rect 75178 298188 75184 298240
rect 75236 298228 75242 298240
rect 131758 298228 131764 298240
rect 75236 298200 131764 298228
rect 75236 298188 75242 298200
rect 131758 298188 131764 298200
rect 131816 298188 131822 298240
rect 73246 298120 73252 298172
rect 73304 298160 73310 298172
rect 159358 298160 159364 298172
rect 73304 298132 159364 298160
rect 73304 298120 73310 298132
rect 159358 298120 159364 298132
rect 159416 298120 159422 298172
rect 169754 298052 169760 298104
rect 169812 298092 169818 298104
rect 170950 298092 170956 298104
rect 169812 298064 170956 298092
rect 169812 298052 169818 298064
rect 170950 298052 170956 298064
rect 171008 298092 171014 298104
rect 176654 298092 176660 298104
rect 171008 298064 176660 298092
rect 171008 298052 171014 298064
rect 176654 298052 176660 298064
rect 176712 298052 176718 298104
rect 502334 298052 502340 298104
rect 502392 298092 502398 298104
rect 502978 298092 502984 298104
rect 502392 298064 502984 298092
rect 502392 298052 502398 298064
rect 502978 298052 502984 298064
rect 503036 298052 503042 298104
rect 158438 297372 158444 297424
rect 158496 297412 158502 297424
rect 176654 297412 176660 297424
rect 158496 297384 176660 297412
rect 158496 297372 158502 297384
rect 176654 297372 176660 297384
rect 176712 297372 176718 297424
rect 129642 297032 129648 297084
rect 129700 297072 129706 297084
rect 158438 297072 158444 297084
rect 129700 297044 158444 297072
rect 129700 297032 129706 297044
rect 158438 297032 158444 297044
rect 158496 297032 158502 297084
rect 87414 296964 87420 297016
rect 87472 297004 87478 297016
rect 133230 297004 133236 297016
rect 87472 296976 133236 297004
rect 87472 296964 87478 296976
rect 133230 296964 133236 296976
rect 133288 296964 133294 297016
rect 83550 296896 83556 296948
rect 83608 296936 83614 296948
rect 133138 296936 133144 296948
rect 83608 296908 133144 296936
rect 83608 296896 83614 296908
rect 133138 296896 133144 296908
rect 133196 296896 133202 296948
rect 104342 296828 104348 296880
rect 104400 296868 104406 296880
rect 156690 296868 156696 296880
rect 104400 296840 156696 296868
rect 104400 296828 104406 296840
rect 156690 296828 156696 296840
rect 156748 296828 156754 296880
rect 66162 296760 66168 296812
rect 66220 296800 66226 296812
rect 140222 296800 140228 296812
rect 66220 296772 140228 296800
rect 66220 296760 66226 296772
rect 140222 296760 140228 296772
rect 140280 296760 140286 296812
rect 68554 296692 68560 296744
rect 68612 296732 68618 296744
rect 157334 296732 157340 296744
rect 68612 296704 157340 296732
rect 68612 296692 68618 296704
rect 157334 296692 157340 296704
rect 157392 296692 157398 296744
rect 327718 296692 327724 296744
rect 327776 296732 327782 296744
rect 502334 296732 502340 296744
rect 327776 296704 502340 296732
rect 327776 296692 327782 296704
rect 502334 296692 502340 296704
rect 502392 296692 502398 296744
rect 84194 295672 84200 295724
rect 84252 295712 84258 295724
rect 84470 295712 84476 295724
rect 84252 295684 84476 295712
rect 84252 295672 84258 295684
rect 84470 295672 84476 295684
rect 84528 295672 84534 295724
rect 111886 295672 111892 295724
rect 111944 295712 111950 295724
rect 151170 295712 151176 295724
rect 111944 295684 151176 295712
rect 111944 295672 111950 295684
rect 151170 295672 151176 295684
rect 151228 295672 151234 295724
rect 78398 295604 78404 295656
rect 78456 295644 78462 295656
rect 78456 295616 93854 295644
rect 78456 295604 78462 295616
rect 82262 295536 82268 295588
rect 82320 295576 82326 295588
rect 88978 295576 88984 295588
rect 82320 295548 88984 295576
rect 82320 295536 82326 295548
rect 88978 295536 88984 295548
rect 89036 295536 89042 295588
rect 93826 295576 93854 295616
rect 117222 295604 117228 295656
rect 117280 295644 117286 295656
rect 164970 295644 164976 295656
rect 117280 295616 164976 295644
rect 117280 295604 117286 295616
rect 164970 295604 164976 295616
rect 165028 295604 165034 295656
rect 137370 295576 137376 295588
rect 93826 295548 137376 295576
rect 137370 295536 137376 295548
rect 137428 295536 137434 295588
rect 84470 295468 84476 295520
rect 84528 295508 84534 295520
rect 145558 295508 145564 295520
rect 84528 295480 145564 295508
rect 84528 295468 84534 295480
rect 145558 295468 145564 295480
rect 145616 295468 145622 295520
rect 32398 295400 32404 295452
rect 32456 295440 32462 295452
rect 101398 295440 101404 295452
rect 32456 295412 84194 295440
rect 32456 295400 32462 295412
rect 84166 295372 84194 295412
rect 84488 295412 101404 295440
rect 84166 295344 84332 295372
rect 84304 295304 84332 295344
rect 84488 295304 84516 295412
rect 101398 295400 101404 295412
rect 101456 295400 101462 295452
rect 105446 295400 105452 295452
rect 105504 295440 105510 295452
rect 171134 295440 171140 295452
rect 105504 295412 171140 295440
rect 105504 295400 105510 295412
rect 171134 295400 171140 295412
rect 171192 295400 171198 295452
rect 88978 295332 88984 295384
rect 89036 295372 89042 295384
rect 156598 295372 156604 295384
rect 89036 295344 156604 295372
rect 89036 295332 89042 295344
rect 156598 295332 156604 295344
rect 156656 295332 156662 295384
rect 295334 295332 295340 295384
rect 295392 295372 295398 295384
rect 302878 295372 302884 295384
rect 295392 295344 302884 295372
rect 295392 295332 295398 295344
rect 302878 295332 302884 295344
rect 302936 295332 302942 295384
rect 84304 295276 84516 295304
rect 79686 294652 79692 294704
rect 79744 294692 79750 294704
rect 104158 294692 104164 294704
rect 79744 294664 104164 294692
rect 79744 294652 79750 294664
rect 104158 294652 104164 294664
rect 104216 294652 104222 294704
rect 70026 294584 70032 294636
rect 70084 294624 70090 294636
rect 117222 294624 117228 294636
rect 70084 294596 117228 294624
rect 70084 294584 70090 294596
rect 117222 294584 117228 294596
rect 117280 294584 117286 294636
rect 300210 294584 300216 294636
rect 300268 294624 300274 294636
rect 492398 294624 492404 294636
rect 300268 294596 492404 294624
rect 300268 294584 300274 294596
rect 492398 294584 492404 294596
rect 492456 294584 492462 294636
rect 80974 294380 80980 294432
rect 81032 294420 81038 294432
rect 135990 294420 135996 294432
rect 81032 294392 135996 294420
rect 81032 294380 81038 294392
rect 135990 294380 135996 294392
rect 136048 294380 136054 294432
rect 106090 294312 106096 294364
rect 106148 294352 106154 294364
rect 123570 294352 123576 294364
rect 106148 294324 123576 294352
rect 106148 294312 106154 294324
rect 123570 294312 123576 294324
rect 123628 294312 123634 294364
rect 114462 294244 114468 294296
rect 114520 294284 114526 294296
rect 140130 294284 140136 294296
rect 114520 294256 140136 294284
rect 114520 294244 114526 294256
rect 140130 294244 140136 294256
rect 140188 294244 140194 294296
rect 82906 294176 82912 294228
rect 82964 294216 82970 294228
rect 116854 294216 116860 294228
rect 82964 294188 116860 294216
rect 82964 294176 82970 294188
rect 116854 294176 116860 294188
rect 116912 294176 116918 294228
rect 93854 294108 93860 294160
rect 93912 294148 93918 294160
rect 138842 294148 138848 294160
rect 93912 294120 138848 294148
rect 93912 294108 93918 294120
rect 138842 294108 138848 294120
rect 138900 294108 138906 294160
rect 67450 294040 67456 294092
rect 67508 294080 67514 294092
rect 79318 294080 79324 294092
rect 67508 294052 79324 294080
rect 67508 294040 67514 294052
rect 79318 294040 79324 294052
rect 79376 294040 79382 294092
rect 49602 293972 49608 294024
rect 49660 294012 49666 294024
rect 96430 294012 96436 294024
rect 49660 293984 96436 294012
rect 49660 293972 49666 293984
rect 96430 293972 96436 293984
rect 96488 293972 96494 294024
rect 103790 293972 103796 294024
rect 103848 294012 103854 294024
rect 104526 294012 104532 294024
rect 103848 293984 104532 294012
rect 103848 293972 103854 293984
rect 104526 293972 104532 293984
rect 104584 293972 104590 294024
rect 114554 293972 114560 294024
rect 114612 294012 114618 294024
rect 115382 294012 115388 294024
rect 114612 293984 115388 294012
rect 114612 293972 114618 293984
rect 115382 293972 115388 293984
rect 115440 293972 115446 294024
rect 117222 293972 117228 294024
rect 117280 294012 117286 294024
rect 173158 294012 173164 294024
rect 117280 293984 173164 294012
rect 117280 293972 117286 293984
rect 173158 293972 173164 293984
rect 173216 293972 173222 294024
rect 295334 293972 295340 294024
rect 295392 294012 295398 294024
rect 302142 294012 302148 294024
rect 295392 293984 302148 294012
rect 295392 293972 295398 293984
rect 302142 293972 302148 293984
rect 302200 293972 302206 294024
rect 75914 293904 75920 293956
rect 75972 293944 75978 293956
rect 76742 293944 76748 293956
rect 75972 293916 76748 293944
rect 75972 293904 75978 293916
rect 76742 293904 76748 293916
rect 76800 293904 76806 293956
rect 84286 293904 84292 293956
rect 84344 293944 84350 293956
rect 85206 293944 85212 293956
rect 84344 293916 85212 293944
rect 84344 293904 84350 293916
rect 85206 293904 85212 293916
rect 85264 293904 85270 293956
rect 85574 293904 85580 293956
rect 85632 293944 85638 293956
rect 86494 293944 86500 293956
rect 85632 293916 86500 293944
rect 85632 293904 85638 293916
rect 86494 293904 86500 293916
rect 86552 293904 86558 293956
rect 88334 293904 88340 293956
rect 88392 293944 88398 293956
rect 89070 293944 89076 293956
rect 88392 293916 89076 293944
rect 88392 293904 88398 293916
rect 89070 293904 89076 293916
rect 89128 293904 89134 293956
rect 92566 292884 92572 292936
rect 92624 292924 92630 292936
rect 120994 292924 121000 292936
rect 92624 292896 121000 292924
rect 92624 292884 92630 292896
rect 120994 292884 121000 292896
rect 121052 292884 121058 292936
rect 110598 292816 110604 292868
rect 110656 292856 110662 292868
rect 126330 292856 126336 292868
rect 110656 292828 126336 292856
rect 110656 292816 110662 292828
rect 126330 292816 126336 292828
rect 126388 292816 126394 292868
rect 88058 292748 88064 292800
rect 88116 292788 88122 292800
rect 129090 292788 129096 292800
rect 88116 292760 129096 292788
rect 88116 292748 88122 292760
rect 129090 292748 129096 292760
rect 129148 292748 129154 292800
rect 53650 292680 53656 292732
rect 53708 292720 53714 292732
rect 71958 292720 71964 292732
rect 53708 292692 71964 292720
rect 53708 292680 53714 292692
rect 71958 292680 71964 292692
rect 72016 292680 72022 292732
rect 91922 292680 91928 292732
rect 91980 292720 91986 292732
rect 134610 292720 134616 292732
rect 91980 292692 134616 292720
rect 91980 292680 91986 292692
rect 134610 292680 134616 292692
rect 134668 292680 134674 292732
rect 53098 292612 53104 292664
rect 53156 292652 53162 292664
rect 92566 292652 92572 292664
rect 53156 292624 92572 292652
rect 53156 292612 53162 292624
rect 92566 292612 92572 292624
rect 92624 292612 92630 292664
rect 109310 292612 109316 292664
rect 109368 292652 109374 292664
rect 162210 292652 162216 292664
rect 109368 292624 162216 292652
rect 109368 292612 109374 292624
rect 162210 292612 162216 292624
rect 162268 292612 162274 292664
rect 3418 292544 3424 292596
rect 3476 292584 3482 292596
rect 46198 292584 46204 292596
rect 3476 292556 46204 292584
rect 3476 292544 3482 292556
rect 46198 292544 46204 292556
rect 46256 292544 46262 292596
rect 68738 292544 68744 292596
rect 68796 292584 68802 292596
rect 141510 292584 141516 292596
rect 68796 292556 141516 292584
rect 68796 292544 68802 292556
rect 141510 292544 141516 292556
rect 141568 292544 141574 292596
rect 319530 292544 319536 292596
rect 319588 292584 319594 292596
rect 520734 292584 520740 292596
rect 319588 292556 520740 292584
rect 319588 292544 319594 292556
rect 520734 292544 520740 292556
rect 520792 292544 520798 292596
rect 71682 292476 71688 292528
rect 71740 292516 71746 292528
rect 111150 292516 111156 292528
rect 71740 292488 111156 292516
rect 71740 292476 71746 292488
rect 111150 292476 111156 292488
rect 111208 292476 111214 292528
rect 121454 292476 121460 292528
rect 121512 292516 121518 292528
rect 126422 292516 126428 292528
rect 121512 292488 126428 292516
rect 121512 292476 121518 292488
rect 126422 292476 126428 292488
rect 126480 292476 126486 292528
rect 117314 291932 117320 291984
rect 117372 291972 117378 291984
rect 119706 291972 119712 291984
rect 117372 291944 119712 291972
rect 117372 291932 117378 291944
rect 119706 291932 119712 291944
rect 119764 291932 119770 291984
rect 101306 291864 101312 291916
rect 101364 291904 101370 291916
rect 101364 291876 103514 291904
rect 101364 291864 101370 291876
rect 103486 291224 103514 291876
rect 112806 291864 112812 291916
rect 112864 291904 112870 291916
rect 112864 291876 113174 291904
rect 112864 291864 112870 291876
rect 113146 291292 113174 291876
rect 116854 291864 116860 291916
rect 116912 291864 116918 291916
rect 119338 291864 119344 291916
rect 119396 291904 119402 291916
rect 119982 291904 119988 291916
rect 119396 291876 119988 291904
rect 119396 291864 119402 291876
rect 119982 291864 119988 291876
rect 120040 291864 120046 291916
rect 116872 291836 116900 291864
rect 147030 291836 147036 291848
rect 116872 291808 147036 291836
rect 147030 291796 147036 291808
rect 147088 291796 147094 291848
rect 160738 291796 160744 291848
rect 160796 291836 160802 291848
rect 176654 291836 176660 291848
rect 160796 291808 176660 291836
rect 160796 291796 160802 291808
rect 176654 291796 176660 291808
rect 176712 291796 176718 291848
rect 119982 291320 119988 291372
rect 120040 291360 120046 291372
rect 129182 291360 129188 291372
rect 120040 291332 129188 291360
rect 120040 291320 120046 291332
rect 129182 291320 129188 291332
rect 129240 291320 129246 291372
rect 583846 291360 583852 291372
rect 567166 291332 583852 291360
rect 127710 291292 127716 291304
rect 113146 291264 127716 291292
rect 127710 291252 127716 291264
rect 127768 291252 127774 291304
rect 345658 291252 345664 291304
rect 345716 291292 345722 291304
rect 567166 291292 567194 291332
rect 583846 291320 583852 291332
rect 583904 291320 583910 291372
rect 345716 291264 567194 291292
rect 345716 291252 345722 291264
rect 131850 291224 131856 291236
rect 103486 291196 131856 291224
rect 131850 291184 131856 291196
rect 131908 291184 131914 291236
rect 323670 291184 323676 291236
rect 323728 291224 323734 291236
rect 566458 291224 566464 291236
rect 323728 291196 566464 291224
rect 323728 291184 323734 291196
rect 566458 291184 566464 291196
rect 566516 291184 566522 291236
rect 31018 290436 31024 290488
rect 31076 290476 31082 290488
rect 68738 290476 68744 290488
rect 31076 290448 68744 290476
rect 31076 290436 31082 290448
rect 68738 290436 68744 290448
rect 68796 290436 68802 290488
rect 362218 289960 362224 290012
rect 362276 290000 362282 290012
rect 533614 290000 533620 290012
rect 362276 289972 533620 290000
rect 362276 289960 362282 289972
rect 533614 289960 533620 289972
rect 533672 289960 533678 290012
rect 121454 289892 121460 289944
rect 121512 289932 121518 289944
rect 149698 289932 149704 289944
rect 121512 289904 149704 289932
rect 121512 289892 121518 289904
rect 149698 289892 149704 289904
rect 149756 289892 149762 289944
rect 318150 289892 318156 289944
rect 318208 289932 318214 289944
rect 583662 289932 583668 289944
rect 318208 289904 583668 289932
rect 318208 289892 318214 289904
rect 583662 289892 583668 289904
rect 583720 289892 583726 289944
rect 56410 289824 56416 289876
rect 56468 289864 56474 289876
rect 67634 289864 67640 289876
rect 56468 289836 67640 289864
rect 56468 289824 56474 289836
rect 67634 289824 67640 289836
rect 67692 289824 67698 289876
rect 121546 289824 121552 289876
rect 121604 289864 121610 289876
rect 164878 289864 164884 289876
rect 121604 289836 164884 289864
rect 121604 289824 121610 289836
rect 164878 289824 164884 289836
rect 164936 289824 164942 289876
rect 169018 289824 169024 289876
rect 169076 289864 169082 289876
rect 176654 289864 176660 289876
rect 169076 289836 176660 289864
rect 169076 289824 169082 289836
rect 176654 289824 176660 289836
rect 176712 289824 176718 289876
rect 302142 289824 302148 289876
rect 302200 289864 302206 289876
rect 449894 289864 449900 289876
rect 302200 289836 449900 289864
rect 302200 289824 302206 289836
rect 449894 289824 449900 289836
rect 449952 289824 449958 289876
rect 121454 289756 121460 289808
rect 121512 289796 121518 289808
rect 162302 289796 162308 289808
rect 121512 289768 162308 289796
rect 121512 289756 121518 289768
rect 162302 289756 162308 289768
rect 162360 289756 162366 289808
rect 4062 289076 4068 289128
rect 4120 289116 4126 289128
rect 67450 289116 67456 289128
rect 4120 289088 67456 289116
rect 4120 289076 4126 289088
rect 67450 289076 67456 289088
rect 67508 289076 67514 289128
rect 369302 288532 369308 288584
rect 369360 288572 369366 288584
rect 418982 288572 418988 288584
rect 369360 288544 418988 288572
rect 369360 288532 369366 288544
rect 418982 288532 418988 288544
rect 419040 288532 419046 288584
rect 52362 288464 52368 288516
rect 52420 288504 52426 288516
rect 67726 288504 67732 288516
rect 52420 288476 67732 288504
rect 52420 288464 52426 288476
rect 67726 288464 67732 288476
rect 67784 288464 67790 288516
rect 385862 288464 385868 288516
rect 385920 288504 385926 288516
rect 566550 288504 566556 288516
rect 385920 288476 566556 288504
rect 385920 288464 385926 288476
rect 566550 288464 566556 288476
rect 566608 288464 566614 288516
rect 50982 288396 50988 288448
rect 51040 288436 51046 288448
rect 67634 288436 67640 288448
rect 51040 288408 67640 288436
rect 51040 288396 51046 288408
rect 67634 288396 67640 288408
rect 67692 288396 67698 288448
rect 356790 288396 356796 288448
rect 356848 288436 356854 288448
rect 583570 288436 583576 288448
rect 356848 288408 583576 288436
rect 356848 288396 356854 288408
rect 583570 288396 583576 288408
rect 583628 288396 583634 288448
rect 121454 288328 121460 288380
rect 121512 288368 121518 288380
rect 126238 288368 126244 288380
rect 121512 288340 126244 288368
rect 121512 288328 121518 288340
rect 126238 288328 126244 288340
rect 126296 288328 126302 288380
rect 296714 287648 296720 287700
rect 296772 287688 296778 287700
rect 406102 287688 406108 287700
rect 296772 287660 406108 287688
rect 296772 287648 296778 287660
rect 406102 287648 406108 287660
rect 406160 287648 406166 287700
rect 413278 287648 413284 287700
rect 413336 287688 413342 287700
rect 456978 287688 456984 287700
rect 413336 287660 456984 287688
rect 413336 287648 413342 287660
rect 456978 287648 456984 287660
rect 457036 287648 457042 287700
rect 468478 287648 468484 287700
rect 468536 287688 468542 287700
rect 486418 287688 486424 287700
rect 468536 287660 486424 287688
rect 468536 287648 468542 287660
rect 486418 287648 486424 287660
rect 486476 287648 486482 287700
rect 121454 287580 121460 287632
rect 121512 287620 121518 287632
rect 122190 287620 122196 287632
rect 121512 287592 122196 287620
rect 121512 287580 121518 287592
rect 122190 287580 122196 287592
rect 122248 287580 122254 287632
rect 337378 287104 337384 287156
rect 337436 287144 337442 287156
rect 571610 287144 571616 287156
rect 337436 287116 571616 287144
rect 337436 287104 337442 287116
rect 571610 287104 571616 287116
rect 571668 287104 571674 287156
rect 59262 287036 59268 287088
rect 59320 287076 59326 287088
rect 67634 287076 67640 287088
rect 59320 287048 67640 287076
rect 59320 287036 59326 287048
rect 67634 287036 67640 287048
rect 67692 287036 67698 287088
rect 121546 287036 121552 287088
rect 121604 287076 121610 287088
rect 167730 287076 167736 287088
rect 121604 287048 167736 287076
rect 121604 287036 121610 287048
rect 167730 287036 167736 287048
rect 167788 287036 167794 287088
rect 342898 287036 342904 287088
rect 342956 287076 342962 287088
rect 583110 287076 583116 287088
rect 342956 287048 583116 287076
rect 342956 287036 342962 287048
rect 583110 287036 583116 287048
rect 583168 287036 583174 287088
rect 153102 286288 153108 286340
rect 153160 286328 153166 286340
rect 171778 286328 171784 286340
rect 153160 286300 171784 286328
rect 153160 286288 153166 286300
rect 171778 286288 171784 286300
rect 171836 286288 171842 286340
rect 363782 285812 363788 285864
rect 363840 285852 363846 285864
rect 514294 285852 514300 285864
rect 363840 285824 514300 285852
rect 363840 285812 363846 285824
rect 514294 285812 514300 285824
rect 514352 285812 514358 285864
rect 54938 285744 54944 285796
rect 54996 285784 55002 285796
rect 67726 285784 67732 285796
rect 54996 285756 67732 285784
rect 54996 285744 55002 285756
rect 67726 285744 67732 285756
rect 67784 285744 67790 285796
rect 121638 285744 121644 285796
rect 121696 285784 121702 285796
rect 153102 285784 153108 285796
rect 121696 285756 153108 285784
rect 121696 285744 121702 285756
rect 153102 285744 153108 285756
rect 153160 285744 153166 285796
rect 370590 285744 370596 285796
rect 370648 285784 370654 285796
rect 536834 285784 536840 285796
rect 370648 285756 536840 285784
rect 370648 285744 370654 285756
rect 536834 285744 536840 285756
rect 536892 285744 536898 285796
rect 41322 285676 41328 285728
rect 41380 285716 41386 285728
rect 67634 285716 67640 285728
rect 41380 285688 67640 285716
rect 41380 285676 41386 285688
rect 67634 285676 67640 285688
rect 67692 285676 67698 285728
rect 123662 285676 123668 285728
rect 123720 285716 123726 285728
rect 162762 285716 162768 285728
rect 123720 285688 162768 285716
rect 123720 285676 123726 285688
rect 162762 285676 162768 285688
rect 162820 285716 162826 285728
rect 176654 285716 176660 285728
rect 162820 285688 176660 285716
rect 162820 285676 162826 285688
rect 176654 285676 176660 285688
rect 176712 285676 176718 285728
rect 295334 285676 295340 285728
rect 295392 285716 295398 285728
rect 298922 285716 298928 285728
rect 295392 285688 298928 285716
rect 295392 285676 295398 285688
rect 298922 285676 298928 285688
rect 298980 285676 298986 285728
rect 381538 285676 381544 285728
rect 381596 285716 381602 285728
rect 582742 285716 582748 285728
rect 381596 285688 582748 285716
rect 381596 285676 381602 285688
rect 582742 285676 582748 285688
rect 582800 285716 582806 285728
rect 583294 285716 583300 285728
rect 582800 285688 583300 285716
rect 582800 285676 582806 285688
rect 583294 285676 583300 285688
rect 583352 285676 583358 285728
rect 121454 285608 121460 285660
rect 121512 285648 121518 285660
rect 175918 285648 175924 285660
rect 121512 285620 175924 285648
rect 121512 285608 121518 285620
rect 175918 285608 175924 285620
rect 175976 285608 175982 285660
rect 471238 284928 471244 284980
rect 471296 284968 471302 284980
rect 527174 284968 527180 284980
rect 471296 284940 527180 284968
rect 471296 284928 471302 284940
rect 527174 284928 527180 284940
rect 527232 284968 527238 284980
rect 530578 284968 530584 284980
rect 527232 284940 530584 284968
rect 527232 284928 527238 284940
rect 530578 284928 530584 284940
rect 530636 284928 530642 284980
rect 531958 284928 531964 284980
rect 532016 284968 532022 284980
rect 546494 284968 546500 284980
rect 532016 284940 546500 284968
rect 532016 284928 532022 284940
rect 546494 284928 546500 284940
rect 546552 284928 546558 284980
rect 387610 284588 387616 284640
rect 387668 284628 387674 284640
rect 392578 284628 392584 284640
rect 387668 284600 392584 284628
rect 387668 284588 387674 284600
rect 392578 284588 392584 284600
rect 392636 284588 392642 284640
rect 366358 284520 366364 284572
rect 366416 284560 366422 284572
rect 428642 284560 428648 284572
rect 366416 284532 428648 284560
rect 366416 284520 366422 284532
rect 428642 284520 428648 284532
rect 428700 284520 428706 284572
rect 365070 284452 365076 284504
rect 365128 284492 365134 284504
rect 473078 284492 473084 284504
rect 365128 284464 473084 284492
rect 365128 284452 365134 284464
rect 473078 284452 473084 284464
rect 473136 284452 473142 284504
rect 371878 284384 371884 284436
rect 371936 284424 371942 284436
rect 575474 284424 575480 284436
rect 371936 284396 575480 284424
rect 371936 284384 371942 284396
rect 575474 284384 575480 284396
rect 575532 284384 575538 284436
rect 57882 284316 57888 284368
rect 57940 284356 57946 284368
rect 67634 284356 67640 284368
rect 57940 284328 67640 284356
rect 57940 284316 57946 284328
rect 67634 284316 67640 284328
rect 67692 284316 67698 284368
rect 301498 284316 301504 284368
rect 301556 284356 301562 284368
rect 302050 284356 302056 284368
rect 301556 284328 302056 284356
rect 301556 284316 301562 284328
rect 302050 284316 302056 284328
rect 302108 284356 302114 284368
rect 583478 284356 583484 284368
rect 302108 284328 583484 284356
rect 302108 284316 302114 284328
rect 583478 284316 583484 284328
rect 583536 284316 583542 284368
rect 66162 284248 66168 284300
rect 66220 284288 66226 284300
rect 67818 284288 67824 284300
rect 66220 284260 67824 284288
rect 66220 284248 66226 284260
rect 67818 284248 67824 284260
rect 67876 284248 67882 284300
rect 574278 283772 574284 283824
rect 574336 283812 574342 283824
rect 574738 283812 574744 283824
rect 574336 283784 574744 283812
rect 574336 283772 574342 283784
rect 574738 283772 574744 283784
rect 574796 283772 574802 283824
rect 120810 283568 120816 283620
rect 120868 283608 120874 283620
rect 155862 283608 155868 283620
rect 120868 283580 155868 283608
rect 120868 283568 120874 283580
rect 155862 283568 155868 283580
rect 155920 283568 155926 283620
rect 389910 283228 389916 283280
rect 389968 283268 389974 283280
rect 441522 283268 441528 283280
rect 389968 283240 441528 283268
rect 389968 283228 389974 283240
rect 441522 283228 441528 283240
rect 441580 283228 441586 283280
rect 359642 283160 359648 283212
rect 359700 283200 359706 283212
rect 507854 283200 507860 283212
rect 359700 283172 507860 283200
rect 359700 283160 359706 283172
rect 507854 283160 507860 283172
rect 507912 283160 507918 283212
rect 371970 283092 371976 283144
rect 372028 283132 372034 283144
rect 574278 283132 574284 283144
rect 372028 283104 574284 283132
rect 372028 283092 372034 283104
rect 574278 283092 574284 283104
rect 574336 283092 574342 283144
rect 373350 283024 373356 283076
rect 373408 283064 373414 283076
rect 581178 283064 581184 283076
rect 373408 283036 581184 283064
rect 373408 283024 373414 283036
rect 581178 283024 581184 283036
rect 581236 283024 581242 283076
rect 341518 282956 341524 283008
rect 341576 282996 341582 283008
rect 555510 282996 555516 283008
rect 341576 282968 555516 282996
rect 341576 282956 341582 282968
rect 555510 282956 555516 282968
rect 555568 282956 555574 283008
rect 45370 282888 45376 282940
rect 45428 282928 45434 282940
rect 67726 282928 67732 282940
rect 45428 282900 67732 282928
rect 45428 282888 45434 282900
rect 67726 282888 67732 282900
rect 67784 282888 67790 282940
rect 121454 282888 121460 282940
rect 121512 282928 121518 282940
rect 142982 282928 142988 282940
rect 121512 282900 142988 282928
rect 121512 282888 121518 282900
rect 142982 282888 142988 282900
rect 143040 282888 143046 282940
rect 155862 282888 155868 282940
rect 155920 282928 155926 282940
rect 176654 282928 176660 282940
rect 155920 282900 176660 282928
rect 155920 282888 155926 282900
rect 176654 282888 176660 282900
rect 176712 282888 176718 282940
rect 295334 282888 295340 282940
rect 295392 282928 295398 282940
rect 569954 282928 569960 282940
rect 295392 282900 569960 282928
rect 295392 282888 295398 282900
rect 569954 282888 569960 282900
rect 570012 282928 570018 282940
rect 573542 282928 573548 282940
rect 570012 282900 573548 282928
rect 570012 282888 570018 282900
rect 573542 282888 573548 282900
rect 573600 282888 573606 282940
rect 64782 282820 64788 282872
rect 64840 282860 64846 282872
rect 67634 282860 67640 282872
rect 64840 282832 67640 282860
rect 64840 282820 64846 282832
rect 67634 282820 67640 282832
rect 67692 282820 67698 282872
rect 120994 282140 121000 282192
rect 121052 282180 121058 282192
rect 158714 282180 158720 282192
rect 121052 282152 158720 282180
rect 121052 282140 121058 282152
rect 158714 282140 158720 282152
rect 158772 282140 158778 282192
rect 374822 281868 374828 281920
rect 374880 281908 374886 281920
rect 438302 281908 438308 281920
rect 374880 281880 438308 281908
rect 374880 281868 374886 281880
rect 438302 281868 438308 281880
rect 438360 281868 438366 281920
rect 374730 281800 374736 281852
rect 374788 281840 374794 281852
rect 482738 281840 482744 281852
rect 374788 281812 482744 281840
rect 374788 281800 374794 281812
rect 482738 281800 482744 281812
rect 482796 281800 482802 281852
rect 369210 281732 369216 281784
rect 369268 281772 369274 281784
rect 523954 281772 523960 281784
rect 369268 281744 523960 281772
rect 369268 281732 369274 281744
rect 523954 281732 523960 281744
rect 524012 281732 524018 281784
rect 377490 281664 377496 281716
rect 377548 281704 377554 281716
rect 567838 281704 567844 281716
rect 377548 281676 567844 281704
rect 377548 281664 377554 281676
rect 567838 281664 567844 281676
rect 567896 281704 567902 281716
rect 568390 281704 568396 281716
rect 567896 281676 568396 281704
rect 567896 281664 567902 281676
rect 568390 281664 568396 281676
rect 568448 281664 568454 281716
rect 384206 281596 384212 281648
rect 384264 281636 384270 281648
rect 576946 281636 576952 281648
rect 384264 281608 576952 281636
rect 384264 281596 384270 281608
rect 576946 281596 576952 281608
rect 577004 281636 577010 281648
rect 577498 281636 577504 281648
rect 577004 281608 577504 281636
rect 577004 281596 577010 281608
rect 577498 281596 577504 281608
rect 577556 281596 577562 281648
rect 121454 281528 121460 281580
rect 121512 281568 121518 281580
rect 157978 281568 157984 281580
rect 121512 281540 157984 281568
rect 121512 281528 121518 281540
rect 157978 281528 157984 281540
rect 158036 281528 158042 281580
rect 158714 281528 158720 281580
rect 158772 281568 158778 281580
rect 159910 281568 159916 281580
rect 158772 281540 159916 281568
rect 158772 281528 158778 281540
rect 159910 281528 159916 281540
rect 159968 281568 159974 281580
rect 176654 281568 176660 281580
rect 159968 281540 176660 281568
rect 159968 281528 159974 281540
rect 176654 281528 176660 281540
rect 176712 281528 176718 281580
rect 295334 281528 295340 281580
rect 295392 281568 295398 281580
rect 295518 281568 295524 281580
rect 295392 281540 295524 281568
rect 295392 281528 295398 281540
rect 295518 281528 295524 281540
rect 295576 281568 295582 281580
rect 356698 281568 356704 281580
rect 295576 281540 356704 281568
rect 295576 281528 295582 281540
rect 356698 281528 356704 281540
rect 356756 281528 356762 281580
rect 362310 281528 362316 281580
rect 362368 281568 362374 281580
rect 582466 281568 582472 281580
rect 362368 281540 582472 281568
rect 362368 281528 362374 281540
rect 582466 281528 582472 281540
rect 582524 281528 582530 281580
rect 157150 281460 157156 281512
rect 157208 281500 157214 281512
rect 157334 281500 157340 281512
rect 157208 281472 157340 281500
rect 157208 281460 157214 281472
rect 157334 281460 157340 281472
rect 157392 281460 157398 281512
rect 121546 280780 121552 280832
rect 121604 280820 121610 280832
rect 167822 280820 167828 280832
rect 121604 280792 167828 280820
rect 121604 280780 121610 280792
rect 167822 280780 167828 280792
rect 167880 280780 167886 280832
rect 169110 280780 169116 280832
rect 169168 280820 169174 280832
rect 175274 280820 175280 280832
rect 169168 280792 175280 280820
rect 169168 280780 169174 280792
rect 175274 280780 175280 280792
rect 175332 280780 175338 280832
rect 377674 280508 377680 280560
rect 377732 280548 377738 280560
rect 397086 280548 397092 280560
rect 377732 280520 397092 280548
rect 377732 280508 377738 280520
rect 397086 280508 397092 280520
rect 397144 280508 397150 280560
rect 367922 280440 367928 280492
rect 367980 280480 367986 280492
rect 409230 280480 409236 280492
rect 367980 280452 409236 280480
rect 367980 280440 367986 280452
rect 409230 280440 409236 280452
rect 409288 280440 409294 280492
rect 376018 280372 376024 280424
rect 376076 280412 376082 280424
rect 469858 280412 469864 280424
rect 376076 280384 469864 280412
rect 376076 280372 376082 280384
rect 469858 280372 469864 280384
rect 469916 280372 469922 280424
rect 297542 280304 297548 280356
rect 297600 280344 297606 280356
rect 425422 280344 425428 280356
rect 297600 280316 425428 280344
rect 297600 280304 297606 280316
rect 425422 280304 425428 280316
rect 425480 280344 425486 280356
rect 573450 280344 573456 280356
rect 425480 280316 573456 280344
rect 425480 280304 425486 280316
rect 573450 280304 573456 280316
rect 573508 280304 573514 280356
rect 389634 280236 389640 280288
rect 389692 280276 389698 280288
rect 574186 280276 574192 280288
rect 389692 280248 574192 280276
rect 389692 280236 389698 280248
rect 574186 280236 574192 280248
rect 574244 280236 574250 280288
rect 53742 280168 53748 280220
rect 53800 280208 53806 280220
rect 67634 280208 67640 280220
rect 53800 280180 67640 280208
rect 53800 280168 53806 280180
rect 67634 280168 67640 280180
rect 67692 280168 67698 280220
rect 121454 280168 121460 280220
rect 121512 280208 121518 280220
rect 138934 280208 138940 280220
rect 121512 280180 138940 280208
rect 121512 280168 121518 280180
rect 138934 280168 138940 280180
rect 138992 280168 138998 280220
rect 157150 280168 157156 280220
rect 157208 280208 157214 280220
rect 157208 280180 158668 280208
rect 157208 280168 157214 280180
rect 158640 280140 158668 280180
rect 326338 280168 326344 280220
rect 326396 280208 326402 280220
rect 581086 280208 581092 280220
rect 326396 280180 581092 280208
rect 326396 280168 326402 280180
rect 581086 280168 581092 280180
rect 581144 280168 581150 280220
rect 176654 280140 176660 280152
rect 158640 280112 176660 280140
rect 176654 280100 176660 280112
rect 176712 280100 176718 280152
rect 378870 279080 378876 279132
rect 378928 279120 378934 279132
rect 393866 279120 393872 279132
rect 378928 279092 393872 279120
rect 378928 279080 378934 279092
rect 393866 279080 393872 279092
rect 393924 279080 393930 279132
rect 381630 279012 381636 279064
rect 381688 279052 381694 279064
rect 403526 279052 403532 279064
rect 381688 279024 403532 279052
rect 381688 279012 381694 279024
rect 403526 279012 403532 279024
rect 403584 279012 403590 279064
rect 300210 278944 300216 278996
rect 300268 278984 300274 278996
rect 447962 278984 447968 278996
rect 300268 278956 447968 278984
rect 300268 278944 300274 278956
rect 447962 278944 447968 278956
rect 448020 278984 448026 278996
rect 583754 278984 583760 278996
rect 448020 278956 583760 278984
rect 448020 278944 448026 278956
rect 583754 278944 583760 278956
rect 583812 278944 583818 278996
rect 373258 278876 373264 278928
rect 373316 278916 373322 278928
rect 400306 278916 400312 278928
rect 373316 278888 400312 278916
rect 373316 278876 373322 278888
rect 400306 278876 400312 278888
rect 400364 278876 400370 278928
rect 421558 278876 421564 278928
rect 421616 278916 421622 278928
rect 421834 278916 421840 278928
rect 421616 278888 421840 278916
rect 421616 278876 421622 278888
rect 421834 278876 421840 278888
rect 421892 278916 421898 278928
rect 581638 278916 581644 278928
rect 421892 278888 581644 278916
rect 421892 278876 421898 278888
rect 581638 278876 581644 278888
rect 581696 278876 581702 278928
rect 121454 278808 121460 278860
rect 121512 278848 121518 278860
rect 151078 278848 151084 278860
rect 121512 278820 151084 278848
rect 121512 278808 121518 278820
rect 151078 278808 151084 278820
rect 151136 278808 151142 278860
rect 158530 278808 158536 278860
rect 158588 278848 158594 278860
rect 171134 278848 171140 278860
rect 158588 278820 171140 278848
rect 158588 278808 158594 278820
rect 171134 278808 171140 278820
rect 171192 278848 171198 278860
rect 171192 278820 172468 278848
rect 171192 278808 171198 278820
rect 35802 278740 35808 278792
rect 35860 278780 35866 278792
rect 67634 278780 67640 278792
rect 35860 278752 67640 278780
rect 35860 278740 35866 278752
rect 67634 278740 67640 278752
rect 67692 278740 67698 278792
rect 121546 278740 121552 278792
rect 121604 278780 121610 278792
rect 171778 278780 171784 278792
rect 121604 278752 171784 278780
rect 121604 278740 121610 278752
rect 171778 278740 171784 278752
rect 171836 278740 171842 278792
rect 172440 278712 172468 278820
rect 295334 278808 295340 278860
rect 295392 278848 295398 278860
rect 298830 278848 298836 278860
rect 295392 278820 298836 278848
rect 295392 278808 295398 278820
rect 298830 278808 298836 278820
rect 298888 278808 298894 278860
rect 391934 278808 391940 278860
rect 391992 278848 391998 278860
rect 580442 278848 580448 278860
rect 391992 278820 580448 278848
rect 391992 278808 391998 278820
rect 580442 278808 580448 278820
rect 580500 278808 580506 278860
rect 379422 278740 379428 278792
rect 379480 278780 379486 278792
rect 583386 278780 583392 278792
rect 379480 278752 583392 278780
rect 379480 278740 379486 278752
rect 583386 278740 583392 278752
rect 583444 278740 583450 278792
rect 176654 278712 176660 278724
rect 172440 278684 176660 278712
rect 176654 278672 176660 278684
rect 176712 278672 176718 278724
rect 501414 278672 501420 278724
rect 501472 278712 501478 278724
rect 502334 278712 502340 278724
rect 501472 278684 502340 278712
rect 501472 278672 501478 278684
rect 502334 278672 502340 278684
rect 502392 278672 502398 278724
rect 538858 278672 538864 278724
rect 538916 278712 538922 278724
rect 543274 278712 543280 278724
rect 538916 278684 543280 278712
rect 538916 278672 538922 278684
rect 543274 278672 543280 278684
rect 543332 278672 543338 278724
rect 563698 278672 563704 278724
rect 563756 278712 563762 278724
rect 565170 278712 565176 278724
rect 563756 278684 565176 278712
rect 563756 278672 563762 278684
rect 565170 278672 565176 278684
rect 565228 278672 565234 278724
rect 577590 278672 577596 278724
rect 577648 278712 577654 278724
rect 580258 278712 580264 278724
rect 577648 278684 580264 278712
rect 577648 278672 577654 278684
rect 580258 278672 580264 278684
rect 580316 278672 580322 278724
rect 352558 278060 352564 278112
rect 352616 278100 352622 278112
rect 384206 278100 384212 278112
rect 352616 278072 384212 278100
rect 352616 278060 352622 278072
rect 384206 278060 384212 278072
rect 384264 278060 384270 278112
rect 314010 277992 314016 278044
rect 314068 278032 314074 278044
rect 385862 278032 385868 278044
rect 314068 278004 385868 278032
rect 314068 277992 314074 278004
rect 385862 277992 385868 278004
rect 385920 277992 385926 278044
rect 65978 277788 65984 277840
rect 66036 277828 66042 277840
rect 68094 277828 68100 277840
rect 66036 277800 68100 277828
rect 66036 277788 66042 277800
rect 68094 277788 68100 277800
rect 68152 277788 68158 277840
rect 389818 277720 389824 277772
rect 389876 277760 389882 277772
rect 549070 277760 549076 277772
rect 389876 277732 549076 277760
rect 389876 277720 389882 277732
rect 549070 277720 549076 277732
rect 549128 277720 549134 277772
rect 364978 277652 364984 277704
rect 365036 277692 365042 277704
rect 431862 277692 431868 277704
rect 365036 277664 431868 277692
rect 365036 277652 365042 277664
rect 431862 277652 431868 277664
rect 431920 277652 431926 277704
rect 452654 277652 452660 277704
rect 452712 277692 452718 277704
rect 489178 277692 489184 277704
rect 452712 277664 489184 277692
rect 452712 277652 452718 277664
rect 489178 277652 489184 277664
rect 489236 277652 489242 277704
rect 385678 277584 385684 277636
rect 385736 277624 385742 277636
rect 453758 277624 453764 277636
rect 385736 277596 453764 277624
rect 385736 277584 385742 277596
rect 453758 277584 453764 277596
rect 453816 277584 453822 277636
rect 486418 277584 486424 277636
rect 486476 277624 486482 277636
rect 576210 277624 576216 277636
rect 486476 277596 576216 277624
rect 486476 277584 486482 277596
rect 576210 277584 576216 277596
rect 576268 277584 576274 277636
rect 380158 277516 380164 277568
rect 380216 277556 380222 277568
rect 495618 277556 495624 277568
rect 380216 277528 495624 277556
rect 380216 277516 380222 277528
rect 495618 277516 495624 277528
rect 495676 277516 495682 277568
rect 121546 277448 121552 277500
rect 121604 277488 121610 277500
rect 133322 277488 133328 277500
rect 121604 277460 133328 277488
rect 121604 277448 121610 277460
rect 133322 277448 133328 277460
rect 133380 277448 133386 277500
rect 385770 277448 385776 277500
rect 385828 277488 385834 277500
rect 517514 277488 517520 277500
rect 385828 277460 517520 277488
rect 385828 277448 385834 277460
rect 517514 277448 517520 277460
rect 517572 277448 517578 277500
rect 63402 277380 63408 277432
rect 63460 277420 63466 277432
rect 67634 277420 67640 277432
rect 63460 277392 67640 277420
rect 63460 277380 63466 277392
rect 67634 277380 67640 277392
rect 67692 277380 67698 277432
rect 121454 277380 121460 277432
rect 121512 277420 121518 277432
rect 163498 277420 163504 277432
rect 121512 277392 163504 277420
rect 121512 277380 121518 277392
rect 163498 277380 163504 277392
rect 163556 277380 163562 277432
rect 566458 277040 566464 277092
rect 566516 277080 566522 277092
rect 568666 277080 568672 277092
rect 566516 277052 568672 277080
rect 566516 277040 566522 277052
rect 568666 277040 568672 277052
rect 568724 277040 568730 277092
rect 301314 276632 301320 276684
rect 301372 276672 301378 276684
rect 381538 276672 381544 276684
rect 301372 276644 381544 276672
rect 301372 276632 301378 276644
rect 381538 276632 381544 276644
rect 381596 276632 381602 276684
rect 382182 276632 382188 276684
rect 382240 276672 382246 276684
rect 391934 276672 391940 276684
rect 382240 276644 391940 276672
rect 382240 276632 382246 276644
rect 391934 276632 391940 276644
rect 391992 276632 391998 276684
rect 566550 276632 566556 276684
rect 566608 276672 566614 276684
rect 571518 276672 571524 276684
rect 566608 276644 571524 276672
rect 566608 276632 566614 276644
rect 571518 276632 571524 276644
rect 571576 276632 571582 276684
rect 410334 276360 410340 276412
rect 410392 276400 410398 276412
rect 582650 276400 582656 276412
rect 410392 276372 582656 276400
rect 410392 276360 410398 276372
rect 582650 276360 582656 276372
rect 582708 276360 582714 276412
rect 385862 276292 385868 276344
rect 385920 276332 385926 276344
rect 466638 276332 466644 276344
rect 385920 276304 466644 276332
rect 385920 276292 385926 276304
rect 466638 276292 466644 276304
rect 466696 276292 466702 276344
rect 382918 276224 382924 276276
rect 382976 276264 382982 276276
rect 530394 276264 530400 276276
rect 382976 276236 530400 276264
rect 382976 276224 382982 276236
rect 530394 276224 530400 276236
rect 530452 276224 530458 276276
rect 367830 276156 367836 276208
rect 367888 276196 367894 276208
rect 412542 276196 412548 276208
rect 367888 276168 412548 276196
rect 367888 276156 367894 276168
rect 412542 276156 412548 276168
rect 412600 276156 412606 276208
rect 52270 276088 52276 276140
rect 52328 276128 52334 276140
rect 67726 276128 67732 276140
rect 52328 276100 67732 276128
rect 52328 276088 52334 276100
rect 67726 276088 67732 276100
rect 67784 276088 67790 276140
rect 121546 276088 121552 276140
rect 121604 276128 121610 276140
rect 147214 276128 147220 276140
rect 121604 276100 147220 276128
rect 121604 276088 121610 276100
rect 147214 276088 147220 276100
rect 147272 276088 147278 276140
rect 383010 276088 383016 276140
rect 383068 276128 383074 276140
rect 570138 276128 570144 276140
rect 383068 276100 570144 276128
rect 383068 276088 383074 276100
rect 570138 276088 570144 276100
rect 570196 276088 570202 276140
rect 48222 276020 48228 276072
rect 48280 276060 48286 276072
rect 67634 276060 67640 276072
rect 48280 276032 67640 276060
rect 48280 276020 48286 276032
rect 67634 276020 67640 276032
rect 67692 276020 67698 276072
rect 121454 276020 121460 276072
rect 121512 276060 121518 276072
rect 170582 276060 170588 276072
rect 121512 276032 170588 276060
rect 121512 276020 121518 276032
rect 170582 276020 170588 276032
rect 170640 276020 170646 276072
rect 172330 276020 172336 276072
rect 172388 276060 172394 276072
rect 175274 276060 175280 276072
rect 172388 276032 175280 276060
rect 172388 276020 172394 276032
rect 175274 276020 175280 276032
rect 175332 276020 175338 276072
rect 295334 276020 295340 276072
rect 295392 276060 295398 276072
rect 300946 276060 300952 276072
rect 295392 276032 300952 276060
rect 295392 276020 295398 276032
rect 300946 276020 300952 276032
rect 301004 276060 301010 276072
rect 301314 276060 301320 276072
rect 301004 276032 301320 276060
rect 301004 276020 301010 276032
rect 301314 276020 301320 276032
rect 301372 276020 301378 276072
rect 353938 276020 353944 276072
rect 353996 276060 354002 276072
rect 354582 276060 354588 276072
rect 353996 276032 354588 276060
rect 353996 276020 354002 276032
rect 354582 276020 354588 276032
rect 354640 276060 354646 276072
rect 571334 276060 571340 276072
rect 354640 276032 571340 276060
rect 354640 276020 354646 276032
rect 571334 276020 571340 276032
rect 571392 276020 571398 276072
rect 175292 275992 175320 276020
rect 177482 275992 177488 276004
rect 175292 275964 177488 275992
rect 177482 275952 177488 275964
rect 177540 275952 177546 276004
rect 363598 275952 363604 276004
rect 363656 275992 363662 276004
rect 364242 275992 364248 276004
rect 363656 275964 364248 275992
rect 363656 275952 363662 275964
rect 364242 275952 364248 275964
rect 364300 275992 364306 276004
rect 410334 275992 410340 276004
rect 364300 275964 410340 275992
rect 364300 275952 364306 275964
rect 410334 275952 410340 275964
rect 410392 275952 410398 276004
rect 405706 275624 415394 275652
rect 295978 275340 295984 275392
rect 296036 275380 296042 275392
rect 405706 275380 405734 275624
rect 409690 275544 409696 275596
rect 409748 275584 409754 275596
rect 409748 275556 411484 275584
rect 409748 275544 409754 275556
rect 296036 275352 405734 275380
rect 296036 275340 296042 275352
rect 370498 275272 370504 275324
rect 370556 275312 370562 275324
rect 389634 275312 389640 275324
rect 370556 275284 389640 275312
rect 370556 275272 370562 275284
rect 389634 275272 389640 275284
rect 389692 275272 389698 275324
rect 411456 275312 411484 275556
rect 415366 275448 415394 275624
rect 452654 275584 452660 275596
rect 431926 275556 452660 275584
rect 415366 275420 418154 275448
rect 418126 275380 418154 275420
rect 431926 275380 431954 275556
rect 452654 275544 452660 275556
rect 452712 275544 452718 275596
rect 418126 275352 431954 275380
rect 580166 275312 580172 275324
rect 411456 275284 580172 275312
rect 580166 275272 580172 275284
rect 580224 275272 580230 275324
rect 389726 275204 389732 275256
rect 389784 275244 389790 275256
rect 389910 275244 389916 275256
rect 389784 275216 389916 275244
rect 389784 275204 389790 275216
rect 389910 275204 389916 275216
rect 389968 275204 389974 275256
rect 64690 274728 64696 274780
rect 64748 274768 64754 274780
rect 67634 274768 67640 274780
rect 64748 274740 67640 274768
rect 64748 274728 64754 274740
rect 67634 274728 67640 274740
rect 67692 274728 67698 274780
rect 121454 274728 121460 274780
rect 121512 274768 121518 274780
rect 126238 274768 126244 274780
rect 121512 274740 126244 274768
rect 121512 274728 121518 274740
rect 126238 274728 126244 274740
rect 126296 274728 126302 274780
rect 121546 274660 121552 274712
rect 121604 274700 121610 274712
rect 145742 274700 145748 274712
rect 121604 274672 145748 274700
rect 121604 274660 121610 274672
rect 145742 274660 145748 274672
rect 145800 274660 145806 274712
rect 295334 274660 295340 274712
rect 295392 274700 295398 274712
rect 298738 274700 298744 274712
rect 295392 274672 298744 274700
rect 295392 274660 295398 274672
rect 298738 274660 298744 274672
rect 298796 274700 298802 274712
rect 298796 274672 299428 274700
rect 298796 274660 298802 274672
rect 121454 274592 121460 274644
rect 121512 274632 121518 274644
rect 166258 274632 166264 274644
rect 121512 274604 166264 274632
rect 121512 274592 121518 274604
rect 166258 274592 166264 274604
rect 166316 274592 166322 274644
rect 299400 274632 299428 274672
rect 385034 274632 385040 274644
rect 299400 274604 385040 274632
rect 385034 274592 385040 274604
rect 385092 274592 385098 274644
rect 22738 273912 22744 273964
rect 22796 273952 22802 273964
rect 60090 273952 60096 273964
rect 22796 273924 60096 273952
rect 22796 273912 22802 273924
rect 60090 273912 60096 273924
rect 60148 273912 60154 273964
rect 61930 273300 61936 273352
rect 61988 273340 61994 273352
rect 67634 273340 67640 273352
rect 61988 273312 67640 273340
rect 61988 273300 61994 273312
rect 67634 273300 67640 273312
rect 67692 273300 67698 273352
rect 60090 273232 60096 273284
rect 60148 273272 60154 273284
rect 60366 273272 60372 273284
rect 60148 273244 60372 273272
rect 60148 273232 60154 273244
rect 60366 273232 60372 273244
rect 60424 273272 60430 273284
rect 67726 273272 67732 273284
rect 60424 273244 67732 273272
rect 60424 273232 60430 273244
rect 67726 273232 67732 273244
rect 67784 273232 67790 273284
rect 121454 273232 121460 273284
rect 121512 273272 121518 273284
rect 141418 273272 141424 273284
rect 121512 273244 141424 273272
rect 121512 273232 121518 273244
rect 141418 273232 141424 273244
rect 141476 273232 141482 273284
rect 345750 273232 345756 273284
rect 345808 273272 345814 273284
rect 386874 273272 386880 273284
rect 345808 273244 386880 273272
rect 345808 273232 345814 273244
rect 386874 273232 386880 273244
rect 386932 273232 386938 273284
rect 120994 272484 121000 272536
rect 121052 272524 121058 272536
rect 124214 272524 124220 272536
rect 121052 272496 124220 272524
rect 121052 272484 121058 272496
rect 124214 272484 124220 272496
rect 124272 272524 124278 272536
rect 160094 272524 160100 272536
rect 124272 272496 160100 272524
rect 124272 272484 124278 272496
rect 160094 272484 160100 272496
rect 160152 272484 160158 272536
rect 121454 272008 121460 272060
rect 121512 272048 121518 272060
rect 125042 272048 125048 272060
rect 121512 272020 125048 272048
rect 121512 272008 121518 272020
rect 125042 272008 125048 272020
rect 125100 272008 125106 272060
rect 64782 271872 64788 271924
rect 64840 271912 64846 271924
rect 67634 271912 67640 271924
rect 64840 271884 67640 271912
rect 64840 271872 64846 271884
rect 67634 271872 67640 271884
rect 67692 271872 67698 271924
rect 160094 271872 160100 271924
rect 160152 271912 160158 271924
rect 161198 271912 161204 271924
rect 160152 271884 161204 271912
rect 160152 271872 160158 271884
rect 161198 271872 161204 271884
rect 161256 271912 161262 271924
rect 176654 271912 176660 271924
rect 161256 271884 176660 271912
rect 161256 271872 161262 271884
rect 176654 271872 176660 271884
rect 176712 271872 176718 271924
rect 295334 271872 295340 271924
rect 295392 271912 295398 271924
rect 306466 271912 306472 271924
rect 295392 271884 306472 271912
rect 295392 271872 295398 271884
rect 306466 271872 306472 271884
rect 306524 271912 306530 271924
rect 381538 271912 381544 271924
rect 306524 271884 381544 271912
rect 306524 271872 306530 271884
rect 381538 271872 381544 271884
rect 381596 271872 381602 271924
rect 64598 271804 64604 271856
rect 64656 271844 64662 271856
rect 67726 271844 67732 271856
rect 64656 271816 67732 271844
rect 64656 271804 64662 271816
rect 67726 271804 67732 271816
rect 67784 271804 67790 271856
rect 325050 271124 325056 271176
rect 325108 271164 325114 271176
rect 350534 271164 350540 271176
rect 325108 271136 350540 271164
rect 325108 271124 325114 271136
rect 350534 271124 350540 271136
rect 350592 271124 350598 271176
rect 46842 270512 46848 270564
rect 46900 270552 46906 270564
rect 67634 270552 67640 270564
rect 46900 270524 67640 270552
rect 46900 270512 46906 270524
rect 67634 270512 67640 270524
rect 67692 270512 67698 270564
rect 121454 270512 121460 270564
rect 121512 270552 121518 270564
rect 130654 270552 130660 270564
rect 121512 270524 130660 270552
rect 121512 270512 121518 270524
rect 130654 270512 130660 270524
rect 130712 270512 130718 270564
rect 140682 269764 140688 269816
rect 140740 269804 140746 269816
rect 169018 269804 169024 269816
rect 140740 269776 169024 269804
rect 140740 269764 140746 269776
rect 169018 269764 169024 269776
rect 169076 269764 169082 269816
rect 366450 269764 366456 269816
rect 366508 269804 366514 269816
rect 387150 269804 387156 269816
rect 366508 269776 387156 269804
rect 366508 269764 366514 269776
rect 387150 269764 387156 269776
rect 387208 269764 387214 269816
rect 121546 269152 121552 269204
rect 121604 269192 121610 269204
rect 125134 269192 125140 269204
rect 121604 269164 125140 269192
rect 121604 269152 121610 269164
rect 125134 269152 125140 269164
rect 125192 269152 125198 269204
rect 49510 269084 49516 269136
rect 49568 269124 49574 269136
rect 67634 269124 67640 269136
rect 49568 269096 67640 269124
rect 49568 269084 49574 269096
rect 67634 269084 67640 269096
rect 67692 269084 67698 269136
rect 121454 269084 121460 269136
rect 121512 269124 121518 269136
rect 143074 269124 143080 269136
rect 121512 269096 143080 269124
rect 121512 269084 121518 269096
rect 143074 269084 143080 269096
rect 143132 269084 143138 269136
rect 295334 269084 295340 269136
rect 295392 269124 295398 269136
rect 325050 269124 325056 269136
rect 295392 269096 325056 269124
rect 295392 269084 295398 269096
rect 325050 269084 325056 269096
rect 325108 269084 325114 269136
rect 66162 268200 66168 268252
rect 66220 268240 66226 268252
rect 68186 268240 68192 268252
rect 66220 268212 68192 268240
rect 66220 268200 66226 268212
rect 68186 268200 68192 268212
rect 68244 268200 68250 268252
rect 13078 267724 13084 267776
rect 13136 267764 13142 267776
rect 57606 267764 57612 267776
rect 13136 267736 57612 267764
rect 13136 267724 13142 267736
rect 57606 267724 57612 267736
rect 57664 267764 57670 267776
rect 67634 267764 67640 267776
rect 57664 267736 67640 267764
rect 57664 267724 57670 267736
rect 67634 267724 67640 267736
rect 67692 267724 67698 267776
rect 161382 267724 161388 267776
rect 161440 267764 161446 267776
rect 176654 267764 176660 267776
rect 161440 267736 176660 267764
rect 161440 267724 161446 267736
rect 176654 267724 176660 267736
rect 176712 267724 176718 267776
rect 57238 267656 57244 267708
rect 57296 267696 57302 267708
rect 68922 267696 68928 267708
rect 57296 267668 68928 267696
rect 57296 267656 57302 267668
rect 68922 267656 68928 267668
rect 68980 267656 68986 267708
rect 62758 267044 62764 267096
rect 62816 267084 62822 267096
rect 63310 267084 63316 267096
rect 62816 267056 63316 267084
rect 62816 267044 62822 267056
rect 63310 267044 63316 267056
rect 63368 267084 63374 267096
rect 67634 267084 67640 267096
rect 63368 267056 67640 267084
rect 63368 267044 63374 267056
rect 67634 267044 67640 267056
rect 67692 267044 67698 267096
rect 298922 267044 298928 267096
rect 298980 267084 298986 267096
rect 328454 267084 328460 267096
rect 298980 267056 328460 267084
rect 298980 267044 298986 267056
rect 328454 267044 328460 267056
rect 328512 267044 328518 267096
rect 306282 266976 306288 267028
rect 306340 267016 306346 267028
rect 389726 267016 389732 267028
rect 306340 266988 389732 267016
rect 306340 266976 306346 266988
rect 389726 266976 389732 266988
rect 389784 266976 389790 267028
rect 3050 266364 3056 266416
rect 3108 266404 3114 266416
rect 25498 266404 25504 266416
rect 3108 266376 25504 266404
rect 3108 266364 3114 266376
rect 25498 266364 25504 266376
rect 25556 266364 25562 266416
rect 121454 266364 121460 266416
rect 121512 266404 121518 266416
rect 166442 266404 166448 266416
rect 121512 266376 166448 266404
rect 121512 266364 121518 266376
rect 166442 266364 166448 266376
rect 166500 266364 166506 266416
rect 165614 266296 165620 266348
rect 165672 266336 165678 266348
rect 176654 266336 176660 266348
rect 165672 266308 176660 266336
rect 165672 266296 165678 266308
rect 176654 266296 176660 266308
rect 176712 266296 176718 266348
rect 45462 265616 45468 265668
rect 45520 265656 45526 265668
rect 60734 265656 60740 265668
rect 45520 265628 60740 265656
rect 45520 265616 45526 265628
rect 60734 265616 60740 265628
rect 60792 265616 60798 265668
rect 60734 265004 60740 265056
rect 60792 265044 60798 265056
rect 61838 265044 61844 265056
rect 60792 265016 61844 265044
rect 60792 265004 60798 265016
rect 61838 265004 61844 265016
rect 61896 265044 61902 265056
rect 67634 265044 67640 265056
rect 61896 265016 67640 265044
rect 61896 265004 61902 265016
rect 67634 265004 67640 265016
rect 67692 265004 67698 265056
rect 48130 264936 48136 264988
rect 48188 264976 48194 264988
rect 67726 264976 67732 264988
rect 48188 264948 67732 264976
rect 48188 264936 48194 264948
rect 67726 264936 67732 264948
rect 67784 264936 67790 264988
rect 121454 264936 121460 264988
rect 121512 264976 121518 264988
rect 166258 264976 166264 264988
rect 121512 264948 166264 264976
rect 121512 264936 121518 264948
rect 166258 264936 166264 264948
rect 166316 264936 166322 264988
rect 59170 264188 59176 264240
rect 59228 264228 59234 264240
rect 67634 264228 67640 264240
rect 59228 264200 67640 264228
rect 59228 264188 59234 264200
rect 67634 264188 67640 264200
rect 67692 264188 67698 264240
rect 295334 264188 295340 264240
rect 295392 264228 295398 264240
rect 331858 264228 331864 264240
rect 295392 264200 331864 264228
rect 295392 264188 295398 264200
rect 331858 264188 331864 264200
rect 331916 264188 331922 264240
rect 50890 263644 50896 263696
rect 50948 263684 50954 263696
rect 67634 263684 67640 263696
rect 50948 263656 67640 263684
rect 50948 263644 50954 263656
rect 67634 263644 67640 263656
rect 67692 263644 67698 263696
rect 121454 263644 121460 263696
rect 121512 263684 121518 263696
rect 136174 263684 136180 263696
rect 121512 263656 136180 263684
rect 121512 263644 121518 263656
rect 136174 263644 136180 263656
rect 136232 263644 136238 263696
rect 21358 263576 21364 263628
rect 21416 263616 21422 263628
rect 59170 263616 59176 263628
rect 21416 263588 59176 263616
rect 21416 263576 21422 263588
rect 59170 263576 59176 263588
rect 59228 263576 59234 263628
rect 121546 263576 121552 263628
rect 121604 263616 121610 263628
rect 163590 263616 163596 263628
rect 121604 263588 163596 263616
rect 121604 263576 121610 263588
rect 163590 263576 163596 263588
rect 163648 263576 163654 263628
rect 121454 263508 121460 263560
rect 121512 263548 121518 263560
rect 146938 263548 146944 263560
rect 121512 263520 146944 263548
rect 121512 263508 121518 263520
rect 146938 263508 146944 263520
rect 146996 263508 147002 263560
rect 140222 262964 140228 263016
rect 140280 263004 140286 263016
rect 162302 263004 162308 263016
rect 140280 262976 162308 263004
rect 140280 262964 140286 262976
rect 162302 262964 162308 262976
rect 162360 262964 162366 263016
rect 146938 262896 146944 262948
rect 146996 262936 147002 262948
rect 169110 262936 169116 262948
rect 146996 262908 169116 262936
rect 146996 262896 147002 262908
rect 169110 262896 169116 262908
rect 169168 262896 169174 262948
rect 36538 262828 36544 262880
rect 36596 262868 36602 262880
rect 57790 262868 57796 262880
rect 36596 262840 57796 262868
rect 36596 262828 36602 262840
rect 57790 262828 57796 262840
rect 57848 262828 57854 262880
rect 122190 262828 122196 262880
rect 122248 262868 122254 262880
rect 169018 262868 169024 262880
rect 122248 262840 169024 262868
rect 122248 262828 122254 262840
rect 169018 262828 169024 262840
rect 169076 262828 169082 262880
rect 57790 262284 57796 262336
rect 57848 262324 57854 262336
rect 67726 262324 67732 262336
rect 57848 262296 67732 262324
rect 57848 262284 57854 262296
rect 67726 262284 67732 262296
rect 67784 262284 67790 262336
rect 56502 262216 56508 262268
rect 56560 262256 56566 262268
rect 67634 262256 67640 262268
rect 56560 262228 67640 262256
rect 56560 262216 56566 262228
rect 67634 262216 67640 262228
rect 67692 262216 67698 262268
rect 121454 262216 121460 262268
rect 121512 262256 121518 262268
rect 141602 262256 141608 262268
rect 121512 262228 141608 262256
rect 121512 262216 121518 262228
rect 141602 262216 141608 262228
rect 141660 262216 141666 262268
rect 331950 262216 331956 262268
rect 332008 262256 332014 262268
rect 386874 262256 386880 262268
rect 332008 262228 386880 262256
rect 332008 262216 332014 262228
rect 386874 262216 386880 262228
rect 386932 262216 386938 262268
rect 121454 261468 121460 261520
rect 121512 261508 121518 261520
rect 143534 261508 143540 261520
rect 121512 261480 143540 261508
rect 121512 261468 121518 261480
rect 143534 261468 143540 261480
rect 143592 261508 143598 261520
rect 144454 261508 144460 261520
rect 143592 261480 144460 261508
rect 143592 261468 143598 261480
rect 144454 261468 144460 261480
rect 144512 261468 144518 261520
rect 162302 261468 162308 261520
rect 162360 261508 162366 261520
rect 162670 261508 162676 261520
rect 162360 261480 162676 261508
rect 162360 261468 162366 261480
rect 162670 261468 162676 261480
rect 162728 261508 162734 261520
rect 176654 261508 176660 261520
rect 162728 261480 176660 261508
rect 162728 261468 162734 261480
rect 176654 261468 176660 261480
rect 176712 261468 176718 261520
rect 295334 261128 295340 261180
rect 295392 261168 295398 261180
rect 297450 261168 297456 261180
rect 295392 261140 297456 261168
rect 295392 261128 295398 261140
rect 297450 261128 297456 261140
rect 297508 261128 297514 261180
rect 66070 260924 66076 260976
rect 66128 260964 66134 260976
rect 68186 260964 68192 260976
rect 66128 260936 68192 260964
rect 66128 260924 66134 260936
rect 68186 260924 68192 260936
rect 68244 260924 68250 260976
rect 56318 260856 56324 260908
rect 56376 260896 56382 260908
rect 67726 260896 67732 260908
rect 56376 260868 67732 260896
rect 56376 260856 56382 260868
rect 67726 260856 67732 260868
rect 67784 260856 67790 260908
rect 121546 260856 121552 260908
rect 121604 260896 121610 260908
rect 155310 260896 155316 260908
rect 121604 260868 155316 260896
rect 121604 260856 121610 260868
rect 155310 260856 155316 260868
rect 155368 260856 155374 260908
rect 39942 260788 39948 260840
rect 40000 260828 40006 260840
rect 67634 260828 67640 260840
rect 40000 260800 67640 260828
rect 40000 260788 40006 260800
rect 67634 260788 67640 260800
rect 67692 260788 67698 260840
rect 360838 260788 360844 260840
rect 360896 260828 360902 260840
rect 386874 260828 386880 260840
rect 360896 260800 386880 260828
rect 360896 260788 360902 260800
rect 386874 260788 386880 260800
rect 386932 260788 386938 260840
rect 572622 260788 572628 260840
rect 572680 260828 572686 260840
rect 581178 260828 581184 260840
rect 572680 260800 581184 260828
rect 572680 260788 572686 260800
rect 581178 260788 581184 260800
rect 581236 260788 581242 260840
rect 575566 260720 575572 260772
rect 575624 260760 575630 260772
rect 576302 260760 576308 260772
rect 575624 260732 576308 260760
rect 575624 260720 575630 260732
rect 576302 260720 576308 260732
rect 576360 260720 576366 260772
rect 122374 260108 122380 260160
rect 122432 260148 122438 260160
rect 165154 260148 165160 260160
rect 122432 260120 165160 260148
rect 122432 260108 122438 260120
rect 165154 260108 165160 260120
rect 165212 260108 165218 260160
rect 121454 259496 121460 259548
rect 121512 259536 121518 259548
rect 146938 259536 146944 259548
rect 121512 259508 146944 259536
rect 121512 259496 121518 259508
rect 146938 259496 146944 259508
rect 146996 259496 147002 259548
rect 63218 259428 63224 259480
rect 63276 259468 63282 259480
rect 67634 259468 67640 259480
rect 63276 259440 67640 259468
rect 63276 259428 63282 259440
rect 67634 259428 67640 259440
rect 67692 259428 67698 259480
rect 121546 259428 121552 259480
rect 121604 259468 121610 259480
rect 153930 259468 153936 259480
rect 121604 259440 153936 259468
rect 121604 259428 121610 259440
rect 153930 259428 153936 259440
rect 153988 259428 153994 259480
rect 166902 259428 166908 259480
rect 166960 259468 166966 259480
rect 176654 259468 176660 259480
rect 166960 259440 176660 259468
rect 166960 259428 166966 259440
rect 176654 259428 176660 259440
rect 176712 259428 176718 259480
rect 576302 258680 576308 258732
rect 576360 258720 576366 258732
rect 580166 258720 580172 258732
rect 576360 258692 580172 258720
rect 576360 258680 576366 258692
rect 580166 258680 580172 258692
rect 580224 258680 580230 258732
rect 60458 258136 60464 258188
rect 60516 258176 60522 258188
rect 67634 258176 67640 258188
rect 60516 258148 67640 258176
rect 60516 258136 60522 258148
rect 67634 258136 67640 258148
rect 67692 258136 67698 258188
rect 121454 258136 121460 258188
rect 121512 258176 121518 258188
rect 148502 258176 148508 258188
rect 121512 258148 148508 258176
rect 121512 258136 121518 258148
rect 148502 258136 148508 258148
rect 148560 258136 148566 258188
rect 54846 258068 54852 258120
rect 54904 258108 54910 258120
rect 67726 258108 67732 258120
rect 54904 258080 67732 258108
rect 54904 258068 54910 258080
rect 67726 258068 67732 258080
rect 67784 258068 67790 258120
rect 121546 258068 121552 258120
rect 121604 258108 121610 258120
rect 167638 258108 167644 258120
rect 121604 258080 167644 258108
rect 121604 258068 121610 258080
rect 167638 258068 167644 258080
rect 167696 258068 167702 258120
rect 60642 258000 60648 258052
rect 60700 258040 60706 258052
rect 67634 258040 67640 258052
rect 60700 258012 67640 258040
rect 60700 258000 60706 258012
rect 67634 258000 67640 258012
rect 67692 258000 67698 258052
rect 17218 257320 17224 257372
rect 17276 257360 17282 257372
rect 60642 257360 60648 257372
rect 17276 257332 60648 257360
rect 17276 257320 17282 257332
rect 60642 257320 60648 257332
rect 60700 257320 60706 257372
rect 156506 257320 156512 257372
rect 156564 257360 156570 257372
rect 179046 257360 179052 257372
rect 156564 257332 179052 257360
rect 156564 257320 156570 257332
rect 179046 257320 179052 257332
rect 179104 257320 179110 257372
rect 121546 256776 121552 256828
rect 121604 256816 121610 256828
rect 144270 256816 144276 256828
rect 121604 256788 144276 256816
rect 121604 256776 121610 256788
rect 144270 256776 144276 256788
rect 144328 256776 144334 256828
rect 55122 256708 55128 256760
rect 55180 256748 55186 256760
rect 67634 256748 67640 256760
rect 55180 256720 67640 256748
rect 55180 256708 55186 256720
rect 67634 256708 67640 256720
rect 67692 256708 67698 256760
rect 121454 256708 121460 256760
rect 121512 256748 121518 256760
rect 175918 256748 175924 256760
rect 121512 256720 175924 256748
rect 121512 256708 121518 256720
rect 175918 256708 175924 256720
rect 175976 256708 175982 256760
rect 360838 256708 360844 256760
rect 360896 256748 360902 256760
rect 363782 256748 363788 256760
rect 360896 256720 363788 256748
rect 360896 256708 360902 256720
rect 363782 256708 363788 256720
rect 363840 256708 363846 256760
rect 121546 255348 121552 255400
rect 121604 255388 121610 255400
rect 149882 255388 149888 255400
rect 121604 255360 149888 255388
rect 121604 255348 121610 255360
rect 149882 255348 149888 255360
rect 149940 255348 149946 255400
rect 60550 255280 60556 255332
rect 60608 255320 60614 255332
rect 67634 255320 67640 255332
rect 60608 255292 67640 255320
rect 60608 255280 60614 255292
rect 67634 255280 67640 255292
rect 67692 255280 67698 255332
rect 121454 255280 121460 255332
rect 121512 255320 121518 255332
rect 159450 255320 159456 255332
rect 121512 255292 159456 255320
rect 121512 255280 121518 255292
rect 159450 255280 159456 255292
rect 159508 255280 159514 255332
rect 355410 255280 355416 255332
rect 355468 255320 355474 255332
rect 386874 255320 386880 255332
rect 355468 255292 386880 255320
rect 355468 255280 355474 255292
rect 386874 255280 386880 255292
rect 386932 255280 386938 255332
rect 2774 254056 2780 254108
rect 2832 254096 2838 254108
rect 4798 254096 4804 254108
rect 2832 254068 4804 254096
rect 2832 254056 2838 254068
rect 4798 254056 4804 254068
rect 4856 254056 4862 254108
rect 157334 253988 157340 254040
rect 157392 254028 157398 254040
rect 158438 254028 158444 254040
rect 157392 254000 158444 254028
rect 157392 253988 157398 254000
rect 158438 253988 158444 254000
rect 158496 254028 158502 254040
rect 176654 254028 176660 254040
rect 158496 254000 176660 254028
rect 158496 253988 158502 254000
rect 176654 253988 176660 254000
rect 176712 253988 176718 254040
rect 63126 253920 63132 253972
rect 63184 253960 63190 253972
rect 67726 253960 67732 253972
rect 63184 253932 67732 253960
rect 63184 253920 63190 253932
rect 67726 253920 67732 253932
rect 67784 253920 67790 253972
rect 121454 253920 121460 253972
rect 121512 253960 121518 253972
rect 171870 253960 171876 253972
rect 121512 253932 171876 253960
rect 121512 253920 121518 253932
rect 171870 253920 171876 253932
rect 171928 253920 171934 253972
rect 295610 253920 295616 253972
rect 295668 253960 295674 253972
rect 298922 253960 298928 253972
rect 295668 253932 298928 253960
rect 295668 253920 295674 253932
rect 298922 253920 298928 253932
rect 298980 253920 298986 253972
rect 60734 253852 60740 253904
rect 60792 253892 60798 253904
rect 62022 253892 62028 253904
rect 60792 253864 62028 253892
rect 60792 253852 60798 253864
rect 62022 253852 62028 253864
rect 62080 253892 62086 253904
rect 67634 253892 67640 253904
rect 62080 253864 67640 253892
rect 62080 253852 62086 253864
rect 67634 253852 67640 253864
rect 67692 253852 67698 253904
rect 302142 253852 302148 253904
rect 302200 253892 302206 253904
rect 306374 253892 306380 253904
rect 302200 253864 306380 253892
rect 302200 253852 302206 253864
rect 306374 253852 306380 253864
rect 306432 253852 306438 253904
rect 26878 253172 26884 253224
rect 26936 253212 26942 253224
rect 60734 253212 60740 253224
rect 26936 253184 60740 253212
rect 26936 253172 26942 253184
rect 60734 253172 60740 253184
rect 60792 253172 60798 253224
rect 64506 253172 64512 253224
rect 64564 253212 64570 253224
rect 68278 253212 68284 253224
rect 64564 253184 68284 253212
rect 64564 253172 64570 253184
rect 68278 253172 68284 253184
rect 68336 253172 68342 253224
rect 298830 253172 298836 253224
rect 298888 253212 298894 253224
rect 299566 253212 299572 253224
rect 298888 253184 299572 253212
rect 298888 253172 298894 253184
rect 299566 253172 299572 253184
rect 299624 253172 299630 253224
rect 121546 252628 121552 252680
rect 121604 252668 121610 252680
rect 152642 252668 152648 252680
rect 121604 252640 152648 252668
rect 121604 252628 121610 252640
rect 152642 252628 152648 252640
rect 152700 252628 152706 252680
rect 121454 252560 121460 252612
rect 121512 252600 121518 252612
rect 170398 252600 170404 252612
rect 121512 252572 170404 252600
rect 121512 252560 121518 252572
rect 170398 252560 170404 252572
rect 170456 252560 170462 252612
rect 327810 252560 327816 252612
rect 327868 252600 327874 252612
rect 386874 252600 386880 252612
rect 327868 252572 386880 252600
rect 327868 252560 327874 252572
rect 386874 252560 386880 252572
rect 386932 252560 386938 252612
rect 297174 252220 297180 252272
rect 297232 252260 297238 252272
rect 301498 252260 301504 252272
rect 297232 252232 301504 252260
rect 297232 252220 297238 252232
rect 301498 252220 301504 252232
rect 301556 252220 301562 252272
rect 60642 251812 60648 251864
rect 60700 251852 60706 251864
rect 68370 251852 68376 251864
rect 60700 251824 68376 251852
rect 60700 251812 60706 251824
rect 68370 251812 68376 251824
rect 68428 251812 68434 251864
rect 121454 251268 121460 251320
rect 121512 251308 121518 251320
rect 137462 251308 137468 251320
rect 121512 251280 137468 251308
rect 121512 251268 121518 251280
rect 137462 251268 137468 251280
rect 137520 251268 137526 251320
rect 121546 251200 121552 251252
rect 121604 251240 121610 251252
rect 174630 251240 174636 251252
rect 121604 251212 174636 251240
rect 121604 251200 121610 251212
rect 174630 251200 174636 251212
rect 174688 251200 174694 251252
rect 572622 251132 572628 251184
rect 572680 251172 572686 251184
rect 582466 251172 582472 251184
rect 572680 251144 582472 251172
rect 572680 251132 572686 251144
rect 582466 251132 582472 251144
rect 582524 251132 582530 251184
rect 120718 250996 120724 251048
rect 120776 251036 120782 251048
rect 124950 251036 124956 251048
rect 120776 251008 124956 251036
rect 120776 250996 120782 251008
rect 124950 250996 124956 251008
rect 125008 250996 125014 251048
rect 64598 249840 64604 249892
rect 64656 249880 64662 249892
rect 67634 249880 67640 249892
rect 64656 249852 67640 249880
rect 64656 249840 64662 249852
rect 67634 249840 67640 249852
rect 67692 249840 67698 249892
rect 59078 249772 59084 249824
rect 59136 249812 59142 249824
rect 67726 249812 67732 249824
rect 59136 249784 67732 249812
rect 59136 249772 59142 249784
rect 67726 249772 67732 249784
rect 67784 249772 67790 249824
rect 121454 249772 121460 249824
rect 121512 249812 121518 249824
rect 131942 249812 131948 249824
rect 121512 249784 131948 249812
rect 121512 249772 121518 249784
rect 131942 249772 131948 249784
rect 132000 249772 132006 249824
rect 55030 249704 55036 249756
rect 55088 249744 55094 249756
rect 67634 249744 67640 249756
rect 55088 249716 67640 249744
rect 55088 249704 55094 249716
rect 67634 249704 67640 249716
rect 67692 249704 67698 249756
rect 57790 248412 57796 248464
rect 57848 248452 57854 248464
rect 67634 248452 67640 248464
rect 57848 248424 67640 248452
rect 57848 248412 57854 248424
rect 67634 248412 67640 248424
rect 67692 248412 67698 248464
rect 121454 248412 121460 248464
rect 121512 248452 121518 248464
rect 174538 248452 174544 248464
rect 121512 248424 174544 248452
rect 121512 248412 121518 248424
rect 174538 248412 174544 248424
rect 174596 248412 174602 248464
rect 572622 248208 572628 248260
rect 572680 248248 572686 248260
rect 576946 248248 576952 248260
rect 572680 248220 576952 248248
rect 572680 248208 572686 248220
rect 576946 248208 576952 248220
rect 577004 248208 577010 248260
rect 122282 247664 122288 247716
rect 122340 247704 122346 247716
rect 166994 247704 167000 247716
rect 122340 247676 167000 247704
rect 122340 247664 122346 247676
rect 166994 247664 167000 247676
rect 167052 247664 167058 247716
rect 301314 247664 301320 247716
rect 301372 247704 301378 247716
rect 307662 247704 307668 247716
rect 301372 247676 307668 247704
rect 301372 247664 301378 247676
rect 307662 247664 307668 247676
rect 307720 247704 307726 247716
rect 378778 247704 378784 247716
rect 307720 247676 378784 247704
rect 307720 247664 307726 247676
rect 378778 247664 378784 247676
rect 378836 247664 378842 247716
rect 62022 247120 62028 247172
rect 62080 247160 62086 247172
rect 67634 247160 67640 247172
rect 62080 247132 67640 247160
rect 62080 247120 62086 247132
rect 67634 247120 67640 247132
rect 67692 247120 67698 247172
rect 59170 247052 59176 247104
rect 59228 247092 59234 247104
rect 67726 247092 67732 247104
rect 59228 247064 67732 247092
rect 59228 247052 59234 247064
rect 67726 247052 67732 247064
rect 67784 247052 67790 247104
rect 121454 247052 121460 247104
rect 121512 247092 121518 247104
rect 126422 247092 126428 247104
rect 121512 247064 126428 247092
rect 121512 247052 121518 247064
rect 126422 247052 126428 247064
rect 126480 247052 126486 247104
rect 295518 247052 295524 247104
rect 295576 247092 295582 247104
rect 301038 247092 301044 247104
rect 295576 247064 301044 247092
rect 295576 247052 295582 247064
rect 301038 247052 301044 247064
rect 301096 247092 301102 247104
rect 301314 247092 301320 247104
rect 301096 247064 301320 247092
rect 301096 247052 301102 247064
rect 301314 247052 301320 247064
rect 301372 247052 301378 247104
rect 379422 246984 379428 247036
rect 379480 247024 379486 247036
rect 386874 247024 386880 247036
rect 379480 246996 386880 247024
rect 379480 246984 379486 246996
rect 386874 246984 386880 246996
rect 386932 246984 386938 247036
rect 353294 246372 353300 246424
rect 353352 246412 353358 246424
rect 379422 246412 379428 246424
rect 353352 246384 379428 246412
rect 353352 246372 353358 246384
rect 379422 246372 379428 246384
rect 379480 246372 379486 246424
rect 295518 246304 295524 246356
rect 295576 246344 295582 246356
rect 298186 246344 298192 246356
rect 295576 246316 298192 246344
rect 295576 246304 295582 246316
rect 298186 246304 298192 246316
rect 298244 246344 298250 246356
rect 358078 246344 358084 246356
rect 298244 246316 358084 246344
rect 298244 246304 298250 246316
rect 358078 246304 358084 246316
rect 358136 246304 358142 246356
rect 121454 245760 121460 245812
rect 121512 245800 121518 245812
rect 140222 245800 140228 245812
rect 121512 245772 140228 245800
rect 121512 245760 121518 245772
rect 140222 245760 140228 245772
rect 140280 245760 140286 245812
rect 121546 245692 121552 245744
rect 121604 245732 121610 245744
rect 147122 245732 147128 245744
rect 121604 245704 147128 245732
rect 121604 245692 121610 245704
rect 147122 245692 147128 245704
rect 147180 245692 147186 245744
rect 124122 245624 124128 245676
rect 124180 245664 124186 245676
rect 176654 245664 176660 245676
rect 124180 245636 176660 245664
rect 124180 245624 124186 245636
rect 176654 245624 176660 245636
rect 176712 245624 176718 245676
rect 50338 245556 50344 245608
rect 50396 245596 50402 245608
rect 68094 245596 68100 245608
rect 50396 245568 68100 245596
rect 50396 245556 50402 245568
rect 68094 245556 68100 245568
rect 68152 245556 68158 245608
rect 582742 245556 582748 245608
rect 582800 245596 582806 245608
rect 583662 245596 583668 245608
rect 582800 245568 583668 245596
rect 582800 245556 582806 245568
rect 583662 245556 583668 245568
rect 583720 245556 583726 245608
rect 342990 244876 342996 244928
rect 343048 244916 343054 244928
rect 387518 244916 387524 244928
rect 343048 244888 387524 244916
rect 343048 244876 343054 244888
rect 387518 244876 387524 244888
rect 387576 244876 387582 244928
rect 121454 244332 121460 244384
rect 121512 244372 121518 244384
rect 160094 244372 160100 244384
rect 121512 244344 160100 244372
rect 121512 244332 121518 244344
rect 160094 244332 160100 244344
rect 160152 244332 160158 244384
rect 65886 244264 65892 244316
rect 65944 244304 65950 244316
rect 68002 244304 68008 244316
rect 65944 244276 68008 244304
rect 65944 244264 65950 244276
rect 68002 244264 68008 244276
rect 68060 244264 68066 244316
rect 121546 244264 121552 244316
rect 121604 244304 121610 244316
rect 173250 244304 173256 244316
rect 121604 244276 173256 244304
rect 121604 244264 121610 244276
rect 173250 244264 173256 244276
rect 173308 244264 173314 244316
rect 577498 244264 577504 244316
rect 577556 244304 577562 244316
rect 582742 244304 582748 244316
rect 577556 244276 582748 244304
rect 577556 244264 577562 244276
rect 582742 244264 582748 244276
rect 582800 244264 582806 244316
rect 121454 244196 121460 244248
rect 121512 244236 121518 244248
rect 140038 244236 140044 244248
rect 121512 244208 140044 244236
rect 121512 244196 121518 244208
rect 140038 244196 140044 244208
rect 140096 244196 140102 244248
rect 295794 244196 295800 244248
rect 295852 244236 295858 244248
rect 353294 244236 353300 244248
rect 295852 244208 353300 244236
rect 295852 244196 295858 244208
rect 353294 244196 353300 244208
rect 353352 244196 353358 244248
rect 363782 243516 363788 243568
rect 363840 243556 363846 243568
rect 364242 243556 364248 243568
rect 363840 243528 364248 243556
rect 363840 243516 363846 243528
rect 364242 243516 364248 243528
rect 364300 243556 364306 243568
rect 386598 243556 386604 243568
rect 364300 243528 386604 243556
rect 364300 243516 364306 243528
rect 386598 243516 386604 243528
rect 386656 243516 386662 243568
rect 121546 242904 121552 242956
rect 121604 242944 121610 242956
rect 166350 242944 166356 242956
rect 121604 242916 166356 242944
rect 121604 242904 121610 242916
rect 166350 242904 166356 242916
rect 166408 242904 166414 242956
rect 121638 242836 121644 242888
rect 121696 242876 121702 242888
rect 130470 242876 130476 242888
rect 121696 242848 130476 242876
rect 121696 242836 121702 242848
rect 130470 242836 130476 242848
rect 130528 242836 130534 242888
rect 120902 242224 120908 242276
rect 120960 242264 120966 242276
rect 149974 242264 149980 242276
rect 120960 242236 149980 242264
rect 120960 242224 120966 242236
rect 149974 242224 149980 242236
rect 150032 242224 150038 242276
rect 121454 242156 121460 242208
rect 121512 242196 121518 242208
rect 160738 242196 160744 242208
rect 121512 242168 160744 242196
rect 121512 242156 121518 242168
rect 160738 242156 160744 242168
rect 160796 242156 160802 242208
rect 296714 242156 296720 242208
rect 296772 242196 296778 242208
rect 333974 242196 333980 242208
rect 296772 242168 333980 242196
rect 296772 242156 296778 242168
rect 333974 242156 333980 242168
rect 334032 242156 334038 242208
rect 337470 242156 337476 242208
rect 337528 242196 337534 242208
rect 387150 242196 387156 242208
rect 337528 242168 387156 242196
rect 337528 242156 337534 242168
rect 387150 242156 387156 242168
rect 387208 242156 387214 242208
rect 61746 241612 61752 241664
rect 61804 241652 61810 241664
rect 67634 241652 67640 241664
rect 61804 241624 67640 241652
rect 61804 241612 61810 241624
rect 67634 241612 67640 241624
rect 67692 241612 67698 241664
rect 168374 241476 168380 241528
rect 168432 241516 168438 241528
rect 169662 241516 169668 241528
rect 168432 241488 169668 241516
rect 168432 241476 168438 241488
rect 169662 241476 169668 241488
rect 169720 241516 169726 241528
rect 177574 241516 177580 241528
rect 169720 241488 177580 241516
rect 169720 241476 169726 241488
rect 177574 241476 177580 241488
rect 177632 241476 177638 241528
rect 161198 241408 161204 241460
rect 161256 241448 161262 241460
rect 377674 241448 377680 241460
rect 161256 241420 377680 241448
rect 161256 241408 161262 241420
rect 377674 241408 377680 241420
rect 377732 241408 377738 241460
rect 572622 241408 572628 241460
rect 572680 241448 572686 241460
rect 582558 241448 582564 241460
rect 572680 241420 582564 241448
rect 572680 241408 572686 241420
rect 582558 241408 582564 241420
rect 582616 241408 582622 241460
rect 141510 240728 141516 240780
rect 141568 240768 141574 240780
rect 141568 240740 184060 240768
rect 141568 240728 141574 240740
rect 184032 240644 184060 240740
rect 298922 240728 298928 240780
rect 298980 240768 298986 240780
rect 335354 240768 335360 240780
rect 298980 240740 335360 240768
rect 298980 240728 298986 240740
rect 335354 240728 335360 240740
rect 335412 240728 335418 240780
rect 173802 240592 173808 240644
rect 173860 240632 173866 240644
rect 180426 240632 180432 240644
rect 173860 240604 180432 240632
rect 173860 240592 173866 240604
rect 180426 240592 180432 240604
rect 180484 240592 180490 240644
rect 184014 240592 184020 240644
rect 184072 240592 184078 240644
rect 291930 240592 291936 240644
rect 291988 240632 291994 240644
rect 293310 240632 293316 240644
rect 291988 240604 293316 240632
rect 291988 240592 291994 240604
rect 293310 240592 293316 240604
rect 293368 240592 293374 240644
rect 3418 240116 3424 240168
rect 3476 240156 3482 240168
rect 14458 240156 14464 240168
rect 3476 240128 14464 240156
rect 3476 240116 3482 240128
rect 14458 240116 14464 240128
rect 14516 240116 14522 240168
rect 121454 240116 121460 240168
rect 121512 240156 121518 240168
rect 148594 240156 148600 240168
rect 121512 240128 148600 240156
rect 121512 240116 121518 240128
rect 148594 240116 148600 240128
rect 148652 240116 148658 240168
rect 363598 240116 363604 240168
rect 363656 240156 363662 240168
rect 386874 240156 386880 240168
rect 363656 240128 386880 240156
rect 363656 240116 363662 240128
rect 386874 240116 386880 240128
rect 386932 240116 386938 240168
rect 159910 240048 159916 240100
rect 159968 240088 159974 240100
rect 362310 240088 362316 240100
rect 159968 240060 362316 240088
rect 159968 240048 159974 240060
rect 362310 240048 362316 240060
rect 362368 240048 362374 240100
rect 180426 239980 180432 240032
rect 180484 240020 180490 240032
rect 359642 240020 359648 240032
rect 180484 239992 359648 240020
rect 180484 239980 180490 239992
rect 359642 239980 359648 239992
rect 359700 239980 359706 240032
rect 166994 239912 167000 239964
rect 167052 239952 167058 239964
rect 298738 239952 298744 239964
rect 167052 239924 298744 239952
rect 167052 239912 167058 239924
rect 298738 239912 298744 239924
rect 298796 239912 298802 239964
rect 179506 239844 179512 239896
rect 179564 239884 179570 239896
rect 180012 239884 180018 239896
rect 179564 239856 180018 239884
rect 179564 239844 179570 239856
rect 180012 239844 180018 239856
rect 180070 239844 180076 239896
rect 289814 239844 289820 239896
rect 289872 239884 289878 239896
rect 294230 239884 294236 239896
rect 289872 239856 294236 239884
rect 289872 239844 289878 239856
rect 294230 239844 294236 239856
rect 294288 239844 294294 239896
rect 63218 239368 63224 239420
rect 63276 239408 63282 239420
rect 76558 239408 76564 239420
rect 63276 239380 76564 239408
rect 63276 239368 63282 239380
rect 76558 239368 76564 239380
rect 76616 239368 76622 239420
rect 111058 239368 111064 239420
rect 111116 239408 111122 239420
rect 295610 239408 295616 239420
rect 111116 239380 295616 239408
rect 111116 239368 111122 239380
rect 295610 239368 295616 239380
rect 295668 239368 295674 239420
rect 121546 238892 121552 238944
rect 121604 238932 121610 238944
rect 148962 238932 148968 238944
rect 121604 238904 148968 238932
rect 121604 238892 121610 238904
rect 148962 238892 148968 238904
rect 149020 238892 149026 238944
rect 110414 238824 110420 238876
rect 110472 238864 110478 238876
rect 110598 238864 110604 238876
rect 110472 238836 110604 238864
rect 110472 238824 110478 238836
rect 110598 238824 110604 238836
rect 110656 238864 110662 238876
rect 142798 238864 142804 238876
rect 110656 238836 142804 238864
rect 110656 238824 110662 238836
rect 142798 238824 142804 238836
rect 142856 238824 142862 238876
rect 148410 238824 148416 238876
rect 148468 238864 148474 238876
rect 195974 238864 195980 238876
rect 148468 238836 195980 238864
rect 148468 238824 148474 238836
rect 195974 238824 195980 238836
rect 196032 238824 196038 238876
rect 61838 238756 61844 238808
rect 61896 238796 61902 238808
rect 180886 238796 180892 238808
rect 61896 238768 180892 238796
rect 61896 238756 61902 238768
rect 180886 238756 180892 238768
rect 180944 238756 180950 238808
rect 255222 238756 255228 238808
rect 255280 238796 255286 238808
rect 387058 238796 387064 238808
rect 255280 238768 387064 238796
rect 255280 238756 255286 238768
rect 387058 238756 387064 238768
rect 387116 238756 387122 238808
rect 25498 238688 25504 238740
rect 25556 238728 25562 238740
rect 86770 238728 86776 238740
rect 25556 238700 86776 238728
rect 25556 238688 25562 238700
rect 86770 238688 86776 238700
rect 86828 238688 86834 238740
rect 114462 238688 114468 238740
rect 114520 238728 114526 238740
rect 125594 238728 125600 238740
rect 114520 238700 125600 238728
rect 114520 238688 114526 238700
rect 125594 238688 125600 238700
rect 125652 238688 125658 238740
rect 172330 238688 172336 238740
rect 172388 238728 172394 238740
rect 374822 238728 374828 238740
rect 172388 238700 374828 238728
rect 172388 238688 172394 238700
rect 374822 238688 374828 238700
rect 374880 238688 374886 238740
rect 81618 238620 81624 238672
rect 81676 238660 81682 238672
rect 279510 238660 279516 238672
rect 81676 238632 279516 238660
rect 81676 238620 81682 238632
rect 279510 238620 279516 238632
rect 279568 238620 279574 238672
rect 287882 238620 287888 238672
rect 287940 238660 287946 238672
rect 377582 238660 377588 238672
rect 287940 238632 377588 238660
rect 287940 238620 287946 238632
rect 377582 238620 377588 238632
rect 377640 238620 377646 238672
rect 58618 238552 58624 238604
rect 58676 238592 58682 238604
rect 82262 238592 82268 238604
rect 58676 238564 82268 238592
rect 58676 238552 58682 238564
rect 82262 238552 82268 238564
rect 82320 238552 82326 238604
rect 82906 238552 82912 238604
rect 82964 238592 82970 238604
rect 111058 238592 111064 238604
rect 82964 238564 111064 238592
rect 82964 238552 82970 238564
rect 111058 238552 111064 238564
rect 111116 238552 111122 238604
rect 117682 238552 117688 238604
rect 117740 238592 117746 238604
rect 250806 238592 250812 238604
rect 117740 238564 250812 238592
rect 117740 238552 117746 238564
rect 250806 238552 250812 238564
rect 250864 238552 250870 238604
rect 273990 238552 273996 238604
rect 274048 238592 274054 238604
rect 377490 238592 377496 238604
rect 274048 238564 377496 238592
rect 274048 238552 274054 238564
rect 377490 238552 377496 238564
rect 377548 238552 377554 238604
rect 86770 238484 86776 238536
rect 86828 238524 86834 238536
rect 210418 238524 210424 238536
rect 86828 238496 210424 238524
rect 86828 238484 86834 238496
rect 210418 238484 210424 238496
rect 210476 238484 210482 238536
rect 278038 238484 278044 238536
rect 278096 238524 278102 238536
rect 365070 238524 365076 238536
rect 278096 238496 365076 238524
rect 278096 238484 278102 238496
rect 365070 238484 365076 238496
rect 365128 238484 365134 238536
rect 118326 238416 118332 238468
rect 118384 238456 118390 238468
rect 240502 238456 240508 238468
rect 118384 238428 240508 238456
rect 118384 238416 118390 238428
rect 240502 238416 240508 238428
rect 240560 238416 240566 238468
rect 250806 238416 250812 238468
rect 250864 238456 250870 238468
rect 300210 238456 300216 238468
rect 250864 238428 300216 238456
rect 250864 238416 250870 238428
rect 300210 238416 300216 238428
rect 300268 238416 300274 238468
rect 89346 238348 89352 238400
rect 89404 238388 89410 238400
rect 138658 238388 138664 238400
rect 89404 238360 138664 238388
rect 89404 238348 89410 238360
rect 138658 238348 138664 238360
rect 138716 238348 138722 238400
rect 204806 238348 204812 238400
rect 204864 238388 204870 238400
rect 255222 238388 255228 238400
rect 204864 238360 255228 238388
rect 204864 238348 204870 238360
rect 255222 238348 255228 238360
rect 255280 238348 255286 238400
rect 263042 238348 263048 238400
rect 263100 238388 263106 238400
rect 297542 238388 297548 238400
rect 263100 238360 297548 238388
rect 263100 238348 263106 238360
rect 297542 238348 297548 238360
rect 297600 238348 297606 238400
rect 77110 238076 77116 238128
rect 77168 238116 77174 238128
rect 106918 238116 106924 238128
rect 77168 238088 106924 238116
rect 77168 238076 77174 238088
rect 106918 238076 106924 238088
rect 106976 238076 106982 238128
rect 253106 238076 253112 238128
rect 253164 238116 253170 238128
rect 263594 238116 263600 238128
rect 253164 238088 263600 238116
rect 253164 238076 253170 238088
rect 263594 238076 263600 238088
rect 263652 238076 263658 238128
rect 63310 238008 63316 238060
rect 63368 238048 63374 238060
rect 117222 238048 117228 238060
rect 63368 238020 117228 238048
rect 63368 238008 63374 238020
rect 117222 238008 117228 238020
rect 117280 238008 117286 238060
rect 236270 238008 236276 238060
rect 236328 238048 236334 238060
rect 273898 238048 273904 238060
rect 236328 238020 273904 238048
rect 236328 238008 236334 238020
rect 273898 238008 273904 238020
rect 273956 238008 273962 238060
rect 79042 237396 79048 237448
rect 79100 237436 79106 237448
rect 86218 237436 86224 237448
rect 79100 237408 86224 237436
rect 79100 237396 79106 237408
rect 86218 237396 86224 237408
rect 86276 237396 86282 237448
rect 14458 237328 14464 237380
rect 14516 237368 14522 237380
rect 103514 237368 103520 237380
rect 14516 237340 103520 237368
rect 14516 237328 14522 237340
rect 103514 237328 103520 237340
rect 103572 237368 103578 237380
rect 104710 237368 104716 237380
rect 103572 237340 104716 237368
rect 103572 237328 103578 237340
rect 104710 237328 104716 237340
rect 104768 237328 104774 237380
rect 113174 237328 113180 237380
rect 113232 237368 113238 237380
rect 354674 237368 354680 237380
rect 113232 237340 354680 237368
rect 113232 237328 113238 237340
rect 354674 237328 354680 237340
rect 354732 237368 354738 237380
rect 355410 237368 355416 237380
rect 354732 237340 355416 237368
rect 354732 237328 354738 237340
rect 355410 237328 355416 237340
rect 355468 237328 355474 237380
rect 109678 237260 109684 237312
rect 109736 237300 109742 237312
rect 140682 237300 140688 237312
rect 109736 237272 140688 237300
rect 109736 237260 109742 237272
rect 140682 237260 140688 237272
rect 140740 237300 140746 237312
rect 365162 237300 365168 237312
rect 140740 237272 365168 237300
rect 140740 237260 140746 237272
rect 365162 237260 365168 237272
rect 365220 237260 365226 237312
rect 99006 237192 99012 237244
rect 99064 237232 99070 237244
rect 120994 237232 121000 237244
rect 99064 237204 121000 237232
rect 99064 237192 99070 237204
rect 120994 237192 121000 237204
rect 121052 237192 121058 237244
rect 157150 237192 157156 237244
rect 157208 237232 157214 237244
rect 345658 237232 345664 237244
rect 157208 237204 345664 237232
rect 157208 237192 157214 237204
rect 345658 237192 345664 237204
rect 345716 237192 345722 237244
rect 175918 237124 175924 237176
rect 175976 237164 175982 237176
rect 295426 237164 295432 237176
rect 175976 237136 295432 237164
rect 175976 237124 175982 237136
rect 295426 237124 295432 237136
rect 295484 237124 295490 237176
rect 269850 237056 269856 237108
rect 269908 237096 269914 237108
rect 319530 237096 319536 237108
rect 269908 237068 319536 237096
rect 269908 237056 269914 237068
rect 319530 237056 319536 237068
rect 319588 237056 319594 237108
rect 169110 236716 169116 236768
rect 169168 236756 169174 236768
rect 192478 236756 192484 236768
rect 169168 236728 192484 236756
rect 169168 236716 169174 236728
rect 192478 236716 192484 236728
rect 192536 236716 192542 236768
rect 64506 236648 64512 236700
rect 64564 236688 64570 236700
rect 98638 236688 98644 236700
rect 64564 236660 98644 236688
rect 64564 236648 64570 236660
rect 98638 236648 98644 236660
rect 98696 236648 98702 236700
rect 167822 236648 167828 236700
rect 167880 236688 167886 236700
rect 273254 236688 273260 236700
rect 167880 236660 273260 236688
rect 167880 236648 167886 236660
rect 273254 236648 273260 236660
rect 273312 236648 273318 236700
rect 67542 235900 67548 235952
rect 67600 235940 67606 235952
rect 381630 235940 381636 235952
rect 67600 235912 381636 235940
rect 67600 235900 67606 235912
rect 381630 235900 381636 235912
rect 381688 235900 381694 235952
rect 4798 235832 4804 235884
rect 4856 235872 4862 235884
rect 112530 235872 112536 235884
rect 4856 235844 112536 235872
rect 4856 235832 4862 235844
rect 112530 235832 112536 235844
rect 112588 235872 112594 235884
rect 128998 235872 129004 235884
rect 112588 235844 129004 235872
rect 112588 235832 112594 235844
rect 128998 235832 129004 235844
rect 129056 235832 129062 235884
rect 154390 235832 154396 235884
rect 154448 235872 154454 235884
rect 373350 235872 373356 235884
rect 154448 235844 373356 235872
rect 154448 235832 154454 235844
rect 373350 235832 373356 235844
rect 373408 235832 373414 235884
rect 119706 235764 119712 235816
rect 119764 235804 119770 235816
rect 323670 235804 323676 235816
rect 119764 235776 323676 235804
rect 119764 235764 119770 235776
rect 323670 235764 323676 235776
rect 323728 235764 323734 235816
rect 72602 235696 72608 235748
rect 72660 235736 72666 235748
rect 123662 235736 123668 235748
rect 72660 235708 123668 235736
rect 72660 235696 72666 235708
rect 123662 235696 123668 235708
rect 123720 235696 123726 235748
rect 162762 235696 162768 235748
rect 162820 235736 162826 235748
rect 366450 235736 366456 235748
rect 162820 235708 366456 235736
rect 162820 235696 162826 235708
rect 366450 235696 366456 235708
rect 366508 235696 366514 235748
rect 91278 235628 91284 235680
rect 91336 235668 91342 235680
rect 129274 235668 129280 235680
rect 91336 235640 129280 235668
rect 91336 235628 91342 235640
rect 129274 235628 129280 235640
rect 129332 235628 129338 235680
rect 174630 235628 174636 235680
rect 174688 235668 174694 235680
rect 273990 235668 273996 235680
rect 174688 235640 273996 235668
rect 174688 235628 174694 235640
rect 273990 235628 273996 235640
rect 274048 235628 274054 235680
rect 113818 235560 113824 235612
rect 113876 235600 113882 235612
rect 152458 235600 152464 235612
rect 113876 235572 152464 235600
rect 113876 235560 113882 235572
rect 152458 235560 152464 235572
rect 152516 235560 152522 235612
rect 265618 235560 265624 235612
rect 265676 235600 265682 235612
rect 310514 235600 310520 235612
rect 265676 235572 310520 235600
rect 265676 235560 265682 235572
rect 310514 235560 310520 235572
rect 310572 235560 310578 235612
rect 56318 235220 56324 235272
rect 56376 235260 56382 235272
rect 116578 235260 116584 235272
rect 56376 235232 116584 235260
rect 56376 235220 56382 235232
rect 116578 235220 116584 235232
rect 116636 235220 116642 235272
rect 380894 234812 380900 234864
rect 380952 234852 380958 234864
rect 381630 234852 381636 234864
rect 380952 234824 381636 234852
rect 380952 234812 380958 234824
rect 381630 234812 381636 234824
rect 381688 234812 381694 234864
rect 63126 234540 63132 234592
rect 63184 234580 63190 234592
rect 263042 234580 263048 234592
rect 63184 234552 263048 234580
rect 63184 234540 63190 234552
rect 263042 234540 263048 234552
rect 263100 234540 263106 234592
rect 572622 234540 572628 234592
rect 572680 234580 572686 234592
rect 581086 234580 581092 234592
rect 572680 234552 581092 234580
rect 572680 234540 572686 234552
rect 581086 234540 581092 234552
rect 581144 234540 581150 234592
rect 69290 234472 69296 234524
rect 69348 234512 69354 234524
rect 219250 234512 219256 234524
rect 69348 234484 219256 234512
rect 69348 234472 69354 234484
rect 219250 234472 219256 234484
rect 219308 234512 219314 234524
rect 369210 234512 369216 234524
rect 219308 234484 369216 234512
rect 219308 234472 219314 234484
rect 369210 234472 369216 234484
rect 369268 234472 369274 234524
rect 95786 234404 95792 234456
rect 95844 234444 95850 234456
rect 126974 234444 126980 234456
rect 95844 234416 126980 234444
rect 95844 234404 95850 234416
rect 126974 234404 126980 234416
rect 127032 234404 127038 234456
rect 140130 233996 140136 234048
rect 140188 234036 140194 234048
rect 273990 234036 273996 234048
rect 140188 234008 273996 234036
rect 140188 233996 140194 234008
rect 273990 233996 273996 234008
rect 274048 233996 274054 234048
rect 69106 233928 69112 233980
rect 69164 233968 69170 233980
rect 69750 233968 69756 233980
rect 69164 233940 69756 233968
rect 69164 233928 69170 233940
rect 69750 233928 69756 233940
rect 69808 233928 69814 233980
rect 74534 233928 74540 233980
rect 74592 233968 74598 233980
rect 75178 233968 75184 233980
rect 74592 233940 75184 233968
rect 74592 233928 74598 233940
rect 75178 233928 75184 233940
rect 75236 233928 75242 233980
rect 80054 233928 80060 233980
rect 80112 233968 80118 233980
rect 80974 233968 80980 233980
rect 80112 233940 80980 233968
rect 80112 233928 80118 233940
rect 80974 233928 80980 233940
rect 81032 233928 81038 233980
rect 84194 233928 84200 233980
rect 84252 233968 84258 233980
rect 84838 233968 84844 233980
rect 84252 233940 84844 233968
rect 84252 233928 84258 233940
rect 84838 233928 84844 233940
rect 84896 233928 84902 233980
rect 95142 233928 95148 233980
rect 95200 233968 95206 233980
rect 120718 233968 120724 233980
rect 95200 233940 120724 233968
rect 95200 233928 95206 233940
rect 120718 233928 120724 233940
rect 120776 233928 120782 233980
rect 242250 233928 242256 233980
rect 242308 233968 242314 233980
rect 386506 233968 386512 233980
rect 242308 233940 386512 233968
rect 242308 233928 242314 233940
rect 386506 233928 386512 233940
rect 386564 233928 386570 233980
rect 64598 233860 64604 233912
rect 64656 233900 64662 233912
rect 64656 233872 84194 233900
rect 64656 233860 64662 233872
rect 84166 233832 84194 233872
rect 86954 233860 86960 233912
rect 87012 233900 87018 233912
rect 88058 233900 88064 233912
rect 87012 233872 88064 233900
rect 87012 233860 87018 233872
rect 88058 233860 88064 233872
rect 88116 233860 88122 233912
rect 95234 233860 95240 233912
rect 95292 233900 95298 233912
rect 96430 233900 96436 233912
rect 95292 233872 96436 233900
rect 95292 233860 95298 233872
rect 96430 233860 96436 233872
rect 96488 233860 96494 233912
rect 100754 233860 100760 233912
rect 100812 233900 100818 233912
rect 101582 233900 101588 233912
rect 100812 233872 101588 233900
rect 100812 233860 100818 233872
rect 101582 233860 101588 233872
rect 101640 233860 101646 233912
rect 107654 233860 107660 233912
rect 107712 233900 107718 233912
rect 108666 233900 108672 233912
rect 107712 233872 108672 233900
rect 107712 233860 107718 233872
rect 108666 233860 108672 233872
rect 108724 233860 108730 233912
rect 114554 233860 114560 233912
rect 114612 233900 114618 233912
rect 115750 233900 115756 233912
rect 114612 233872 115756 233900
rect 114612 233860 114618 233872
rect 115750 233860 115756 233872
rect 115808 233860 115814 233912
rect 148962 233860 148968 233912
rect 149020 233900 149026 233912
rect 311158 233900 311164 233912
rect 149020 233872 311164 233900
rect 149020 233860 149026 233872
rect 311158 233860 311164 233872
rect 311216 233860 311222 233912
rect 361022 233860 361028 233912
rect 361080 233900 361086 233912
rect 386782 233900 386788 233912
rect 361080 233872 386788 233900
rect 361080 233860 361086 233872
rect 386782 233860 386788 233872
rect 386840 233860 386846 233912
rect 95878 233832 95884 233844
rect 84166 233804 95884 233832
rect 95878 233792 95884 233804
rect 95936 233792 95942 233844
rect 61654 233180 61660 233232
rect 61712 233220 61718 233232
rect 341518 233220 341524 233232
rect 61712 233192 341524 233220
rect 61712 233180 61718 233192
rect 341518 233180 341524 233192
rect 341576 233180 341582 233232
rect 86126 233112 86132 233164
rect 86184 233152 86190 233164
rect 157242 233152 157248 233164
rect 86184 233124 157248 233152
rect 86184 233112 86190 233124
rect 157242 233112 157248 233124
rect 157300 233112 157306 233164
rect 184014 233112 184020 233164
rect 184072 233152 184078 233164
rect 295610 233152 295616 233164
rect 184072 233124 295616 233152
rect 184072 233112 184078 233124
rect 295610 233112 295616 233124
rect 295668 233112 295674 233164
rect 325694 233152 325700 233164
rect 316006 233124 325700 233152
rect 76466 233044 76472 233096
rect 76524 233084 76530 233096
rect 134518 233084 134524 233096
rect 76524 233056 134524 233084
rect 76524 233044 76530 233056
rect 134518 233044 134524 233056
rect 134576 233044 134582 233096
rect 144362 233044 144368 233096
rect 144420 233084 144426 233096
rect 254670 233084 254676 233096
rect 144420 233056 254676 233084
rect 144420 233044 144426 233056
rect 254670 233044 254676 233056
rect 254728 233044 254734 233096
rect 273254 233044 273260 233096
rect 273312 233084 273318 233096
rect 316006 233084 316034 233124
rect 325694 233112 325700 233124
rect 325752 233152 325758 233164
rect 326338 233152 326344 233164
rect 325752 233124 326344 233152
rect 325752 233112 325758 233124
rect 326338 233112 326344 233124
rect 326396 233112 326402 233164
rect 273312 233056 316034 233084
rect 273312 233044 273318 233056
rect 70670 232568 70676 232620
rect 70728 232608 70734 232620
rect 88978 232608 88984 232620
rect 70728 232580 88984 232608
rect 70728 232568 70734 232580
rect 88978 232568 88984 232580
rect 89036 232568 89042 232620
rect 170490 232568 170496 232620
rect 170548 232608 170554 232620
rect 186958 232608 186964 232620
rect 170548 232580 186964 232608
rect 170548 232568 170554 232580
rect 186958 232568 186964 232580
rect 187016 232568 187022 232620
rect 1302 232500 1308 232552
rect 1360 232540 1366 232552
rect 120074 232540 120080 232552
rect 1360 232512 120080 232540
rect 1360 232500 1366 232512
rect 120074 232500 120080 232512
rect 120132 232500 120138 232552
rect 155310 232500 155316 232552
rect 155368 232540 155374 232552
rect 275278 232540 275284 232552
rect 155368 232512 275284 232540
rect 155368 232500 155374 232512
rect 275278 232500 275284 232512
rect 275336 232500 275342 232552
rect 129274 231752 129280 231804
rect 129332 231792 129338 231804
rect 367922 231792 367928 231804
rect 129332 231764 367928 231792
rect 129332 231752 129338 231764
rect 367922 231752 367928 231764
rect 367980 231752 367986 231804
rect 82262 231684 82268 231736
rect 82320 231724 82326 231736
rect 278038 231724 278044 231736
rect 82320 231696 278044 231724
rect 82320 231684 82326 231696
rect 278038 231684 278044 231696
rect 278096 231684 278102 231736
rect 279510 231684 279516 231736
rect 279568 231724 279574 231736
rect 280062 231724 280068 231736
rect 279568 231696 280068 231724
rect 279568 231684 279574 231696
rect 280062 231684 280068 231696
rect 280120 231724 280126 231736
rect 309134 231724 309140 231736
rect 280120 231696 309140 231724
rect 280120 231684 280126 231696
rect 309134 231684 309140 231696
rect 309192 231684 309198 231736
rect 104710 231616 104716 231668
rect 104768 231656 104774 231668
rect 293218 231656 293224 231668
rect 104768 231628 293224 231656
rect 104768 231616 104774 231628
rect 293218 231616 293224 231628
rect 293276 231616 293282 231668
rect 91922 231548 91928 231600
rect 91980 231588 91986 231600
rect 135898 231588 135904 231600
rect 91980 231560 135904 231588
rect 91980 231548 91986 231560
rect 135898 231548 135904 231560
rect 135956 231548 135962 231600
rect 149882 231548 149888 231600
rect 149940 231588 149946 231600
rect 189074 231588 189080 231600
rect 149940 231560 189080 231588
rect 149940 231548 149946 231560
rect 189074 231548 189080 231560
rect 189132 231588 189138 231600
rect 189718 231588 189724 231600
rect 189132 231560 189724 231588
rect 189132 231548 189138 231560
rect 189718 231548 189724 231560
rect 189776 231548 189782 231600
rect 215202 231548 215208 231600
rect 215260 231588 215266 231600
rect 363690 231588 363696 231600
rect 215260 231560 363696 231588
rect 215260 231548 215266 231560
rect 363690 231548 363696 231560
rect 363748 231548 363754 231600
rect 173250 231140 173256 231192
rect 173308 231180 173314 231192
rect 246298 231180 246304 231192
rect 173308 231152 246304 231180
rect 173308 231140 173314 231152
rect 246298 231140 246304 231152
rect 246356 231140 246362 231192
rect 88702 231072 88708 231124
rect 88760 231112 88766 231124
rect 315390 231112 315396 231124
rect 88760 231084 315396 231112
rect 88760 231072 88766 231084
rect 315390 231072 315396 231084
rect 315448 231072 315454 231124
rect 107378 230392 107384 230444
rect 107436 230432 107442 230444
rect 151722 230432 151728 230444
rect 107436 230404 151728 230432
rect 107436 230392 107442 230404
rect 151722 230392 151728 230404
rect 151780 230392 151786 230444
rect 169662 230392 169668 230444
rect 169720 230432 169726 230444
rect 371878 230432 371884 230444
rect 169720 230404 371884 230432
rect 169720 230392 169726 230404
rect 371878 230392 371884 230404
rect 371936 230392 371942 230444
rect 158438 230324 158444 230376
rect 158496 230364 158502 230376
rect 327718 230364 327724 230376
rect 158496 230336 327724 230364
rect 158496 230324 158502 230336
rect 327718 230324 327724 230336
rect 327776 230324 327782 230376
rect 233878 230256 233884 230308
rect 233936 230296 233942 230308
rect 353938 230296 353944 230308
rect 233936 230268 353944 230296
rect 233936 230256 233942 230268
rect 353938 230256 353944 230268
rect 353996 230256 354002 230308
rect 163590 230188 163596 230240
rect 163648 230228 163654 230240
rect 269850 230228 269856 230240
rect 163648 230200 269856 230228
rect 163648 230188 163654 230200
rect 269850 230188 269856 230200
rect 269908 230188 269914 230240
rect 166442 229848 166448 229900
rect 166500 229888 166506 229900
rect 203610 229888 203616 229900
rect 166500 229860 203616 229888
rect 166500 229848 166506 229860
rect 203610 229848 203616 229860
rect 203668 229848 203674 229900
rect 151722 229780 151728 229832
rect 151780 229820 151786 229832
rect 242158 229820 242164 229832
rect 151780 229792 242164 229820
rect 151780 229780 151786 229792
rect 242158 229780 242164 229792
rect 242216 229780 242222 229832
rect 65978 229712 65984 229764
rect 66036 229752 66042 229764
rect 380342 229752 380348 229764
rect 66036 229724 380348 229752
rect 66036 229712 66042 229724
rect 380342 229712 380348 229724
rect 380400 229752 380406 229764
rect 386414 229752 386420 229764
rect 380400 229724 386420 229752
rect 380400 229712 380406 229724
rect 386414 229712 386420 229724
rect 386472 229712 386478 229764
rect 83550 229032 83556 229084
rect 83608 229072 83614 229084
rect 130378 229072 130384 229084
rect 83608 229044 130384 229072
rect 83608 229032 83614 229044
rect 130378 229032 130384 229044
rect 130436 229032 130442 229084
rect 162670 229032 162676 229084
rect 162728 229072 162734 229084
rect 387794 229072 387800 229084
rect 162728 229044 387800 229072
rect 162728 229032 162734 229044
rect 387794 229032 387800 229044
rect 387852 229032 387858 229084
rect 60366 228964 60372 229016
rect 60424 229004 60430 229016
rect 242250 229004 242256 229016
rect 60424 228976 242256 229004
rect 60424 228964 60430 228976
rect 242250 228964 242256 228976
rect 242308 228964 242314 229016
rect 167730 228896 167736 228948
rect 167788 228936 167794 228948
rect 333238 228936 333244 228948
rect 167788 228908 333244 228936
rect 167788 228896 167794 228908
rect 333238 228896 333244 228908
rect 333296 228896 333302 228948
rect 137370 228828 137376 228880
rect 137428 228868 137434 228880
rect 223574 228868 223580 228880
rect 137428 228840 223580 228868
rect 137428 228828 137434 228840
rect 223574 228828 223580 228840
rect 223632 228868 223638 228880
rect 352558 228868 352564 228880
rect 223632 228840 352564 228868
rect 223632 228828 223638 228840
rect 352558 228828 352564 228840
rect 352616 228828 352622 228880
rect 387150 228692 387156 228744
rect 387208 228732 387214 228744
rect 387702 228732 387708 228744
rect 387208 228704 387708 228732
rect 387208 228692 387214 228704
rect 387702 228692 387708 228704
rect 387760 228692 387766 228744
rect 387794 228420 387800 228472
rect 387852 228460 387858 228472
rect 388438 228460 388444 228472
rect 387852 228432 388444 228460
rect 387852 228420 387858 228432
rect 388438 228420 388444 228432
rect 388496 228420 388502 228472
rect 7558 228352 7564 228404
rect 7616 228392 7622 228404
rect 83550 228392 83556 228404
rect 7616 228364 83556 228392
rect 7616 228352 7622 228364
rect 83550 228352 83556 228364
rect 83608 228352 83614 228404
rect 332686 228284 332692 228336
rect 332744 228324 332750 228336
rect 333238 228324 333244 228336
rect 332744 228296 333244 228324
rect 332744 228284 332750 228296
rect 333238 228284 333244 228296
rect 333296 228284 333302 228336
rect 52362 227672 52368 227724
rect 52420 227712 52426 227724
rect 345014 227712 345020 227724
rect 52420 227684 345020 227712
rect 52420 227672 52426 227684
rect 345014 227672 345020 227684
rect 345072 227712 345078 227724
rect 345750 227712 345756 227724
rect 345072 227684 345756 227712
rect 345072 227672 345078 227684
rect 345750 227672 345756 227684
rect 345808 227672 345814 227724
rect 160738 227604 160744 227656
rect 160796 227644 160802 227656
rect 318150 227644 318156 227656
rect 160796 227616 318156 227644
rect 160796 227604 160802 227616
rect 318150 227604 318156 227616
rect 318208 227604 318214 227656
rect 572622 227332 572628 227384
rect 572680 227372 572686 227384
rect 576854 227372 576860 227384
rect 572680 227344 576860 227372
rect 572680 227332 572686 227344
rect 576854 227332 576860 227344
rect 576912 227332 576918 227384
rect 177666 227264 177672 227316
rect 177724 227304 177730 227316
rect 196618 227304 196624 227316
rect 177724 227276 196624 227304
rect 177724 227264 177730 227276
rect 196618 227264 196624 227276
rect 196676 227264 196682 227316
rect 61746 227196 61752 227248
rect 61804 227236 61810 227248
rect 197998 227236 198004 227248
rect 61804 227208 198004 227236
rect 61804 227196 61810 227208
rect 197998 227196 198004 227208
rect 198056 227196 198062 227248
rect 195974 227128 195980 227180
rect 196032 227168 196038 227180
rect 353938 227168 353944 227180
rect 196032 227140 353944 227168
rect 196032 227128 196038 227140
rect 353938 227128 353944 227140
rect 353996 227128 354002 227180
rect 48130 227060 48136 227112
rect 48188 227100 48194 227112
rect 269758 227100 269764 227112
rect 48188 227072 269764 227100
rect 48188 227060 48194 227072
rect 269758 227060 269764 227072
rect 269816 227060 269822 227112
rect 67358 226992 67364 227044
rect 67416 227032 67422 227044
rect 386966 227032 386972 227044
rect 67416 227004 386972 227032
rect 67416 226992 67422 227004
rect 386966 226992 386972 227004
rect 387024 226992 387030 227044
rect 48222 226244 48228 226296
rect 48280 226284 48286 226296
rect 361022 226284 361028 226296
rect 48280 226256 361028 226284
rect 48280 226244 48286 226256
rect 361022 226244 361028 226256
rect 361080 226244 361086 226296
rect 133322 226176 133328 226228
rect 133380 226216 133386 226228
rect 378870 226216 378876 226228
rect 133380 226188 378876 226216
rect 133380 226176 133386 226188
rect 378870 226176 378876 226188
rect 378928 226176 378934 226228
rect 158530 226108 158536 226160
rect 158588 226148 158594 226160
rect 342898 226148 342904 226160
rect 158588 226120 342904 226148
rect 158588 226108 158594 226120
rect 342898 226108 342904 226120
rect 342956 226108 342962 226160
rect 54846 225632 54852 225684
rect 54904 225672 54910 225684
rect 160738 225672 160744 225684
rect 54904 225644 160744 225672
rect 54904 225632 54910 225644
rect 160738 225632 160744 225644
rect 160796 225632 160802 225684
rect 170582 225632 170588 225684
rect 170640 225672 170646 225684
rect 243538 225672 243544 225684
rect 170640 225644 243544 225672
rect 170640 225632 170646 225644
rect 243538 225632 243544 225644
rect 243596 225632 243602 225684
rect 271874 225632 271880 225684
rect 271932 225672 271938 225684
rect 294138 225672 294144 225684
rect 271932 225644 294144 225672
rect 271932 225632 271938 225644
rect 294138 225632 294144 225644
rect 294196 225632 294202 225684
rect 100294 225564 100300 225616
rect 100352 225604 100358 225616
rect 222838 225604 222844 225616
rect 100352 225576 222844 225604
rect 100352 225564 100358 225576
rect 222838 225564 222844 225576
rect 222896 225564 222902 225616
rect 256694 225564 256700 225616
rect 256752 225604 256758 225616
rect 268378 225604 268384 225616
rect 256752 225576 268384 225604
rect 256752 225564 256758 225576
rect 268378 225564 268384 225576
rect 268436 225564 268442 225616
rect 291838 225564 291844 225616
rect 291896 225604 291902 225616
rect 316034 225604 316040 225616
rect 291896 225576 316040 225604
rect 291896 225564 291902 225576
rect 316034 225564 316040 225576
rect 316092 225564 316098 225616
rect 360286 225428 360292 225480
rect 360344 225468 360350 225480
rect 361022 225468 361028 225480
rect 360344 225440 361028 225468
rect 360344 225428 360350 225440
rect 361022 225428 361028 225440
rect 361080 225428 361086 225480
rect 378134 225156 378140 225208
rect 378192 225196 378198 225208
rect 378870 225196 378876 225208
rect 378192 225168 378876 225196
rect 378192 225156 378198 225168
rect 378870 225156 378876 225168
rect 378928 225156 378934 225208
rect 149974 224884 149980 224936
rect 150032 224924 150038 224936
rect 360194 224924 360200 224936
rect 150032 224896 360200 224924
rect 150032 224884 150038 224896
rect 360194 224884 360200 224896
rect 360252 224884 360258 224936
rect 148502 224816 148508 224868
rect 148560 224856 148566 224868
rect 276014 224856 276020 224868
rect 148560 224828 276020 224856
rect 148560 224816 148566 224828
rect 276014 224816 276020 224828
rect 276072 224816 276078 224868
rect 347130 224816 347136 224868
rect 347188 224856 347194 224868
rect 347774 224856 347780 224868
rect 347188 224828 347780 224856
rect 347188 224816 347194 224828
rect 347774 224816 347780 224828
rect 347832 224816 347838 224868
rect 360194 224476 360200 224528
rect 360252 224516 360258 224528
rect 360838 224516 360844 224528
rect 360252 224488 360844 224516
rect 360252 224476 360258 224488
rect 360838 224476 360844 224488
rect 360896 224476 360902 224528
rect 276014 224408 276020 224460
rect 276072 224448 276078 224460
rect 276658 224448 276664 224460
rect 276072 224420 276664 224448
rect 276072 224408 276078 224420
rect 276658 224408 276664 224420
rect 276716 224408 276722 224460
rect 59078 223524 59084 223576
rect 59136 223564 59142 223576
rect 327166 223564 327172 223576
rect 59136 223536 327172 223564
rect 59136 223524 59142 223536
rect 327166 223524 327172 223536
rect 327224 223564 327230 223576
rect 327810 223564 327816 223576
rect 327224 223536 327816 223564
rect 327224 223524 327230 223536
rect 327810 223524 327816 223536
rect 327868 223524 327874 223576
rect 385126 223564 385132 223576
rect 373966 223536 385132 223564
rect 153838 223456 153844 223508
rect 153896 223496 153902 223508
rect 373966 223496 373994 223536
rect 385126 223524 385132 223536
rect 385184 223564 385190 223576
rect 385862 223564 385868 223576
rect 385184 223536 385868 223564
rect 385184 223524 385190 223536
rect 385862 223524 385868 223536
rect 385920 223524 385926 223576
rect 153896 223468 373994 223496
rect 153896 223456 153902 223468
rect 145742 223388 145748 223440
rect 145800 223428 145806 223440
rect 298186 223428 298192 223440
rect 145800 223400 298192 223428
rect 145800 223388 145806 223400
rect 298186 223388 298192 223400
rect 298244 223388 298250 223440
rect 125134 222912 125140 222964
rect 125192 222952 125198 222964
rect 220078 222952 220084 222964
rect 125192 222924 220084 222952
rect 125192 222912 125198 222924
rect 220078 222912 220084 222924
rect 220136 222912 220142 222964
rect 56410 222844 56416 222896
rect 56468 222884 56474 222896
rect 117958 222884 117964 222896
rect 56468 222856 117964 222884
rect 56468 222844 56474 222856
rect 117958 222844 117964 222856
rect 118016 222844 118022 222896
rect 165154 222844 165160 222896
rect 165212 222884 165218 222896
rect 278130 222884 278136 222896
rect 165212 222856 278136 222884
rect 165212 222844 165218 222856
rect 278130 222844 278136 222856
rect 278188 222844 278194 222896
rect 45370 222096 45376 222148
rect 45428 222136 45434 222148
rect 342346 222136 342352 222148
rect 45428 222108 342352 222136
rect 45428 222096 45434 222108
rect 342346 222096 342352 222108
rect 342404 222136 342410 222148
rect 342990 222136 342996 222148
rect 342404 222108 342996 222136
rect 342404 222096 342410 222108
rect 342990 222096 342996 222108
rect 343048 222096 343054 222148
rect 162302 222028 162308 222080
rect 162360 222068 162366 222080
rect 263594 222068 263600 222080
rect 162360 222040 263600 222068
rect 162360 222028 162366 222040
rect 263594 222028 263600 222040
rect 263652 222068 263658 222080
rect 264238 222068 264244 222080
rect 263652 222040 264244 222068
rect 263652 222028 263658 222040
rect 264238 222028 264244 222040
rect 264296 222028 264302 222080
rect 310422 222028 310428 222080
rect 310480 222068 310486 222080
rect 314010 222068 314016 222080
rect 310480 222040 314016 222068
rect 310480 222028 310486 222040
rect 314010 222028 314016 222040
rect 314068 222028 314074 222080
rect 141418 221620 141424 221672
rect 141476 221660 141482 221672
rect 211890 221660 211896 221672
rect 141476 221632 211896 221660
rect 141476 221620 141482 221632
rect 211890 221620 211896 221632
rect 211948 221620 211954 221672
rect 131850 221552 131856 221604
rect 131908 221592 131914 221604
rect 247678 221592 247684 221604
rect 131908 221564 247684 221592
rect 131908 221552 131914 221564
rect 247678 221552 247684 221564
rect 247736 221552 247742 221604
rect 87414 221484 87420 221536
rect 87472 221524 87478 221536
rect 207658 221524 207664 221536
rect 87472 221496 207664 221524
rect 87472 221484 87478 221496
rect 207658 221484 207664 221496
rect 207716 221484 207722 221536
rect 3418 221416 3424 221468
rect 3476 221456 3482 221468
rect 120166 221456 120172 221468
rect 3476 221428 120172 221456
rect 3476 221416 3482 221428
rect 120166 221416 120172 221428
rect 120224 221416 120230 221468
rect 151170 221416 151176 221468
rect 151228 221456 151234 221468
rect 310422 221456 310428 221468
rect 151228 221428 310428 221456
rect 151228 221416 151234 221428
rect 310422 221416 310428 221428
rect 310480 221416 310486 221468
rect 144454 220736 144460 220788
rect 144512 220776 144518 220788
rect 386874 220776 386880 220788
rect 144512 220748 386880 220776
rect 144512 220736 144518 220748
rect 386874 220736 386880 220748
rect 386932 220736 386938 220788
rect 156690 220668 156696 220720
rect 156748 220708 156754 220720
rect 385034 220708 385040 220720
rect 156748 220680 385040 220708
rect 156748 220668 156754 220680
rect 385034 220668 385040 220680
rect 385092 220708 385098 220720
rect 385770 220708 385776 220720
rect 385092 220680 385776 220708
rect 385092 220668 385098 220680
rect 385770 220668 385776 220680
rect 385828 220668 385834 220720
rect 102870 220192 102876 220244
rect 102928 220232 102934 220244
rect 252738 220232 252744 220244
rect 102928 220204 252744 220232
rect 102928 220192 102934 220204
rect 252738 220192 252744 220204
rect 252796 220192 252802 220244
rect 69198 220124 69204 220176
rect 69256 220164 69262 220176
rect 251174 220164 251180 220176
rect 69256 220136 251180 220164
rect 69256 220124 69262 220136
rect 251174 220124 251180 220136
rect 251232 220124 251238 220176
rect 50890 220056 50896 220108
rect 50948 220096 50954 220108
rect 356054 220096 356060 220108
rect 50948 220068 356060 220096
rect 50948 220056 50954 220068
rect 356054 220056 356060 220068
rect 356112 220056 356118 220108
rect 153930 219376 153936 219428
rect 153988 219416 153994 219428
rect 363782 219416 363788 219428
rect 153988 219388 363788 219416
rect 153988 219376 153994 219388
rect 363782 219376 363788 219388
rect 363840 219376 363846 219428
rect 576210 219376 576216 219428
rect 576268 219416 576274 219428
rect 580074 219416 580080 219428
rect 576268 219388 580080 219416
rect 576268 219376 576274 219388
rect 580074 219376 580080 219388
rect 580132 219376 580138 219428
rect 155862 219308 155868 219360
rect 155920 219348 155926 219360
rect 360930 219348 360936 219360
rect 155920 219320 360936 219348
rect 155920 219308 155926 219320
rect 360930 219308 360936 219320
rect 360988 219308 360994 219360
rect 57698 218832 57704 218884
rect 57756 218872 57762 218884
rect 162762 218872 162768 218884
rect 57756 218844 162768 218872
rect 57756 218832 57762 218844
rect 162762 218832 162768 218844
rect 162820 218832 162826 218884
rect 53650 218764 53656 218816
rect 53708 218804 53714 218816
rect 153838 218804 153844 218816
rect 53708 218776 153844 218804
rect 53708 218764 53714 218776
rect 153838 218764 153844 218776
rect 153896 218764 153902 218816
rect 160738 218764 160744 218816
rect 160796 218804 160802 218816
rect 274634 218804 274640 218816
rect 160796 218776 274640 218804
rect 160796 218764 160802 218776
rect 274634 218764 274640 218776
rect 274692 218764 274698 218816
rect 137462 218696 137468 218748
rect 137520 218736 137526 218748
rect 338206 218736 338212 218748
rect 137520 218708 338212 218736
rect 137520 218696 137526 218708
rect 338206 218696 338212 218708
rect 338264 218696 338270 218748
rect 153102 217948 153108 218000
rect 153160 217988 153166 218000
rect 270494 217988 270500 218000
rect 153160 217960 270500 217988
rect 153160 217948 153166 217960
rect 270494 217948 270500 217960
rect 270552 217948 270558 218000
rect 114554 217472 114560 217524
rect 114612 217512 114618 217524
rect 289078 217512 289084 217524
rect 114612 217484 289084 217512
rect 114612 217472 114618 217484
rect 289078 217472 289084 217484
rect 289136 217472 289142 217524
rect 77386 217404 77392 217456
rect 77444 217444 77450 217456
rect 252830 217444 252836 217456
rect 77444 217416 252836 217444
rect 77444 217404 77450 217416
rect 252830 217404 252836 217416
rect 252888 217404 252894 217456
rect 280890 217404 280896 217456
rect 280948 217444 280954 217456
rect 311894 217444 311900 217456
rect 280948 217416 311900 217444
rect 280948 217404 280954 217416
rect 311894 217404 311900 217416
rect 311952 217404 311958 217456
rect 52270 217336 52276 217388
rect 52328 217376 52334 217388
rect 233878 217376 233884 217388
rect 52328 217348 233884 217376
rect 52328 217336 52334 217348
rect 233878 217336 233884 217348
rect 233936 217336 233942 217388
rect 248414 217336 248420 217388
rect 248472 217376 248478 217388
rect 291194 217376 291200 217388
rect 248472 217348 291200 217376
rect 248472 217336 248478 217348
rect 291194 217336 291200 217348
rect 291252 217336 291258 217388
rect 169018 217268 169024 217320
rect 169076 217308 169082 217320
rect 357986 217308 357992 217320
rect 169076 217280 357992 217308
rect 169076 217268 169082 217280
rect 357986 217268 357992 217280
rect 358044 217268 358050 217320
rect 270494 216656 270500 216708
rect 270552 216696 270558 216708
rect 271230 216696 271236 216708
rect 270552 216668 271236 216696
rect 270552 216656 270558 216668
rect 271230 216656 271236 216668
rect 271288 216656 271294 216708
rect 242158 216588 242164 216640
rect 242216 216628 242222 216640
rect 387518 216628 387524 216640
rect 242216 216600 387524 216628
rect 242216 216588 242222 216600
rect 387518 216588 387524 216600
rect 387576 216588 387582 216640
rect 357986 216520 357992 216572
rect 358044 216560 358050 216572
rect 358170 216560 358176 216572
rect 358044 216532 358176 216560
rect 358044 216520 358050 216532
rect 358170 216520 358176 216532
rect 358228 216560 358234 216572
rect 373258 216560 373264 216572
rect 358228 216532 373264 216560
rect 358228 216520 358234 216532
rect 373258 216520 373264 216532
rect 373316 216520 373322 216572
rect 141602 216112 141608 216164
rect 141660 216152 141666 216164
rect 261478 216152 261484 216164
rect 141660 216124 261484 216152
rect 141660 216112 141666 216124
rect 261478 216112 261484 216124
rect 261536 216112 261542 216164
rect 104986 216044 104992 216096
rect 105044 216084 105050 216096
rect 283650 216084 283656 216096
rect 105044 216056 283656 216084
rect 105044 216044 105050 216056
rect 283650 216044 283656 216056
rect 283708 216044 283714 216096
rect 70394 215976 70400 216028
rect 70452 216016 70458 216028
rect 249794 216016 249800 216028
rect 70452 215988 249800 216016
rect 70452 215976 70458 215988
rect 249794 215976 249800 215988
rect 249852 215976 249858 216028
rect 92566 215908 92572 215960
rect 92624 215948 92630 215960
rect 314010 215948 314016 215960
rect 92624 215920 314016 215948
rect 92624 215908 92630 215920
rect 314010 215908 314016 215920
rect 314068 215908 314074 215960
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 21358 215268 21364 215280
rect 3384 215240 21364 215268
rect 3384 215228 3390 215240
rect 21358 215228 21364 215240
rect 21416 215228 21422 215280
rect 162762 215228 162768 215280
rect 162820 215268 162826 215280
rect 287698 215268 287704 215280
rect 162820 215240 287704 215268
rect 162820 215228 162826 215240
rect 287698 215228 287704 215240
rect 287756 215228 287762 215280
rect 155218 214752 155224 214804
rect 155276 214792 155282 214804
rect 256694 214792 256700 214804
rect 155276 214764 256700 214792
rect 155276 214752 155282 214764
rect 256694 214752 256700 214764
rect 256752 214752 256758 214804
rect 100846 214684 100852 214736
rect 100904 214724 100910 214736
rect 263594 214724 263600 214736
rect 100904 214696 263600 214724
rect 100904 214684 100910 214696
rect 263594 214684 263600 214696
rect 263652 214684 263658 214736
rect 325050 214684 325056 214736
rect 325108 214724 325114 214736
rect 349154 214724 349160 214736
rect 325108 214696 349160 214724
rect 325108 214684 325114 214696
rect 349154 214684 349160 214696
rect 349212 214684 349218 214736
rect 96706 214616 96712 214668
rect 96764 214656 96770 214668
rect 336734 214656 336740 214668
rect 96764 214628 336740 214656
rect 96764 214616 96770 214628
rect 336734 214616 336740 214628
rect 336792 214616 336798 214668
rect 76558 214548 76564 214600
rect 76616 214588 76622 214600
rect 330478 214588 330484 214600
rect 76616 214560 330484 214588
rect 76616 214548 76622 214560
rect 330478 214548 330484 214560
rect 330536 214548 330542 214600
rect 64690 213868 64696 213920
rect 64748 213908 64754 213920
rect 331306 213908 331312 213920
rect 64748 213880 331312 213908
rect 64748 213868 64754 213880
rect 331306 213868 331312 213880
rect 331364 213908 331370 213920
rect 331950 213908 331956 213920
rect 331364 213880 331956 213908
rect 331364 213868 331370 213880
rect 331950 213868 331956 213880
rect 332008 213868 332014 213920
rect 130562 213324 130568 213376
rect 130620 213364 130626 213376
rect 191098 213364 191104 213376
rect 130620 213336 191104 213364
rect 130620 213324 130626 213336
rect 191098 213324 191104 213336
rect 191156 213324 191162 213376
rect 202138 213324 202144 213376
rect 202196 213364 202202 213376
rect 283558 213364 283564 213376
rect 202196 213336 283564 213364
rect 202196 213324 202202 213336
rect 283558 213324 283564 213336
rect 283616 213324 283622 213376
rect 127710 213256 127716 213308
rect 127768 213296 127774 213308
rect 270494 213296 270500 213308
rect 127768 213268 270500 213296
rect 127768 213256 127774 213268
rect 270494 213256 270500 213268
rect 270552 213256 270558 213308
rect 60458 213188 60464 213240
rect 60516 213228 60522 213240
rect 238018 213228 238024 213240
rect 60516 213200 238024 213228
rect 60516 213188 60522 213200
rect 238018 213188 238024 213200
rect 238076 213188 238082 213240
rect 273990 213188 273996 213240
rect 274048 213228 274054 213240
rect 346394 213228 346400 213240
rect 274048 213200 346400 213228
rect 274048 213188 274054 213200
rect 346394 213188 346400 213200
rect 346452 213228 346458 213240
rect 347682 213228 347688 213240
rect 346452 213200 347688 213228
rect 346452 213188 346458 213200
rect 347682 213188 347688 213200
rect 347740 213188 347746 213240
rect 347682 212508 347688 212560
rect 347740 212548 347746 212560
rect 386874 212548 386880 212560
rect 347740 212520 386880 212548
rect 347740 212508 347746 212520
rect 386874 212508 386880 212520
rect 386932 212508 386938 212560
rect 572622 212508 572628 212560
rect 572680 212548 572686 212560
rect 582742 212548 582748 212560
rect 572680 212520 582748 212548
rect 572680 212508 572686 212520
rect 582742 212508 582748 212520
rect 582800 212508 582806 212560
rect 148594 211964 148600 212016
rect 148652 212004 148658 212016
rect 242158 212004 242164 212016
rect 148652 211976 242164 212004
rect 148652 211964 148658 211976
rect 242158 211964 242164 211976
rect 242216 211964 242222 212016
rect 111794 211896 111800 211948
rect 111852 211936 111858 211948
rect 273254 211936 273260 211948
rect 111852 211908 273260 211936
rect 111852 211896 111858 211908
rect 273254 211896 273260 211908
rect 273312 211896 273318 211948
rect 92474 211828 92480 211880
rect 92532 211868 92538 211880
rect 259546 211868 259552 211880
rect 92532 211840 259552 211868
rect 92532 211828 92538 211840
rect 259546 211828 259552 211840
rect 259604 211828 259610 211880
rect 88978 211760 88984 211812
rect 89036 211800 89042 211812
rect 312538 211800 312544 211812
rect 89036 211772 312544 211800
rect 89036 211760 89042 211772
rect 312538 211760 312544 211772
rect 312596 211760 312602 211812
rect 323578 211760 323584 211812
rect 323636 211800 323642 211812
rect 340966 211800 340972 211812
rect 323636 211772 340972 211800
rect 323636 211760 323642 211772
rect 340966 211760 340972 211772
rect 341024 211760 341030 211812
rect 344278 211760 344284 211812
rect 344336 211800 344342 211812
rect 387150 211800 387156 211812
rect 344336 211772 387156 211800
rect 344336 211760 344342 211772
rect 387150 211760 387156 211772
rect 387208 211760 387214 211812
rect 572622 211080 572628 211132
rect 572680 211120 572686 211132
rect 583570 211120 583576 211132
rect 572680 211092 583576 211120
rect 572680 211080 572686 211092
rect 583570 211080 583576 211092
rect 583628 211080 583634 211132
rect 142890 210672 142896 210724
rect 142948 210712 142954 210724
rect 229738 210712 229744 210724
rect 142948 210684 229744 210712
rect 142948 210672 142954 210684
rect 229738 210672 229744 210684
rect 229796 210672 229802 210724
rect 95878 210604 95884 210656
rect 95936 210644 95942 210656
rect 166166 210644 166172 210656
rect 95936 210616 166172 210644
rect 95936 210604 95942 210616
rect 166166 210604 166172 210616
rect 166224 210604 166230 210656
rect 203518 210604 203524 210656
rect 203576 210644 203582 210656
rect 340138 210644 340144 210656
rect 203576 210616 340144 210644
rect 203576 210604 203582 210616
rect 340138 210604 340144 210616
rect 340196 210604 340202 210656
rect 137278 210536 137284 210588
rect 137336 210576 137342 210588
rect 277394 210576 277400 210588
rect 137336 210548 277400 210576
rect 137336 210536 137342 210548
rect 277394 210536 277400 210548
rect 277452 210536 277458 210588
rect 103606 210468 103612 210520
rect 103664 210508 103670 210520
rect 352558 210508 352564 210520
rect 103664 210480 352564 210508
rect 103664 210468 103670 210480
rect 352558 210468 352564 210480
rect 352616 210468 352622 210520
rect 78674 210400 78680 210452
rect 78732 210440 78738 210452
rect 329834 210440 329840 210452
rect 78732 210412 329840 210440
rect 78732 210400 78738 210412
rect 329834 210400 329840 210412
rect 329892 210400 329898 210452
rect 80146 209380 80152 209432
rect 80204 209420 80210 209432
rect 162302 209420 162308 209432
rect 80204 209392 162308 209420
rect 80204 209380 80210 209392
rect 162302 209380 162308 209392
rect 162360 209380 162366 209432
rect 144178 209312 144184 209364
rect 144236 209352 144242 209364
rect 280154 209352 280160 209364
rect 144236 209324 280160 209352
rect 144236 209312 144242 209324
rect 280154 209312 280160 209324
rect 280212 209312 280218 209364
rect 86218 209244 86224 209296
rect 86276 209284 86282 209296
rect 240778 209284 240784 209296
rect 86276 209256 240784 209284
rect 86276 209244 86282 209256
rect 240778 209244 240784 209256
rect 240836 209244 240842 209296
rect 136082 209176 136088 209228
rect 136140 209216 136146 209228
rect 327074 209216 327080 209228
rect 136140 209188 327080 209216
rect 136140 209176 136146 209188
rect 327074 209176 327080 209188
rect 327132 209216 327138 209228
rect 327902 209216 327908 209228
rect 327132 209188 327908 209216
rect 327132 209176 327138 209188
rect 327902 209176 327908 209188
rect 327960 209176 327966 209228
rect 49510 209108 49516 209160
rect 49568 209148 49574 209160
rect 269298 209148 269304 209160
rect 49568 209120 269304 209148
rect 49568 209108 49574 209120
rect 269298 209108 269304 209120
rect 269356 209108 269362 209160
rect 107746 209040 107752 209092
rect 107804 209080 107810 209092
rect 335538 209080 335544 209092
rect 107804 209052 335544 209080
rect 107804 209040 107810 209052
rect 335538 209040 335544 209052
rect 335596 209040 335602 209092
rect 327902 208360 327908 208412
rect 327960 208400 327966 208412
rect 386874 208400 386880 208412
rect 327960 208372 386880 208400
rect 327960 208360 327966 208372
rect 386874 208360 386880 208372
rect 386932 208360 386938 208412
rect 149698 207816 149704 207868
rect 149756 207856 149762 207868
rect 259454 207856 259460 207868
rect 149756 207828 259460 207856
rect 149756 207816 149762 207828
rect 259454 207816 259460 207828
rect 259512 207816 259518 207868
rect 86954 207748 86960 207800
rect 87012 207788 87018 207800
rect 252646 207788 252652 207800
rect 87012 207760 252652 207788
rect 87012 207748 87018 207760
rect 252646 207748 252652 207760
rect 252704 207748 252710 207800
rect 84378 207680 84384 207732
rect 84436 207720 84442 207732
rect 267734 207720 267740 207732
rect 84436 207692 267740 207720
rect 84436 207680 84442 207692
rect 267734 207680 267740 207692
rect 267792 207680 267798 207732
rect 60550 207612 60556 207664
rect 60608 207652 60614 207664
rect 336826 207652 336832 207664
rect 60608 207624 336832 207652
rect 60608 207612 60614 207624
rect 336826 207612 336832 207624
rect 336884 207612 336890 207664
rect 572438 206932 572444 206984
rect 572496 206972 572502 206984
rect 575474 206972 575480 206984
rect 572496 206944 575480 206972
rect 572496 206932 572502 206944
rect 575474 206932 575480 206944
rect 575532 206932 575538 206984
rect 143074 206524 143080 206576
rect 143132 206564 143138 206576
rect 265066 206564 265072 206576
rect 143132 206536 265072 206564
rect 143132 206524 143138 206536
rect 265066 206524 265072 206536
rect 265124 206524 265130 206576
rect 89806 206456 89812 206508
rect 89864 206496 89870 206508
rect 249886 206496 249892 206508
rect 89864 206468 249892 206496
rect 89864 206456 89870 206468
rect 249886 206456 249892 206468
rect 249944 206456 249950 206508
rect 65886 206388 65892 206440
rect 65944 206428 65950 206440
rect 255406 206428 255412 206440
rect 65944 206400 255412 206428
rect 65944 206388 65950 206400
rect 255406 206388 255412 206400
rect 255464 206388 255470 206440
rect 281534 206388 281540 206440
rect 281592 206428 281598 206440
rect 342254 206428 342260 206440
rect 281592 206400 342260 206428
rect 281592 206388 281598 206400
rect 342254 206388 342260 206400
rect 342312 206388 342318 206440
rect 118694 206320 118700 206372
rect 118752 206360 118758 206372
rect 315482 206360 315488 206372
rect 118752 206332 315488 206360
rect 118752 206320 118758 206332
rect 315482 206320 315488 206332
rect 315540 206320 315546 206372
rect 57882 206252 57888 206304
rect 57940 206292 57946 206304
rect 300210 206292 300216 206304
rect 57940 206264 300216 206292
rect 57940 206252 57946 206264
rect 300210 206252 300216 206264
rect 300268 206252 300274 206304
rect 351270 205640 351276 205692
rect 351328 205680 351334 205692
rect 386874 205680 386880 205692
rect 351328 205652 386880 205680
rect 351328 205640 351334 205652
rect 386874 205640 386880 205652
rect 386932 205640 386938 205692
rect 576210 205640 576216 205692
rect 576268 205680 576274 205692
rect 580902 205680 580908 205692
rect 576268 205652 580908 205680
rect 576268 205640 576274 205652
rect 580902 205640 580908 205652
rect 580960 205640 580966 205692
rect 162118 205164 162124 205216
rect 162176 205204 162182 205216
rect 225598 205204 225604 205216
rect 162176 205176 225604 205204
rect 162176 205164 162182 205176
rect 225598 205164 225604 205176
rect 225656 205164 225662 205216
rect 107654 205096 107660 205148
rect 107712 205136 107718 205148
rect 167730 205136 167736 205148
rect 107712 205108 167736 205136
rect 107712 205096 107718 205108
rect 167730 205096 167736 205108
rect 167788 205096 167794 205148
rect 224954 205096 224960 205148
rect 225012 205136 225018 205148
rect 308490 205136 308496 205148
rect 225012 205108 308496 205136
rect 225012 205096 225018 205108
rect 308490 205096 308496 205108
rect 308548 205096 308554 205148
rect 166166 205028 166172 205080
rect 166224 205068 166230 205080
rect 281534 205068 281540 205080
rect 166224 205040 281540 205068
rect 166224 205028 166230 205040
rect 281534 205028 281540 205040
rect 281592 205028 281598 205080
rect 53742 204960 53748 205012
rect 53800 205000 53806 205012
rect 238110 205000 238116 205012
rect 53800 204972 238116 205000
rect 53800 204960 53806 204972
rect 238110 204960 238116 204972
rect 238168 204960 238174 205012
rect 134702 204892 134708 204944
rect 134760 204932 134766 204944
rect 340138 204932 340144 204944
rect 134760 204904 340144 204932
rect 134760 204892 134766 204904
rect 340138 204892 340144 204904
rect 340196 204892 340202 204944
rect 571518 203872 571524 203924
rect 571576 203912 571582 203924
rect 574278 203912 574284 203924
rect 571576 203884 574284 203912
rect 571576 203872 571582 203884
rect 574278 203872 574284 203884
rect 574336 203872 574342 203924
rect 145558 203736 145564 203788
rect 145616 203776 145622 203788
rect 235258 203776 235264 203788
rect 145616 203748 235264 203776
rect 145616 203736 145622 203748
rect 235258 203736 235264 203748
rect 235316 203736 235322 203788
rect 73246 203668 73252 203720
rect 73304 203708 73310 203720
rect 148410 203708 148416 203720
rect 73304 203680 148416 203708
rect 73304 203668 73310 203680
rect 148410 203668 148416 203680
rect 148468 203668 148474 203720
rect 149790 203668 149796 203720
rect 149848 203708 149854 203720
rect 278774 203708 278780 203720
rect 149848 203680 278780 203708
rect 149848 203668 149854 203680
rect 278774 203668 278780 203680
rect 278832 203668 278838 203720
rect 315298 203668 315304 203720
rect 315356 203708 315362 203720
rect 360838 203708 360844 203720
rect 315356 203680 360844 203708
rect 315356 203668 315362 203680
rect 360838 203668 360844 203680
rect 360896 203668 360902 203720
rect 129182 203600 129188 203652
rect 129240 203640 129246 203652
rect 347866 203640 347872 203652
rect 129240 203612 347872 203640
rect 129240 203600 129246 203612
rect 347866 203600 347872 203612
rect 347924 203600 347930 203652
rect 69014 203532 69020 203584
rect 69072 203572 69078 203584
rect 324314 203572 324320 203584
rect 69072 203544 324320 203572
rect 69072 203532 69078 203544
rect 324314 203532 324320 203544
rect 324372 203532 324378 203584
rect 147030 202376 147036 202428
rect 147088 202416 147094 202428
rect 239398 202416 239404 202428
rect 147088 202388 239404 202416
rect 147088 202376 147094 202388
rect 239398 202376 239404 202388
rect 239456 202376 239462 202428
rect 129090 202308 129096 202360
rect 129148 202348 129154 202360
rect 232498 202348 232504 202360
rect 129148 202320 232504 202348
rect 129148 202308 129154 202320
rect 232498 202308 232504 202320
rect 232556 202308 232562 202360
rect 245654 202308 245660 202360
rect 245712 202348 245718 202360
rect 309870 202348 309876 202360
rect 245712 202320 309876 202348
rect 245712 202308 245718 202320
rect 309870 202308 309876 202320
rect 309928 202308 309934 202360
rect 126330 202240 126336 202292
rect 126388 202280 126394 202292
rect 264974 202280 264980 202292
rect 126388 202252 264980 202280
rect 126388 202240 126394 202252
rect 264974 202240 264980 202252
rect 265032 202240 265038 202292
rect 110506 202172 110512 202224
rect 110564 202212 110570 202224
rect 255590 202212 255596 202224
rect 110564 202184 255596 202212
rect 110564 202172 110570 202184
rect 255590 202172 255596 202184
rect 255648 202172 255654 202224
rect 340138 202172 340144 202224
rect 340196 202212 340202 202224
rect 386874 202212 386880 202224
rect 340196 202184 386880 202212
rect 340196 202172 340202 202184
rect 386874 202172 386880 202184
rect 386932 202172 386938 202224
rect 159358 202104 159364 202156
rect 159416 202144 159422 202156
rect 347958 202144 347964 202156
rect 159416 202116 347964 202144
rect 159416 202104 159422 202116
rect 347958 202104 347964 202116
rect 348016 202104 348022 202156
rect 96614 200948 96620 201000
rect 96672 200988 96678 201000
rect 160094 200988 160100 201000
rect 96672 200960 160100 200988
rect 96672 200948 96678 200960
rect 160094 200948 160100 200960
rect 160152 200948 160158 201000
rect 136174 200880 136180 200932
rect 136232 200920 136238 200932
rect 262306 200920 262312 200932
rect 136232 200892 262312 200920
rect 136232 200880 136238 200892
rect 262306 200880 262312 200892
rect 262364 200880 262370 200932
rect 140222 200812 140228 200864
rect 140280 200852 140286 200864
rect 269206 200852 269212 200864
rect 140280 200824 269212 200852
rect 140280 200812 140286 200824
rect 269206 200812 269212 200824
rect 269264 200812 269270 200864
rect 103698 200744 103704 200796
rect 103756 200784 103762 200796
rect 322934 200784 322940 200796
rect 103756 200756 322940 200784
rect 103756 200744 103762 200756
rect 322934 200744 322940 200756
rect 322992 200744 322998 200796
rect 100754 199588 100760 199640
rect 100812 199628 100818 199640
rect 255498 199628 255504 199640
rect 100812 199600 255504 199628
rect 100812 199588 100818 199600
rect 255498 199588 255504 199600
rect 255556 199588 255562 199640
rect 318058 199588 318064 199640
rect 318116 199628 318122 199640
rect 335446 199628 335452 199640
rect 318116 199600 335452 199628
rect 318116 199588 318122 199600
rect 335446 199588 335452 199600
rect 335504 199588 335510 199640
rect 162210 199520 162216 199572
rect 162268 199560 162274 199572
rect 318150 199560 318156 199572
rect 162268 199532 318156 199560
rect 162268 199520 162274 199532
rect 318150 199520 318156 199532
rect 318208 199520 318214 199572
rect 116578 199452 116584 199504
rect 116636 199492 116642 199504
rect 333238 199492 333244 199504
rect 116636 199464 333244 199492
rect 116636 199452 116642 199464
rect 333238 199452 333244 199464
rect 333296 199452 333302 199504
rect 120718 199384 120724 199436
rect 120776 199424 120782 199436
rect 340230 199424 340236 199436
rect 120776 199396 340236 199424
rect 120776 199384 120782 199396
rect 340230 199384 340236 199396
rect 340288 199384 340294 199436
rect 572622 198636 572628 198688
rect 572680 198676 572686 198688
rect 579706 198676 579712 198688
rect 572680 198648 579712 198676
rect 572680 198636 572686 198648
rect 579706 198636 579712 198648
rect 579764 198636 579770 198688
rect 151078 198228 151084 198280
rect 151136 198268 151142 198280
rect 233970 198268 233976 198280
rect 151136 198240 233976 198268
rect 151136 198228 151142 198240
rect 233970 198228 233976 198240
rect 234028 198228 234034 198280
rect 261478 198228 261484 198280
rect 261536 198268 261542 198280
rect 334158 198268 334164 198280
rect 261536 198240 334164 198268
rect 261536 198228 261542 198240
rect 334158 198228 334164 198240
rect 334216 198228 334222 198280
rect 138934 198160 138940 198212
rect 138992 198200 138998 198212
rect 260926 198200 260932 198212
rect 138992 198172 260932 198200
rect 138992 198160 138998 198172
rect 260926 198160 260932 198172
rect 260984 198160 260990 198212
rect 269758 198160 269764 198212
rect 269816 198200 269822 198212
rect 347774 198200 347780 198212
rect 269816 198172 347780 198200
rect 269816 198160 269822 198172
rect 347774 198160 347780 198172
rect 347832 198160 347838 198212
rect 133230 198092 133236 198144
rect 133288 198132 133294 198144
rect 277486 198132 277492 198144
rect 133288 198104 277492 198132
rect 133288 198092 133294 198104
rect 277486 198092 277492 198104
rect 277544 198092 277550 198144
rect 57790 198024 57796 198076
rect 57848 198064 57854 198076
rect 276106 198064 276112 198076
rect 57848 198036 276112 198064
rect 57848 198024 57854 198036
rect 276106 198024 276112 198036
rect 276164 198024 276170 198076
rect 99374 197956 99380 198008
rect 99432 197996 99438 198008
rect 345290 197996 345296 198008
rect 99432 197968 345296 197996
rect 99432 197956 99438 197968
rect 345290 197956 345296 197968
rect 345348 197956 345354 198008
rect 300118 197276 300124 197328
rect 300176 197316 300182 197328
rect 382182 197316 382188 197328
rect 300176 197288 382188 197316
rect 300176 197276 300182 197288
rect 382182 197276 382188 197288
rect 382240 197316 382246 197328
rect 386874 197316 386880 197328
rect 382240 197288 386880 197316
rect 382240 197276 382246 197288
rect 386874 197276 386880 197288
rect 386932 197276 386938 197328
rect 152642 196868 152648 196920
rect 152700 196908 152706 196920
rect 262398 196908 262404 196920
rect 152700 196880 262404 196908
rect 152700 196868 152706 196880
rect 262398 196868 262404 196880
rect 262456 196868 262462 196920
rect 124858 196800 124864 196852
rect 124916 196840 124922 196852
rect 273346 196840 273352 196852
rect 124916 196812 273352 196840
rect 124916 196800 124922 196812
rect 273346 196800 273352 196812
rect 273404 196800 273410 196852
rect 80054 196732 80060 196784
rect 80112 196772 80118 196784
rect 319530 196772 319536 196784
rect 80112 196744 319536 196772
rect 80112 196732 80118 196744
rect 319530 196732 319536 196744
rect 319588 196732 319594 196784
rect 93946 196664 93952 196716
rect 94004 196704 94010 196716
rect 343726 196704 343732 196716
rect 94004 196676 343732 196704
rect 94004 196664 94010 196676
rect 343726 196664 343732 196676
rect 343784 196664 343790 196716
rect 69106 196596 69112 196648
rect 69164 196636 69170 196648
rect 320818 196636 320824 196648
rect 69164 196608 320824 196636
rect 69164 196596 69170 196608
rect 320818 196596 320824 196608
rect 320876 196596 320882 196648
rect 130654 195440 130660 195492
rect 130712 195480 130718 195492
rect 196710 195480 196716 195492
rect 130712 195452 196716 195480
rect 130712 195440 130718 195452
rect 196710 195440 196716 195452
rect 196768 195440 196774 195492
rect 160094 195372 160100 195424
rect 160152 195412 160158 195424
rect 261018 195412 261024 195424
rect 160152 195384 261024 195412
rect 160152 195372 160158 195384
rect 261018 195372 261024 195384
rect 261076 195372 261082 195424
rect 192478 195304 192484 195356
rect 192536 195344 192542 195356
rect 370590 195344 370596 195356
rect 192536 195316 370596 195344
rect 192536 195304 192542 195316
rect 370590 195304 370596 195316
rect 370648 195304 370654 195356
rect 153838 195236 153844 195288
rect 153896 195276 153902 195288
rect 338850 195276 338856 195288
rect 153896 195248 338856 195276
rect 153896 195236 153902 195248
rect 338850 195236 338856 195248
rect 338908 195236 338914 195288
rect 147122 194080 147128 194132
rect 147180 194120 147186 194132
rect 270586 194120 270592 194132
rect 147180 194092 270592 194120
rect 147180 194080 147186 194092
rect 270586 194080 270592 194092
rect 270644 194080 270650 194132
rect 134610 194012 134616 194064
rect 134668 194052 134674 194064
rect 258166 194052 258172 194064
rect 134668 194024 258172 194052
rect 134668 194012 134674 194024
rect 258166 194012 258172 194024
rect 258224 194012 258230 194064
rect 63402 193944 63408 193996
rect 63460 193984 63466 193996
rect 160738 193984 160744 193996
rect 63460 193956 160744 193984
rect 63460 193944 63466 193956
rect 160738 193944 160744 193956
rect 160796 193944 160802 193996
rect 227714 193944 227720 193996
rect 227772 193984 227778 193996
rect 351914 193984 351920 193996
rect 227772 193956 351920 193984
rect 227772 193944 227778 193956
rect 351914 193944 351920 193956
rect 351972 193944 351978 193996
rect 115934 193876 115940 193928
rect 115992 193916 115998 193928
rect 249058 193916 249064 193928
rect 115992 193888 249064 193916
rect 115992 193876 115998 193888
rect 249058 193876 249064 193888
rect 249116 193876 249122 193928
rect 74626 193808 74632 193860
rect 74684 193848 74690 193860
rect 321646 193848 321652 193860
rect 74684 193820 321652 193848
rect 74684 193808 74690 193820
rect 321646 193808 321652 193820
rect 321704 193808 321710 193860
rect 330478 193808 330484 193860
rect 330536 193848 330542 193860
rect 386414 193848 386420 193860
rect 330536 193820 386420 193848
rect 330536 193808 330542 193820
rect 386414 193808 386420 193820
rect 386472 193808 386478 193860
rect 583846 193128 583852 193180
rect 583904 193128 583910 193180
rect 583864 192976 583892 193128
rect 583846 192924 583852 192976
rect 583904 192924 583910 192976
rect 246298 192856 246304 192908
rect 246356 192896 246362 192908
rect 349338 192896 349344 192908
rect 246356 192868 349344 192896
rect 246356 192856 246362 192868
rect 349338 192856 349344 192868
rect 349396 192856 349402 192908
rect 148318 192788 148324 192840
rect 148376 192828 148382 192840
rect 271966 192828 271972 192840
rect 148376 192800 271972 192828
rect 148376 192788 148382 192800
rect 271966 192788 271972 192800
rect 272024 192788 272030 192840
rect 120810 192720 120816 192772
rect 120868 192760 120874 192772
rect 246390 192760 246396 192772
rect 120868 192732 246396 192760
rect 120868 192720 120874 192732
rect 246390 192720 246396 192732
rect 246448 192720 246454 192772
rect 89714 192652 89720 192704
rect 89772 192692 89778 192704
rect 249978 192692 249984 192704
rect 89772 192664 249984 192692
rect 89772 192652 89778 192664
rect 249978 192652 249984 192664
rect 250036 192652 250042 192704
rect 189718 192584 189724 192636
rect 189776 192624 189782 192636
rect 354030 192624 354036 192636
rect 189776 192596 354036 192624
rect 189776 192584 189782 192596
rect 354030 192584 354036 192596
rect 354088 192584 354094 192636
rect 138750 192516 138756 192568
rect 138808 192556 138814 192568
rect 345198 192556 345204 192568
rect 138808 192528 345204 192556
rect 138808 192516 138814 192528
rect 345198 192516 345204 192528
rect 345256 192516 345262 192568
rect 71774 192448 71780 192500
rect 71832 192488 71838 192500
rect 343818 192488 343824 192500
rect 71832 192460 343824 192488
rect 71832 192448 71838 192460
rect 343818 192448 343824 192460
rect 343876 192448 343882 192500
rect 306282 191836 306288 191888
rect 306340 191876 306346 191888
rect 334066 191876 334072 191888
rect 306340 191848 334072 191876
rect 306340 191836 306374 191848
rect 334066 191836 334072 191848
rect 334124 191836 334130 191888
rect 278130 191768 278136 191820
rect 278188 191808 278194 191820
rect 306346 191808 306374 191836
rect 278188 191780 306374 191808
rect 278188 191768 278194 191780
rect 571702 191700 571708 191752
rect 571760 191740 571766 191752
rect 574186 191740 574192 191752
rect 571760 191712 574192 191740
rect 571760 191700 571766 191712
rect 574186 191700 574192 191712
rect 574244 191700 574250 191752
rect 231854 191360 231860 191412
rect 231912 191400 231918 191412
rect 278038 191400 278044 191412
rect 231912 191372 278044 191400
rect 231912 191360 231918 191372
rect 278038 191360 278044 191372
rect 278096 191360 278102 191412
rect 163498 191292 163504 191344
rect 163556 191332 163562 191344
rect 324406 191332 324412 191344
rect 163556 191304 324412 191332
rect 163556 191292 163562 191304
rect 324406 191292 324412 191304
rect 324464 191292 324470 191344
rect 56502 191224 56508 191276
rect 56560 191264 56566 191276
rect 242250 191264 242256 191276
rect 56560 191236 242256 191264
rect 56560 191224 56566 191236
rect 242250 191224 242256 191236
rect 242308 191224 242314 191276
rect 273898 191224 273904 191276
rect 273956 191264 273962 191276
rect 358078 191264 358084 191276
rect 273956 191236 358084 191264
rect 273956 191224 273962 191236
rect 358078 191224 358084 191236
rect 358136 191224 358142 191276
rect 142982 191156 142988 191208
rect 143040 191196 143046 191208
rect 358814 191196 358820 191208
rect 143040 191168 358820 191196
rect 143040 191156 143046 191168
rect 358814 191156 358820 191168
rect 358872 191156 358878 191208
rect 84286 191088 84292 191140
rect 84344 191128 84350 191140
rect 321554 191128 321560 191140
rect 84344 191100 321560 191128
rect 84344 191088 84350 191100
rect 321554 191088 321560 191100
rect 321612 191088 321618 191140
rect 324958 191088 324964 191140
rect 325016 191128 325022 191140
rect 329098 191128 329104 191140
rect 325016 191100 329104 191128
rect 325016 191088 325022 191100
rect 329098 191088 329104 191100
rect 329156 191088 329162 191140
rect 102042 190476 102048 190528
rect 102100 190516 102106 190528
rect 192478 190516 192484 190528
rect 102100 190488 192484 190516
rect 102100 190476 102106 190488
rect 192478 190476 192484 190488
rect 192536 190476 192542 190528
rect 324406 190408 324412 190460
rect 324464 190448 324470 190460
rect 380250 190448 380256 190460
rect 324464 190420 380256 190448
rect 324464 190408 324470 190420
rect 380250 190408 380256 190420
rect 380308 190408 380314 190460
rect 333238 190340 333244 190392
rect 333296 190380 333302 190392
rect 387058 190380 387064 190392
rect 333296 190352 387064 190380
rect 333296 190340 333302 190352
rect 387058 190340 387064 190352
rect 387116 190340 387122 190392
rect 126422 190000 126428 190052
rect 126480 190040 126486 190052
rect 246482 190040 246488 190052
rect 126480 190012 246488 190040
rect 126480 190000 126486 190012
rect 246482 190000 246488 190012
rect 246540 190000 246546 190052
rect 152550 189932 152556 189984
rect 152608 189972 152614 189984
rect 273438 189972 273444 189984
rect 152608 189944 273444 189972
rect 152608 189932 152614 189944
rect 273438 189932 273444 189944
rect 273496 189932 273502 189984
rect 117958 189864 117964 189916
rect 118016 189904 118022 189916
rect 209038 189904 209044 189916
rect 118016 189876 209044 189904
rect 118016 189864 118022 189876
rect 209038 189864 209044 189876
rect 209096 189864 209102 189916
rect 210418 189864 210424 189916
rect 210476 189904 210482 189916
rect 332042 189904 332048 189916
rect 210476 189876 332048 189904
rect 210476 189864 210482 189876
rect 332042 189864 332048 189876
rect 332100 189864 332106 189916
rect 40678 189796 40684 189848
rect 40736 189836 40742 189848
rect 109678 189836 109684 189848
rect 40736 189808 109684 189836
rect 40736 189796 40742 189808
rect 109678 189796 109684 189808
rect 109736 189796 109742 189848
rect 171778 189796 171784 189848
rect 171836 189836 171842 189848
rect 324498 189836 324504 189848
rect 171836 189808 324504 189836
rect 171836 189796 171842 189808
rect 324498 189796 324504 189808
rect 324556 189796 324562 189848
rect 62022 189728 62028 189780
rect 62080 189768 62086 189780
rect 259638 189768 259644 189780
rect 62080 189740 259644 189768
rect 62080 189728 62086 189740
rect 259638 189728 259644 189740
rect 259696 189728 259702 189780
rect 103422 189048 103428 189100
rect 103480 189088 103486 189100
rect 171962 189088 171968 189100
rect 103480 189060 171968 189088
rect 103480 189048 103486 189060
rect 171962 189048 171968 189060
rect 172020 189048 172026 189100
rect 3418 188980 3424 189032
rect 3476 189020 3482 189032
rect 53098 189020 53104 189032
rect 3476 188992 53104 189020
rect 3476 188980 3482 188992
rect 53098 188980 53104 188992
rect 53156 188980 53162 189032
rect 324498 188980 324504 189032
rect 324556 189020 324562 189032
rect 325050 189020 325056 189032
rect 324556 188992 325056 189020
rect 324556 188980 324562 188992
rect 325050 188980 325056 188992
rect 325108 189020 325114 189032
rect 383010 189020 383016 189032
rect 325108 188992 383016 189020
rect 325108 188980 325114 188992
rect 383010 188980 383016 188992
rect 383068 188980 383074 189032
rect 243538 188572 243544 188624
rect 243596 188612 243602 188624
rect 330478 188612 330484 188624
rect 243596 188584 330484 188612
rect 243596 188572 243602 188584
rect 330478 188572 330484 188584
rect 330536 188572 330542 188624
rect 156598 188504 156604 188556
rect 156656 188544 156662 188556
rect 246298 188544 246304 188556
rect 156656 188516 246304 188544
rect 156656 188504 156662 188516
rect 246298 188504 246304 188516
rect 246356 188504 246362 188556
rect 138842 188436 138848 188488
rect 138900 188476 138906 188488
rect 247770 188476 247776 188488
rect 138900 188448 247776 188476
rect 138900 188436 138906 188448
rect 247770 188436 247776 188448
rect 247828 188436 247834 188488
rect 144270 188368 144276 188420
rect 144328 188408 144334 188420
rect 262214 188408 262220 188420
rect 144328 188380 262220 188408
rect 144328 188368 144334 188380
rect 262214 188368 262220 188380
rect 262272 188368 262278 188420
rect 135990 188300 135996 188352
rect 136048 188340 136054 188352
rect 274726 188340 274732 188352
rect 136048 188312 274732 188340
rect 136048 188300 136054 188312
rect 274726 188300 274732 188312
rect 274784 188300 274790 188352
rect 100662 187688 100668 187740
rect 100720 187728 100726 187740
rect 171778 187728 171784 187740
rect 100720 187700 171784 187728
rect 100720 187688 100726 187700
rect 171778 187688 171784 187700
rect 171836 187688 171842 187740
rect 329190 187620 329196 187672
rect 329248 187660 329254 187672
rect 386782 187660 386788 187672
rect 329248 187632 386788 187660
rect 329248 187620 329254 187632
rect 386782 187620 386788 187632
rect 386840 187620 386846 187672
rect 572622 187620 572628 187672
rect 572680 187660 572686 187672
rect 583478 187660 583484 187672
rect 572680 187632 583484 187660
rect 572680 187620 572686 187632
rect 583478 187620 583484 187632
rect 583536 187620 583542 187672
rect 330478 187552 330484 187604
rect 330536 187592 330542 187604
rect 370498 187592 370504 187604
rect 330536 187564 370504 187592
rect 330536 187552 330542 187564
rect 370498 187552 370504 187564
rect 370556 187552 370562 187604
rect 161382 187144 161388 187196
rect 161440 187184 161446 187196
rect 195238 187184 195244 187196
rect 161440 187156 195244 187184
rect 161440 187144 161446 187156
rect 195238 187144 195244 187156
rect 195296 187144 195302 187196
rect 104894 187076 104900 187128
rect 104952 187116 104958 187128
rect 188338 187116 188344 187128
rect 104952 187088 188344 187116
rect 104952 187076 104958 187088
rect 188338 187076 188344 187088
rect 188396 187076 188402 187128
rect 162302 187008 162308 187060
rect 162360 187048 162366 187060
rect 327258 187048 327264 187060
rect 162360 187020 327264 187048
rect 162360 187008 162366 187020
rect 327258 187008 327264 187020
rect 327316 187008 327322 187060
rect 95234 186940 95240 186992
rect 95292 186980 95298 186992
rect 320174 186980 320180 186992
rect 95292 186952 320180 186980
rect 95292 186940 95298 186952
rect 320174 186940 320180 186952
rect 320232 186940 320238 186992
rect 126882 186328 126888 186380
rect 126940 186368 126946 186380
rect 169110 186368 169116 186380
rect 126940 186340 169116 186368
rect 126940 186328 126946 186340
rect 169110 186328 169116 186340
rect 169168 186328 169174 186380
rect 131942 185852 131948 185904
rect 132000 185892 132006 185904
rect 243538 185892 243544 185904
rect 132000 185864 243544 185892
rect 132000 185852 132006 185864
rect 243538 185852 243544 185864
rect 243596 185852 243602 185904
rect 170398 185784 170404 185836
rect 170456 185824 170462 185836
rect 324958 185824 324964 185836
rect 170456 185796 324964 185824
rect 170456 185784 170462 185796
rect 324958 185784 324964 185796
rect 325016 185784 325022 185836
rect 60642 185716 60648 185768
rect 60700 185756 60706 185768
rect 254026 185756 254032 185768
rect 60700 185728 254032 185756
rect 60700 185716 60706 185728
rect 254026 185716 254032 185728
rect 254084 185716 254090 185768
rect 102134 185648 102140 185700
rect 102192 185688 102198 185700
rect 323118 185688 323124 185700
rect 102192 185660 323124 185688
rect 102192 185648 102198 185660
rect 323118 185648 323124 185660
rect 323176 185648 323182 185700
rect 66070 185580 66076 185632
rect 66128 185620 66134 185632
rect 324498 185620 324504 185632
rect 66128 185592 324504 185620
rect 66128 185580 66134 185592
rect 324498 185580 324504 185592
rect 324556 185580 324562 185632
rect 329190 185580 329196 185632
rect 329248 185620 329254 185632
rect 386874 185620 386880 185632
rect 329248 185592 386880 185620
rect 329248 185580 329254 185592
rect 386874 185580 386880 185592
rect 386932 185580 386938 185632
rect 115842 184968 115848 185020
rect 115900 185008 115906 185020
rect 170490 185008 170496 185020
rect 115900 184980 170496 185008
rect 115900 184968 115906 184980
rect 170490 184968 170496 184980
rect 170548 184968 170554 185020
rect 122742 184900 122748 184952
rect 122800 184940 122806 184952
rect 211982 184940 211988 184952
rect 122800 184912 211988 184940
rect 122800 184900 122806 184912
rect 211982 184900 211988 184912
rect 212040 184900 212046 184952
rect 571426 184832 571432 184884
rect 571484 184872 571490 184884
rect 574094 184872 574100 184884
rect 571484 184844 574100 184872
rect 571484 184832 571490 184844
rect 574094 184832 574100 184844
rect 574152 184832 574158 184884
rect 160002 184424 160008 184476
rect 160060 184464 160066 184476
rect 189718 184464 189724 184476
rect 160060 184436 189724 184464
rect 160060 184424 160066 184436
rect 189718 184424 189724 184436
rect 189776 184424 189782 184476
rect 126238 184356 126244 184408
rect 126296 184396 126302 184408
rect 266538 184396 266544 184408
rect 126296 184368 266544 184396
rect 126296 184356 126302 184368
rect 266538 184356 266544 184368
rect 266596 184356 266602 184408
rect 148410 184288 148416 184340
rect 148468 184328 148474 184340
rect 337470 184328 337476 184340
rect 148468 184300 337476 184328
rect 148468 184288 148474 184300
rect 337470 184288 337476 184300
rect 337528 184288 337534 184340
rect 84194 184220 84200 184272
rect 84252 184260 84258 184272
rect 321830 184260 321836 184272
rect 84252 184232 321836 184260
rect 84252 184220 84258 184232
rect 321830 184220 321836 184232
rect 321888 184220 321894 184272
rect 77294 184152 77300 184204
rect 77352 184192 77358 184204
rect 318058 184192 318064 184204
rect 77352 184164 318064 184192
rect 77352 184152 77358 184164
rect 318058 184152 318064 184164
rect 318116 184152 318122 184204
rect 119982 183540 119988 183592
rect 120040 183580 120046 183592
rect 170674 183580 170680 183592
rect 120040 183552 170680 183580
rect 120040 183540 120046 183552
rect 170674 183540 170680 183552
rect 170732 183540 170738 183592
rect 237374 182996 237380 183048
rect 237432 183036 237438 183048
rect 271138 183036 271144 183048
rect 237432 183008 271144 183036
rect 237432 182996 237438 183008
rect 271138 182996 271144 183008
rect 271196 182996 271202 183048
rect 93854 182928 93860 182980
rect 93912 182968 93918 182980
rect 253934 182968 253940 182980
rect 93912 182940 253940 182968
rect 93912 182928 93918 182940
rect 253934 182928 253940 182940
rect 253992 182928 253998 182980
rect 283650 182928 283656 182980
rect 283708 182968 283714 182980
rect 342530 182968 342536 182980
rect 283708 182940 342536 182968
rect 283708 182928 283714 182940
rect 342530 182928 342536 182940
rect 342588 182928 342594 182980
rect 167638 182860 167644 182912
rect 167696 182900 167702 182912
rect 339494 182900 339500 182912
rect 167696 182872 339500 182900
rect 167696 182860 167702 182872
rect 339494 182860 339500 182872
rect 339552 182860 339558 182912
rect 106918 182792 106924 182844
rect 106976 182832 106982 182844
rect 350626 182832 350632 182844
rect 106976 182804 350632 182832
rect 106976 182792 106982 182804
rect 350626 182792 350632 182804
rect 350684 182792 350690 182844
rect 130746 182248 130752 182300
rect 130804 182288 130810 182300
rect 206370 182288 206376 182300
rect 130804 182260 206376 182288
rect 130804 182248 130810 182260
rect 206370 182248 206376 182260
rect 206428 182248 206434 182300
rect 110690 182180 110696 182232
rect 110748 182220 110754 182232
rect 214558 182220 214564 182232
rect 110748 182192 214564 182220
rect 110748 182180 110754 182192
rect 214558 182180 214564 182192
rect 214616 182180 214622 182232
rect 341518 182180 341524 182232
rect 341576 182220 341582 182232
rect 386414 182220 386420 182232
rect 341576 182192 386420 182220
rect 341576 182180 341582 182192
rect 386414 182180 386420 182192
rect 386472 182180 386478 182232
rect 222838 181636 222844 181688
rect 222896 181676 222902 181688
rect 266446 181676 266452 181688
rect 222896 181648 266452 181676
rect 222896 181636 222902 181648
rect 266446 181636 266452 181648
rect 266504 181636 266510 181688
rect 311158 181636 311164 181688
rect 311216 181676 311222 181688
rect 341058 181676 341064 181688
rect 311216 181648 341064 181676
rect 311216 181636 311222 181648
rect 341058 181636 341064 181648
rect 341116 181636 341122 181688
rect 211062 181568 211068 181620
rect 211120 181608 211126 181620
rect 220814 181608 220820 181620
rect 211120 181580 220820 181608
rect 211120 181568 211126 181580
rect 220814 181568 220820 181580
rect 220872 181568 220878 181620
rect 225598 181568 225604 181620
rect 225656 181608 225662 181620
rect 335630 181608 335636 181620
rect 225656 181580 335636 181608
rect 225656 181568 225662 181580
rect 335630 181568 335636 181580
rect 335688 181568 335694 181620
rect 171870 181500 171876 181552
rect 171928 181540 171934 181552
rect 251266 181540 251272 181552
rect 171928 181512 251272 181540
rect 171928 181500 171934 181512
rect 251266 181500 251272 181512
rect 251324 181500 251330 181552
rect 271230 181500 271236 181552
rect 271288 181540 271294 181552
rect 381630 181540 381636 181552
rect 271288 181512 381636 181540
rect 271288 181500 271294 181512
rect 381630 181500 381636 181512
rect 381688 181500 381694 181552
rect 154482 181432 154488 181484
rect 154540 181472 154546 181484
rect 197998 181472 198004 181484
rect 154540 181444 198004 181472
rect 154540 181432 154546 181444
rect 197998 181432 198004 181444
rect 198056 181432 198062 181484
rect 203610 181432 203616 181484
rect 203668 181472 203674 181484
rect 356882 181472 356888 181484
rect 203668 181444 356888 181472
rect 203668 181432 203674 181444
rect 356882 181432 356888 181444
rect 356940 181432 356946 181484
rect 121086 180956 121092 181008
rect 121144 180996 121150 181008
rect 166534 180996 166540 181008
rect 121144 180968 166540 180996
rect 121144 180956 121150 180968
rect 166534 180956 166540 180968
rect 166592 180956 166598 181008
rect 112990 180888 112996 180940
rect 113048 180928 113054 180940
rect 167730 180928 167736 180940
rect 113048 180900 167736 180928
rect 113048 180888 113054 180900
rect 167730 180888 167736 180900
rect 167788 180888 167794 180940
rect 128078 180820 128084 180872
rect 128136 180860 128142 180872
rect 214650 180860 214656 180872
rect 128136 180832 214656 180860
rect 128136 180820 128142 180832
rect 214650 180820 214656 180832
rect 214708 180820 214714 180872
rect 242158 180412 242164 180464
rect 242216 180452 242222 180464
rect 256786 180452 256792 180464
rect 242216 180424 256792 180452
rect 242216 180412 242222 180424
rect 256786 180412 256792 180424
rect 256844 180412 256850 180464
rect 240778 180344 240784 180396
rect 240836 180384 240842 180396
rect 258350 180384 258356 180396
rect 240836 180356 258356 180384
rect 240836 180344 240842 180356
rect 258350 180344 258356 180356
rect 258408 180344 258414 180396
rect 166902 180276 166908 180328
rect 166960 180316 166966 180328
rect 182818 180316 182824 180328
rect 166960 180288 182824 180316
rect 166960 180276 166966 180288
rect 182818 180276 182824 180288
rect 182876 180276 182882 180328
rect 238110 180276 238116 180328
rect 238168 180316 238174 180328
rect 263686 180316 263692 180328
rect 238168 180288 263692 180316
rect 238168 180276 238174 180288
rect 263686 180276 263692 180288
rect 263744 180276 263750 180328
rect 315390 180276 315396 180328
rect 315448 180316 315454 180328
rect 346486 180316 346492 180328
rect 315448 180288 346492 180316
rect 315448 180276 315454 180288
rect 346486 180276 346492 180288
rect 346544 180276 346550 180328
rect 158622 180208 158628 180260
rect 158680 180248 158686 180260
rect 184198 180248 184204 180260
rect 158680 180220 184204 180248
rect 158680 180208 158686 180220
rect 184198 180208 184204 180220
rect 184256 180208 184262 180260
rect 209038 180208 209044 180260
rect 209096 180248 209102 180260
rect 272058 180248 272064 180260
rect 209096 180220 272064 180248
rect 209096 180208 209102 180220
rect 272058 180208 272064 180220
rect 272116 180208 272122 180260
rect 300210 180208 300216 180260
rect 300268 180248 300274 180260
rect 345106 180248 345112 180260
rect 300268 180220 345112 180248
rect 300268 180208 300274 180220
rect 345106 180208 345112 180220
rect 345164 180208 345170 180260
rect 66162 180140 66168 180192
rect 66220 180180 66226 180192
rect 251358 180180 251364 180192
rect 66220 180152 251364 180180
rect 66220 180140 66226 180152
rect 251358 180140 251364 180152
rect 251416 180140 251422 180192
rect 280062 180140 280068 180192
rect 280120 180180 280126 180192
rect 380434 180180 380440 180192
rect 280120 180152 380440 180180
rect 280120 180140 280126 180152
rect 380434 180140 380440 180152
rect 380492 180140 380498 180192
rect 68922 180072 68928 180124
rect 68980 180112 68986 180124
rect 321738 180112 321744 180124
rect 68980 180084 321744 180112
rect 68980 180072 68986 180084
rect 321738 180072 321744 180084
rect 321796 180072 321802 180124
rect 132034 179528 132040 179580
rect 132092 179568 132098 179580
rect 165338 179568 165344 179580
rect 132092 179540 165344 179568
rect 132092 179528 132098 179540
rect 165338 179528 165344 179540
rect 165396 179528 165402 179580
rect 110230 179460 110236 179512
rect 110288 179500 110294 179512
rect 167822 179500 167828 179512
rect 110288 179472 167828 179500
rect 110288 179460 110294 179472
rect 167822 179460 167828 179472
rect 167880 179460 167886 179512
rect 114370 179392 114376 179444
rect 114428 179432 114434 179444
rect 210418 179432 210424 179444
rect 114428 179404 210424 179432
rect 114428 179392 114434 179404
rect 210418 179392 210424 179404
rect 210476 179392 210482 179444
rect 246482 178984 246488 179036
rect 246540 179024 246546 179036
rect 252554 179024 252560 179036
rect 246540 178996 252560 179024
rect 246540 178984 246546 178996
rect 252554 178984 252560 178996
rect 252612 178984 252618 179036
rect 247770 178916 247776 178968
rect 247828 178956 247834 178968
rect 249334 178956 249340 178968
rect 247828 178928 249340 178956
rect 247828 178916 247834 178928
rect 249334 178916 249340 178928
rect 249392 178916 249398 178968
rect 233970 178848 233976 178900
rect 234028 178888 234034 178900
rect 249426 178888 249432 178900
rect 234028 178860 249432 178888
rect 234028 178848 234034 178860
rect 249426 178848 249432 178860
rect 249484 178848 249490 178900
rect 220078 178780 220084 178832
rect 220136 178820 220142 178832
rect 265158 178820 265164 178832
rect 220136 178792 265164 178820
rect 220136 178780 220142 178792
rect 265158 178780 265164 178792
rect 265216 178780 265222 178832
rect 317322 178780 317328 178832
rect 317380 178820 317386 178832
rect 337378 178820 337384 178832
rect 317380 178792 337384 178820
rect 317380 178780 317386 178792
rect 337378 178780 337384 178792
rect 337436 178780 337442 178832
rect 211890 178712 211896 178764
rect 211948 178752 211954 178764
rect 258074 178752 258080 178764
rect 211948 178724 258080 178752
rect 211948 178712 211954 178724
rect 258074 178712 258080 178724
rect 258132 178712 258138 178764
rect 289078 178712 289084 178764
rect 289136 178752 289142 178764
rect 325786 178752 325792 178764
rect 289136 178724 325792 178752
rect 289136 178712 289142 178724
rect 325786 178712 325792 178724
rect 325844 178712 325850 178764
rect 146938 178644 146944 178696
rect 146996 178684 147002 178696
rect 254118 178684 254124 178696
rect 146996 178656 254124 178684
rect 146996 178644 147002 178656
rect 254118 178644 254124 178656
rect 254176 178644 254182 178696
rect 305638 178644 305644 178696
rect 305696 178684 305702 178696
rect 363690 178684 363696 178696
rect 305696 178656 363696 178684
rect 305696 178644 305702 178656
rect 363690 178644 363696 178656
rect 363748 178644 363754 178696
rect 318058 178508 318064 178560
rect 318116 178548 318122 178560
rect 323026 178548 323032 178560
rect 318116 178520 323032 178548
rect 318116 178508 318122 178520
rect 323026 178508 323032 178520
rect 323084 178508 323090 178560
rect 148226 178236 148232 178288
rect 148284 178276 148290 178288
rect 166442 178276 166448 178288
rect 148284 178248 166448 178276
rect 148284 178236 148290 178248
rect 166442 178236 166448 178248
rect 166500 178236 166506 178288
rect 123018 178168 123024 178220
rect 123076 178208 123082 178220
rect 169294 178208 169300 178220
rect 123076 178180 169300 178208
rect 123076 178168 123082 178180
rect 169294 178168 169300 178180
rect 169352 178168 169358 178220
rect 118418 178100 118424 178152
rect 118476 178140 118482 178152
rect 166626 178140 166632 178152
rect 118476 178112 166632 178140
rect 118476 178100 118482 178112
rect 166626 178100 166632 178112
rect 166684 178100 166690 178152
rect 129458 178032 129464 178084
rect 129516 178072 129522 178084
rect 214190 178072 214196 178084
rect 129516 178044 214196 178072
rect 129516 178032 129522 178044
rect 214190 178032 214196 178044
rect 214248 178032 214254 178084
rect 326430 177964 326436 178016
rect 326488 178004 326494 178016
rect 386874 178004 386880 178016
rect 326488 177976 386880 178004
rect 326488 177964 326494 177976
rect 386874 177964 386880 177976
rect 386932 177964 386938 178016
rect 572070 177964 572076 178016
rect 572128 178004 572134 178016
rect 576302 178004 576308 178016
rect 572128 177976 576308 178004
rect 572128 177964 572134 177976
rect 576302 177964 576308 177976
rect 576360 177964 576366 178016
rect 258166 177760 258172 177812
rect 258224 177800 258230 177812
rect 258224 177772 267734 177800
rect 258224 177760 258230 177772
rect 242250 177556 242256 177608
rect 242308 177596 242314 177608
rect 258258 177596 258264 177608
rect 242308 177568 258264 177596
rect 242308 177556 242314 177568
rect 258258 177556 258264 177568
rect 258316 177556 258322 177608
rect 171042 177488 171048 177540
rect 171100 177528 171106 177540
rect 215938 177528 215944 177540
rect 171100 177500 215944 177528
rect 171100 177488 171106 177500
rect 215938 177488 215944 177500
rect 215996 177488 216002 177540
rect 239398 177488 239404 177540
rect 239456 177528 239462 177540
rect 256970 177528 256976 177540
rect 239456 177500 256976 177528
rect 239456 177488 239462 177500
rect 256970 177488 256976 177500
rect 257028 177488 257034 177540
rect 196710 177420 196716 177472
rect 196768 177460 196774 177472
rect 249242 177460 249248 177472
rect 196768 177432 249248 177460
rect 196768 177420 196774 177432
rect 249242 177420 249248 177432
rect 249300 177420 249306 177472
rect 267706 177460 267734 177772
rect 314010 177556 314016 177608
rect 314068 177596 314074 177608
rect 332778 177596 332784 177608
rect 314068 177568 332784 177596
rect 314068 177556 314074 177568
rect 332778 177556 332784 177568
rect 332836 177556 332842 177608
rect 311250 177488 311256 177540
rect 311308 177528 311314 177540
rect 338758 177528 338764 177540
rect 311308 177500 338764 177528
rect 311308 177488 311314 177500
rect 338758 177488 338764 177500
rect 338816 177488 338822 177540
rect 269114 177460 269120 177472
rect 267706 177432 269120 177460
rect 269114 177420 269120 177432
rect 269172 177420 269178 177472
rect 275278 177420 275284 177472
rect 275336 177460 275342 177472
rect 328546 177460 328552 177472
rect 275336 177432 328552 177460
rect 275336 177420 275342 177432
rect 328546 177420 328552 177432
rect 328604 177420 328610 177472
rect 164878 177352 164884 177404
rect 164936 177392 164942 177404
rect 251450 177392 251456 177404
rect 164936 177364 251456 177392
rect 164936 177352 164942 177364
rect 251450 177352 251456 177364
rect 251508 177352 251514 177404
rect 264238 177352 264244 177404
rect 264296 177392 264302 177404
rect 365070 177392 365076 177404
rect 264296 177364 365076 177392
rect 264296 177352 264302 177364
rect 365070 177352 365076 177364
rect 365128 177352 365134 177404
rect 166350 177284 166356 177336
rect 166408 177324 166414 177336
rect 325878 177324 325884 177336
rect 166408 177296 325884 177324
rect 166408 177284 166414 177296
rect 325878 177284 325884 177296
rect 325936 177284 325942 177336
rect 104618 177012 104624 177064
rect 104676 177052 104682 177064
rect 170582 177052 170588 177064
rect 104676 177024 170588 177052
rect 104676 177012 104682 177024
rect 170582 177012 170588 177024
rect 170640 177012 170646 177064
rect 133138 176944 133144 176996
rect 133196 176984 133202 176996
rect 164510 176984 164516 176996
rect 133196 176956 164516 176984
rect 133196 176944 133202 176956
rect 164510 176944 164516 176956
rect 164568 176944 164574 176996
rect 128170 176876 128176 176928
rect 128228 176916 128234 176928
rect 165430 176916 165436 176928
rect 128228 176888 165436 176916
rect 128228 176876 128234 176888
rect 165430 176876 165436 176888
rect 165488 176876 165494 176928
rect 108114 176808 108120 176860
rect 108172 176848 108178 176860
rect 169018 176848 169024 176860
rect 108172 176820 169024 176848
rect 108172 176808 108178 176820
rect 169018 176808 169024 176820
rect 169076 176808 169082 176860
rect 107010 176740 107016 176792
rect 107068 176780 107074 176792
rect 171870 176780 171876 176792
rect 107068 176752 171876 176780
rect 107068 176740 107074 176752
rect 171870 176740 171876 176752
rect 171928 176740 171934 176792
rect 158990 176672 158996 176724
rect 159048 176712 159054 176724
rect 166258 176712 166264 176724
rect 159048 176684 166264 176712
rect 159048 176672 159054 176684
rect 166258 176672 166264 176684
rect 166316 176672 166322 176724
rect 135714 176604 135720 176656
rect 135772 176644 135778 176656
rect 213914 176644 213920 176656
rect 135772 176616 213920 176644
rect 135772 176604 135778 176616
rect 213914 176604 213920 176616
rect 213972 176604 213978 176656
rect 235258 176604 235264 176656
rect 235316 176644 235322 176656
rect 248046 176644 248052 176656
rect 235316 176616 248052 176644
rect 235316 176604 235322 176616
rect 248046 176604 248052 176616
rect 248104 176604 248110 176656
rect 324314 176604 324320 176656
rect 324372 176644 324378 176656
rect 380342 176644 380348 176656
rect 324372 176616 380348 176644
rect 324372 176604 324378 176616
rect 380342 176604 380348 176616
rect 380400 176604 380406 176656
rect 246298 176536 246304 176588
rect 246356 176576 246362 176588
rect 255314 176576 255320 176588
rect 246356 176548 255320 176576
rect 246356 176536 246362 176548
rect 255314 176536 255320 176548
rect 255372 176536 255378 176588
rect 134426 176196 134432 176248
rect 134484 176236 134490 176248
rect 165522 176236 165528 176248
rect 134484 176208 165528 176236
rect 134484 176196 134490 176208
rect 165522 176196 165528 176208
rect 165580 176196 165586 176248
rect 124490 176128 124496 176180
rect 124548 176168 124554 176180
rect 167914 176168 167920 176180
rect 124548 176140 167920 176168
rect 124548 176128 124554 176140
rect 167914 176128 167920 176140
rect 167972 176128 167978 176180
rect 319530 176128 319536 176180
rect 319588 176168 319594 176180
rect 334250 176168 334256 176180
rect 319588 176140 334256 176168
rect 319588 176128 319594 176140
rect 334250 176128 334256 176140
rect 334308 176128 334314 176180
rect 116946 176060 116952 176112
rect 117004 176100 117010 176112
rect 169202 176100 169208 176112
rect 117004 176072 169208 176100
rect 117004 176060 117010 176072
rect 169202 176060 169208 176072
rect 169260 176060 169266 176112
rect 312538 176060 312544 176112
rect 312596 176100 312602 176112
rect 327350 176100 327356 176112
rect 312596 176072 327356 176100
rect 312596 176060 312602 176072
rect 327350 176060 327356 176072
rect 327408 176060 327414 176112
rect 98362 175992 98368 176044
rect 98420 176032 98426 176044
rect 170398 176032 170404 176044
rect 98420 176004 170404 176032
rect 98420 175992 98426 176004
rect 170398 175992 170404 176004
rect 170456 175992 170462 176044
rect 307018 175992 307024 176044
rect 307076 176032 307082 176044
rect 343634 176032 343640 176044
rect 307076 176004 343640 176032
rect 307076 175992 307082 176004
rect 343634 175992 343640 176004
rect 343692 175992 343698 176044
rect 4798 175924 4804 175976
rect 4856 175964 4862 175976
rect 110414 175964 110420 175976
rect 4856 175936 110420 175964
rect 4856 175924 4862 175936
rect 110414 175924 110420 175936
rect 110472 175924 110478 175976
rect 160738 175924 160744 175976
rect 160796 175964 160802 175976
rect 259730 175964 259736 175976
rect 160796 175936 259736 175964
rect 160796 175924 160802 175936
rect 259730 175924 259736 175936
rect 259788 175924 259794 175976
rect 283558 175924 283564 175976
rect 283616 175964 283622 175976
rect 329926 175964 329932 175976
rect 283616 175936 329932 175964
rect 283616 175924 283622 175936
rect 329926 175924 329932 175936
rect 329984 175924 329990 175976
rect 243538 175788 243544 175840
rect 243596 175828 243602 175840
rect 249150 175828 249156 175840
rect 243596 175800 249156 175828
rect 243596 175788 243602 175800
rect 249150 175788 249156 175800
rect 249208 175788 249214 175840
rect 164510 175176 164516 175228
rect 164568 175216 164574 175228
rect 214006 175216 214012 175228
rect 164568 175188 214012 175216
rect 164568 175176 164574 175188
rect 214006 175176 214012 175188
rect 214064 175176 214070 175228
rect 324314 175176 324320 175228
rect 324372 175216 324378 175228
rect 360286 175216 360292 175228
rect 324372 175188 360292 175216
rect 324372 175176 324378 175188
rect 360286 175176 360292 175188
rect 360344 175176 360350 175228
rect 165522 175108 165528 175160
rect 165580 175148 165586 175160
rect 213914 175148 213920 175160
rect 165580 175120 213920 175148
rect 165580 175108 165586 175120
rect 213914 175108 213920 175120
rect 213972 175108 213978 175160
rect 3694 163480 3700 163532
rect 3752 163520 3758 163532
rect 4062 163520 4068 163532
rect 3752 163492 4068 163520
rect 3752 163480 3758 163492
rect 4062 163480 4068 163492
rect 4120 163520 4126 163532
rect 66898 163520 66904 163532
rect 4120 163492 66904 163520
rect 4120 163480 4126 163492
rect 66898 163480 66904 163492
rect 66956 163480 66962 163532
rect 3418 150356 3424 150408
rect 3476 150396 3482 150408
rect 31018 150396 31024 150408
rect 3476 150368 31024 150396
rect 3476 150356 3482 150368
rect 31018 150356 31024 150368
rect 31076 150356 31082 150408
rect 3234 137912 3240 137964
rect 3292 137952 3298 137964
rect 17218 137952 17224 137964
rect 3292 137924 17224 137952
rect 3292 137912 3298 137924
rect 17218 137912 17224 137924
rect 17276 137912 17282 137964
rect 60642 128324 60648 128376
rect 60700 128364 60706 128376
rect 66070 128364 66076 128376
rect 60700 128336 66076 128364
rect 60700 128324 60706 128336
rect 66070 128324 66076 128336
rect 66128 128324 66134 128376
rect 57882 125604 57888 125656
rect 57940 125644 57946 125656
rect 66162 125644 66168 125656
rect 57940 125616 66168 125644
rect 57940 125604 57946 125616
rect 66162 125604 66168 125616
rect 66220 125604 66226 125656
rect 63310 122816 63316 122868
rect 63368 122856 63374 122868
rect 66070 122856 66076 122868
rect 63368 122828 66076 122856
rect 63368 122816 63374 122828
rect 66070 122816 66076 122828
rect 66128 122816 66134 122868
rect 63402 121456 63408 121508
rect 63460 121496 63466 121508
rect 66162 121496 66168 121508
rect 63460 121468 66168 121496
rect 63460 121456 63466 121468
rect 66162 121456 66168 121468
rect 66220 121456 66226 121508
rect 2774 110712 2780 110764
rect 2832 110752 2838 110764
rect 4798 110752 4804 110764
rect 2832 110724 4804 110752
rect 2832 110712 2838 110724
rect 4798 110712 4804 110724
rect 4856 110712 4862 110764
rect 3418 97588 3424 97640
rect 3476 97628 3482 97640
rect 7558 97628 7564 97640
rect 3476 97600 7564 97628
rect 3476 97588 3482 97600
rect 7558 97588 7564 97600
rect 7616 97588 7622 97640
rect 165430 174496 165436 174548
rect 165488 174536 165494 174548
rect 214098 174536 214104 174548
rect 165488 174508 214104 174536
rect 165488 174496 165494 174508
rect 214098 174496 214104 174508
rect 214156 174496 214162 174548
rect 283742 174020 283748 174072
rect 283800 174060 283806 174072
rect 307294 174060 307300 174072
rect 283800 174032 307300 174060
rect 283800 174020 283806 174032
rect 307294 174020 307300 174032
rect 307352 174020 307358 174072
rect 274082 173952 274088 174004
rect 274140 173992 274146 174004
rect 306742 173992 306748 174004
rect 274140 173964 306748 173992
rect 274140 173952 274146 173964
rect 306742 173952 306748 173964
rect 306800 173952 306806 174004
rect 264238 173884 264244 173936
rect 264296 173924 264302 173936
rect 307662 173924 307668 173936
rect 264296 173896 307668 173924
rect 264296 173884 264302 173896
rect 307662 173884 307668 173896
rect 307720 173884 307726 173936
rect 165338 173816 165344 173868
rect 165396 173856 165402 173868
rect 213914 173856 213920 173868
rect 165396 173828 213920 173856
rect 165396 173816 165402 173828
rect 213914 173816 213920 173828
rect 213972 173816 213978 173868
rect 354030 173816 354036 173868
rect 354088 173856 354094 173868
rect 387150 173856 387156 173868
rect 354088 173828 387156 173856
rect 354088 173816 354094 173828
rect 387150 173816 387156 173828
rect 387208 173856 387214 173868
rect 387610 173856 387616 173868
rect 387208 173828 387616 173856
rect 387208 173816 387214 173828
rect 387610 173816 387616 173828
rect 387668 173816 387674 173868
rect 206370 173748 206376 173800
rect 206428 173788 206434 173800
rect 214006 173788 214012 173800
rect 206428 173760 214012 173788
rect 206428 173748 206434 173760
rect 214006 173748 214012 173760
rect 214064 173748 214070 173800
rect 283650 172660 283656 172712
rect 283708 172700 283714 172712
rect 307570 172700 307576 172712
rect 283708 172672 307576 172700
rect 283708 172660 283714 172672
rect 307570 172660 307576 172672
rect 307628 172660 307634 172712
rect 269758 172592 269764 172644
rect 269816 172632 269822 172644
rect 307294 172632 307300 172644
rect 269816 172604 307300 172632
rect 269816 172592 269822 172604
rect 307294 172592 307300 172604
rect 307352 172592 307358 172644
rect 261662 172524 261668 172576
rect 261720 172564 261726 172576
rect 307662 172564 307668 172576
rect 261720 172536 307668 172564
rect 261720 172524 261726 172536
rect 307662 172524 307668 172536
rect 307720 172524 307726 172576
rect 324314 172456 324320 172508
rect 324372 172496 324378 172508
rect 385126 172496 385132 172508
rect 324372 172468 385132 172496
rect 324372 172456 324378 172468
rect 385126 172456 385132 172468
rect 385184 172456 385190 172508
rect 251818 171844 251824 171896
rect 251876 171884 251882 171896
rect 258074 171884 258080 171896
rect 251876 171856 258080 171884
rect 251876 171844 251882 171856
rect 258074 171844 258080 171856
rect 258132 171844 258138 171896
rect 166994 171776 167000 171828
rect 167052 171816 167058 171828
rect 214650 171816 214656 171828
rect 167052 171788 214656 171816
rect 167052 171776 167058 171788
rect 214650 171776 214656 171788
rect 214708 171776 214714 171828
rect 289446 171232 289452 171284
rect 289504 171272 289510 171284
rect 306926 171272 306932 171284
rect 289504 171244 306932 171272
rect 289504 171232 289510 171244
rect 306926 171232 306932 171244
rect 306984 171232 306990 171284
rect 268470 171164 268476 171216
rect 268528 171204 268534 171216
rect 307662 171204 307668 171216
rect 268528 171176 307668 171204
rect 268528 171164 268534 171176
rect 307662 171164 307668 171176
rect 307720 171164 307726 171216
rect 262858 171096 262864 171148
rect 262916 171136 262922 171148
rect 306558 171136 306564 171148
rect 262916 171108 306564 171136
rect 262916 171096 262922 171108
rect 306558 171096 306564 171108
rect 306616 171096 306622 171148
rect 324866 171096 324872 171148
rect 324924 171136 324930 171148
rect 354030 171136 354036 171148
rect 324924 171108 354036 171136
rect 324924 171096 324930 171108
rect 354030 171096 354036 171108
rect 354088 171096 354094 171148
rect 169110 171028 169116 171080
rect 169168 171068 169174 171080
rect 213914 171068 213920 171080
rect 169168 171040 213920 171068
rect 169168 171028 169174 171040
rect 213914 171028 213920 171040
rect 213972 171028 213978 171080
rect 251726 171028 251732 171080
rect 251784 171068 251790 171080
rect 256694 171068 256700 171080
rect 251784 171040 256700 171068
rect 251784 171028 251790 171040
rect 256694 171028 256700 171040
rect 256752 171028 256758 171080
rect 324314 171028 324320 171080
rect 324372 171068 324378 171080
rect 382274 171068 382280 171080
rect 324372 171040 382280 171068
rect 324372 171028 324378 171040
rect 382274 171028 382280 171040
rect 382332 171028 382338 171080
rect 356882 170280 356888 170332
rect 356940 170320 356946 170332
rect 359642 170320 359648 170332
rect 356940 170292 359648 170320
rect 356940 170280 356946 170292
rect 359642 170280 359648 170292
rect 359700 170280 359706 170332
rect 282270 169872 282276 169924
rect 282328 169912 282334 169924
rect 307662 169912 307668 169924
rect 282328 169884 307668 169912
rect 282328 169872 282334 169884
rect 307662 169872 307668 169884
rect 307720 169872 307726 169924
rect 251818 169804 251824 169856
rect 251876 169844 251882 169856
rect 259638 169844 259644 169856
rect 251876 169816 259644 169844
rect 251876 169804 251882 169816
rect 259638 169804 259644 169816
rect 259696 169804 259702 169856
rect 265618 169804 265624 169856
rect 265676 169844 265682 169856
rect 307294 169844 307300 169856
rect 265676 169816 307300 169844
rect 265676 169804 265682 169816
rect 307294 169804 307300 169816
rect 307352 169804 307358 169856
rect 257338 169736 257344 169788
rect 257396 169776 257402 169788
rect 306742 169776 306748 169788
rect 257396 169748 306748 169776
rect 257396 169736 257402 169748
rect 306742 169736 306748 169748
rect 306800 169736 306806 169788
rect 324314 169736 324320 169788
rect 324372 169776 324378 169788
rect 356790 169776 356796 169788
rect 324372 169748 356796 169776
rect 324372 169736 324378 169748
rect 356790 169736 356796 169748
rect 356848 169736 356854 169788
rect 572622 169736 572628 169788
rect 572680 169776 572686 169788
rect 576854 169776 576860 169788
rect 572680 169748 576860 169776
rect 572680 169736 572686 169748
rect 576854 169736 576860 169748
rect 576912 169736 576918 169788
rect 167914 169668 167920 169720
rect 167972 169708 167978 169720
rect 213914 169708 213920 169720
rect 167972 169680 213920 169708
rect 167972 169668 167978 169680
rect 213914 169668 213920 169680
rect 213972 169668 213978 169720
rect 324498 169668 324504 169720
rect 324556 169708 324562 169720
rect 329190 169708 329196 169720
rect 324556 169680 329196 169708
rect 324556 169668 324562 169680
rect 329190 169668 329196 169680
rect 329248 169668 329254 169720
rect 332042 169668 332048 169720
rect 332100 169708 332106 169720
rect 386874 169708 386880 169720
rect 332100 169680 386880 169708
rect 332100 169668 332106 169680
rect 386874 169668 386880 169680
rect 386932 169668 386938 169720
rect 169294 169600 169300 169652
rect 169352 169640 169358 169652
rect 214006 169640 214012 169652
rect 169352 169612 214012 169640
rect 169352 169600 169358 169612
rect 214006 169600 214012 169612
rect 214064 169600 214070 169652
rect 252462 169600 252468 169652
rect 252520 169640 252526 169652
rect 261018 169640 261024 169652
rect 252520 169612 261024 169640
rect 252520 169600 252526 169612
rect 261018 169600 261024 169612
rect 261076 169600 261082 169652
rect 324314 168988 324320 169040
rect 324372 169028 324378 169040
rect 327258 169028 327264 169040
rect 324372 169000 327264 169028
rect 324372 168988 324378 169000
rect 327258 168988 327264 169000
rect 327316 169028 327322 169040
rect 331950 169028 331956 169040
rect 327316 169000 331956 169028
rect 327316 168988 327322 169000
rect 331950 168988 331956 169000
rect 332008 168988 332014 169040
rect 279418 168444 279424 168496
rect 279476 168484 279482 168496
rect 306742 168484 306748 168496
rect 279476 168456 306748 168484
rect 279476 168444 279482 168456
rect 306742 168444 306748 168456
rect 306800 168444 306806 168496
rect 258902 168376 258908 168428
rect 258960 168416 258966 168428
rect 307294 168416 307300 168428
rect 258960 168388 307300 168416
rect 258960 168376 258966 168388
rect 307294 168376 307300 168388
rect 307352 168376 307358 168428
rect 166534 168308 166540 168360
rect 166592 168348 166598 168360
rect 213914 168348 213920 168360
rect 166592 168320 213920 168348
rect 166592 168308 166598 168320
rect 213914 168308 213920 168320
rect 213972 168308 213978 168360
rect 252370 168308 252376 168360
rect 252428 168348 252434 168360
rect 262398 168348 262404 168360
rect 252428 168320 262404 168348
rect 252428 168308 252434 168320
rect 262398 168308 262404 168320
rect 262456 168308 262462 168360
rect 324314 168308 324320 168360
rect 324372 168348 324378 168360
rect 380894 168348 380900 168360
rect 324372 168320 380900 168348
rect 324372 168308 324378 168320
rect 380894 168308 380900 168320
rect 380952 168308 380958 168360
rect 211982 168240 211988 168292
rect 212040 168280 212046 168292
rect 214006 168280 214012 168292
rect 212040 168252 214012 168280
rect 212040 168240 212046 168252
rect 214006 168240 214012 168252
rect 214064 168240 214070 168292
rect 324406 168240 324412 168292
rect 324464 168280 324470 168292
rect 324682 168280 324688 168292
rect 324464 168252 324688 168280
rect 324464 168240 324470 168252
rect 324682 168240 324688 168252
rect 324740 168280 324746 168292
rect 376018 168280 376024 168292
rect 324740 168252 376024 168280
rect 324740 168240 324746 168252
rect 376018 168240 376024 168252
rect 376076 168240 376082 168292
rect 252462 168172 252468 168224
rect 252520 168212 252526 168224
rect 256970 168212 256976 168224
rect 252520 168184 256976 168212
rect 252520 168172 252526 168184
rect 256970 168172 256976 168184
rect 257028 168172 257034 168224
rect 271230 167628 271236 167680
rect 271288 167668 271294 167680
rect 307570 167668 307576 167680
rect 271288 167640 307576 167668
rect 271288 167628 271294 167640
rect 307570 167628 307576 167640
rect 307628 167628 307634 167680
rect 252462 167220 252468 167272
rect 252520 167260 252526 167272
rect 258166 167260 258172 167272
rect 252520 167232 258172 167260
rect 252520 167220 252526 167232
rect 258166 167220 258172 167232
rect 258224 167220 258230 167272
rect 279602 167084 279608 167136
rect 279660 167124 279666 167136
rect 307662 167124 307668 167136
rect 279660 167096 307668 167124
rect 279660 167084 279666 167096
rect 307662 167084 307668 167096
rect 307720 167084 307726 167136
rect 262950 167016 262956 167068
rect 263008 167056 263014 167068
rect 307478 167056 307484 167068
rect 263008 167028 307484 167056
rect 263008 167016 263014 167028
rect 307478 167016 307484 167028
rect 307536 167016 307542 167068
rect 166626 166948 166632 167000
rect 166684 166988 166690 167000
rect 214098 166988 214104 167000
rect 166684 166960 214104 166988
rect 166684 166948 166690 166960
rect 214098 166948 214104 166960
rect 214156 166948 214162 167000
rect 252462 166948 252468 167000
rect 252520 166988 252526 167000
rect 258258 166988 258264 167000
rect 252520 166960 258264 166988
rect 252520 166948 252526 166960
rect 258258 166948 258264 166960
rect 258316 166948 258322 167000
rect 324314 166948 324320 167000
rect 324372 166988 324378 167000
rect 344278 166988 344284 167000
rect 324372 166960 344284 166988
rect 324372 166948 324378 166960
rect 344278 166948 344284 166960
rect 344336 166948 344342 167000
rect 169202 166880 169208 166932
rect 169260 166920 169266 166932
rect 214006 166920 214012 166932
rect 169260 166892 214012 166920
rect 169260 166880 169266 166892
rect 214006 166880 214012 166892
rect 214064 166880 214070 166932
rect 170674 166812 170680 166864
rect 170732 166852 170738 166864
rect 213914 166852 213920 166864
rect 170732 166824 213920 166852
rect 170732 166812 170738 166824
rect 213914 166812 213920 166824
rect 213972 166812 213978 166864
rect 252370 166812 252376 166864
rect 252428 166852 252434 166864
rect 256786 166852 256792 166864
rect 252428 166824 256792 166852
rect 252428 166812 252434 166824
rect 256786 166812 256792 166824
rect 256844 166812 256850 166864
rect 252278 166268 252284 166320
rect 252336 166308 252342 166320
rect 259546 166308 259552 166320
rect 252336 166280 259552 166308
rect 252336 166268 252342 166280
rect 259546 166268 259552 166280
rect 259604 166268 259610 166320
rect 337470 166268 337476 166320
rect 337528 166308 337534 166320
rect 386874 166308 386880 166320
rect 337528 166280 386880 166308
rect 337528 166268 337534 166280
rect 386874 166268 386880 166280
rect 386932 166268 386938 166320
rect 278222 165724 278228 165776
rect 278280 165764 278286 165776
rect 306558 165764 306564 165776
rect 278280 165736 306564 165764
rect 278280 165724 278286 165736
rect 306558 165724 306564 165736
rect 306616 165724 306622 165776
rect 268562 165656 268568 165708
rect 268620 165696 268626 165708
rect 307662 165696 307668 165708
rect 268620 165668 307668 165696
rect 268620 165656 268626 165668
rect 307662 165656 307668 165668
rect 307720 165656 307726 165708
rect 257522 165588 257528 165640
rect 257580 165628 257586 165640
rect 307478 165628 307484 165640
rect 257580 165600 307484 165628
rect 257580 165588 257586 165600
rect 307478 165588 307484 165600
rect 307536 165588 307542 165640
rect 572346 165588 572352 165640
rect 572404 165628 572410 165640
rect 574094 165628 574100 165640
rect 572404 165600 574100 165628
rect 572404 165588 572410 165600
rect 574094 165588 574100 165600
rect 574152 165588 574158 165640
rect 170490 165520 170496 165572
rect 170548 165560 170554 165572
rect 213914 165560 213920 165572
rect 170548 165532 213920 165560
rect 170548 165520 170554 165532
rect 213914 165520 213920 165532
rect 213972 165520 213978 165572
rect 252462 165520 252468 165572
rect 252520 165560 252526 165572
rect 264974 165560 264980 165572
rect 252520 165532 264980 165560
rect 252520 165520 252526 165532
rect 264974 165520 264980 165532
rect 265032 165520 265038 165572
rect 252462 164976 252468 165028
rect 252520 165016 252526 165028
rect 259730 165016 259736 165028
rect 252520 164988 259736 165016
rect 252520 164976 252526 164988
rect 259730 164976 259736 164988
rect 259788 164976 259794 165028
rect 264422 164840 264428 164892
rect 264480 164880 264486 164892
rect 307294 164880 307300 164892
rect 264480 164852 307300 164880
rect 264480 164840 264486 164852
rect 307294 164840 307300 164852
rect 307352 164840 307358 164892
rect 292022 164296 292028 164348
rect 292080 164336 292086 164348
rect 307570 164336 307576 164348
rect 292080 164308 307576 164336
rect 292080 164296 292086 164308
rect 307570 164296 307576 164308
rect 307628 164296 307634 164348
rect 324314 164296 324320 164348
rect 324372 164336 324378 164348
rect 337378 164336 337384 164348
rect 324372 164308 337384 164336
rect 324372 164296 324378 164308
rect 337378 164296 337384 164308
rect 337436 164296 337442 164348
rect 275278 164228 275284 164280
rect 275336 164268 275342 164280
rect 307662 164268 307668 164280
rect 275336 164240 307668 164268
rect 275336 164228 275342 164240
rect 307662 164228 307668 164240
rect 307720 164228 307726 164280
rect 323394 164228 323400 164280
rect 323452 164268 323458 164280
rect 380250 164268 380256 164280
rect 323452 164240 380256 164268
rect 323452 164228 323458 164240
rect 380250 164228 380256 164240
rect 380308 164228 380314 164280
rect 167730 164160 167736 164212
rect 167788 164200 167794 164212
rect 213914 164200 213920 164212
rect 167788 164172 213920 164200
rect 167788 164160 167794 164172
rect 213914 164160 213920 164172
rect 213972 164160 213978 164212
rect 252186 164160 252192 164212
rect 252244 164200 252250 164212
rect 262306 164200 262312 164212
rect 252244 164172 262312 164200
rect 252244 164160 252250 164172
rect 262306 164160 262312 164172
rect 262364 164160 262370 164212
rect 324314 164160 324320 164212
rect 324372 164200 324378 164212
rect 333238 164200 333244 164212
rect 324372 164172 333244 164200
rect 324372 164160 324378 164172
rect 333238 164160 333244 164172
rect 333296 164160 333302 164212
rect 210418 164092 210424 164144
rect 210476 164132 210482 164144
rect 214006 164132 214012 164144
rect 210476 164104 214012 164132
rect 210476 164092 210482 164104
rect 214006 164092 214012 164104
rect 214064 164092 214070 164144
rect 324406 164092 324412 164144
rect 324464 164132 324470 164144
rect 330570 164132 330576 164144
rect 324464 164104 330576 164132
rect 324464 164092 324470 164104
rect 330570 164092 330576 164104
rect 330628 164092 330634 164144
rect 260374 163480 260380 163532
rect 260432 163520 260438 163532
rect 307386 163520 307392 163532
rect 260432 163492 307392 163520
rect 260432 163480 260438 163492
rect 307386 163480 307392 163492
rect 307444 163480 307450 163532
rect 289262 162936 289268 162988
rect 289320 162976 289326 162988
rect 307478 162976 307484 162988
rect 289320 162948 307484 162976
rect 289320 162936 289326 162948
rect 307478 162936 307484 162948
rect 307536 162936 307542 162988
rect 261478 162868 261484 162920
rect 261536 162908 261542 162920
rect 307662 162908 307668 162920
rect 261536 162880 307668 162908
rect 261536 162868 261542 162880
rect 307662 162868 307668 162880
rect 307720 162868 307726 162920
rect 167822 162800 167828 162852
rect 167880 162840 167886 162852
rect 213914 162840 213920 162852
rect 167880 162812 213920 162840
rect 167880 162800 167886 162812
rect 213914 162800 213920 162812
rect 213972 162800 213978 162852
rect 252094 162800 252100 162852
rect 252152 162840 252158 162852
rect 265158 162840 265164 162852
rect 252152 162812 265164 162840
rect 252152 162800 252158 162812
rect 265158 162800 265164 162812
rect 265216 162800 265222 162852
rect 380434 162800 380440 162852
rect 380492 162840 380498 162852
rect 386874 162840 386880 162852
rect 380492 162812 386880 162840
rect 380492 162800 380498 162812
rect 386874 162800 386880 162812
rect 386932 162800 386938 162852
rect 252462 162732 252468 162784
rect 252520 162772 252526 162784
rect 263686 162772 263692 162784
rect 252520 162744 263692 162772
rect 252520 162732 252526 162744
rect 263686 162732 263692 162744
rect 263744 162732 263750 162784
rect 260834 162120 260840 162172
rect 260892 162160 260898 162172
rect 284938 162160 284944 162172
rect 260892 162132 284944 162160
rect 260892 162120 260898 162132
rect 284938 162120 284944 162132
rect 284996 162120 285002 162172
rect 325878 162120 325884 162172
rect 325936 162160 325942 162172
rect 369210 162160 369216 162172
rect 325936 162132 369216 162160
rect 325936 162120 325942 162132
rect 369210 162120 369216 162132
rect 369268 162120 369274 162172
rect 251542 162052 251548 162104
rect 251600 162092 251606 162104
rect 252830 162092 252836 162104
rect 251600 162064 252836 162092
rect 251600 162052 251606 162064
rect 252830 162052 252836 162064
rect 252888 162052 252894 162104
rect 287698 161576 287704 161628
rect 287756 161616 287762 161628
rect 306742 161616 306748 161628
rect 287756 161588 306748 161616
rect 287756 161576 287762 161588
rect 306742 161576 306748 161588
rect 306800 161576 306806 161628
rect 281074 161508 281080 161560
rect 281132 161548 281138 161560
rect 307662 161548 307668 161560
rect 281132 161520 307668 161548
rect 281132 161508 281138 161520
rect 307662 161508 307668 161520
rect 307720 161508 307726 161560
rect 260098 161440 260104 161492
rect 260156 161480 260162 161492
rect 307478 161480 307484 161492
rect 260156 161452 307484 161480
rect 260156 161440 260162 161452
rect 307478 161440 307484 161452
rect 307536 161440 307542 161492
rect 169018 161372 169024 161424
rect 169076 161412 169082 161424
rect 213914 161412 213920 161424
rect 169076 161384 213920 161412
rect 169076 161372 169082 161384
rect 213914 161372 213920 161384
rect 213972 161372 213978 161424
rect 171870 161304 171876 161356
rect 171928 161344 171934 161356
rect 214006 161344 214012 161356
rect 171928 161316 214012 161344
rect 171928 161304 171934 161316
rect 214006 161304 214012 161316
rect 214064 161304 214070 161356
rect 177758 160692 177764 160744
rect 177816 160732 177822 160744
rect 216030 160732 216036 160744
rect 177816 160704 216036 160732
rect 177816 160692 177822 160704
rect 216030 160692 216036 160704
rect 216088 160692 216094 160744
rect 324314 160692 324320 160744
rect 324372 160732 324378 160744
rect 331490 160732 331496 160744
rect 324372 160704 331496 160732
rect 324372 160692 324378 160704
rect 331490 160692 331496 160704
rect 331548 160692 331554 160744
rect 251542 160216 251548 160268
rect 251600 160256 251606 160268
rect 254210 160256 254216 160268
rect 251600 160228 254216 160256
rect 251600 160216 251606 160228
rect 254210 160216 254216 160228
rect 254268 160216 254274 160268
rect 297542 160216 297548 160268
rect 297600 160256 297606 160268
rect 307662 160256 307668 160268
rect 297600 160228 307668 160256
rect 297600 160216 297606 160228
rect 307662 160216 307668 160228
rect 307720 160216 307726 160268
rect 263134 160148 263140 160200
rect 263192 160188 263198 160200
rect 306742 160188 306748 160200
rect 263192 160160 306748 160188
rect 263192 160148 263198 160160
rect 306742 160148 306748 160160
rect 306800 160148 306806 160200
rect 257430 160080 257436 160132
rect 257488 160120 257494 160132
rect 307570 160120 307576 160132
rect 257488 160092 307576 160120
rect 257488 160080 257494 160092
rect 307570 160080 307576 160092
rect 307628 160080 307634 160132
rect 170582 160012 170588 160064
rect 170640 160052 170646 160064
rect 213914 160052 213920 160064
rect 170640 160024 213920 160052
rect 170640 160012 170646 160024
rect 213914 160012 213920 160024
rect 213972 160012 213978 160064
rect 324314 159332 324320 159384
rect 324372 159372 324378 159384
rect 327350 159372 327356 159384
rect 324372 159344 327356 159372
rect 324372 159332 324378 159344
rect 327350 159332 327356 159344
rect 327408 159372 327414 159384
rect 367922 159372 367928 159384
rect 327408 159344 367928 159372
rect 327408 159332 327414 159344
rect 367922 159332 367928 159344
rect 367980 159332 367986 159384
rect 289078 158856 289084 158908
rect 289136 158896 289142 158908
rect 307662 158896 307668 158908
rect 289136 158868 307668 158896
rect 289136 158856 289142 158868
rect 307662 158856 307668 158868
rect 307720 158856 307726 158908
rect 261570 158788 261576 158840
rect 261628 158828 261634 158840
rect 307570 158828 307576 158840
rect 261628 158800 307576 158828
rect 261628 158788 261634 158800
rect 307570 158788 307576 158800
rect 307628 158788 307634 158840
rect 253290 158720 253296 158772
rect 253348 158760 253354 158772
rect 307478 158760 307484 158772
rect 253348 158732 307484 158760
rect 253348 158720 253354 158732
rect 307478 158720 307484 158732
rect 307536 158720 307542 158772
rect 359642 158720 359648 158772
rect 359700 158760 359706 158772
rect 380342 158760 380348 158772
rect 359700 158732 380348 158760
rect 359700 158720 359706 158732
rect 380342 158720 380348 158732
rect 380400 158720 380406 158772
rect 572622 158720 572628 158772
rect 572680 158760 572686 158772
rect 575474 158760 575480 158772
rect 572680 158732 575480 158760
rect 572680 158720 572686 158732
rect 575474 158720 575480 158732
rect 575532 158720 575538 158772
rect 171962 158652 171968 158704
rect 172020 158692 172026 158704
rect 213914 158692 213920 158704
rect 172020 158664 213920 158692
rect 172020 158652 172026 158664
rect 213914 158652 213920 158664
rect 213972 158652 213978 158704
rect 252462 158652 252468 158704
rect 252520 158692 252526 158704
rect 273438 158692 273444 158704
rect 252520 158664 273444 158692
rect 252520 158652 252526 158664
rect 273438 158652 273444 158664
rect 273496 158652 273502 158704
rect 324406 158652 324412 158704
rect 324464 158692 324470 158704
rect 360194 158692 360200 158704
rect 324464 158664 360200 158692
rect 324464 158652 324470 158664
rect 360194 158652 360200 158664
rect 360252 158652 360258 158704
rect 324314 158584 324320 158636
rect 324372 158624 324378 158636
rect 359642 158624 359648 158636
rect 324372 158596 359648 158624
rect 324372 158584 324378 158596
rect 359642 158584 359648 158596
rect 359700 158584 359706 158636
rect 279694 157972 279700 158024
rect 279752 158012 279758 158024
rect 307294 158012 307300 158024
rect 279752 157984 307300 158012
rect 279752 157972 279758 157984
rect 307294 157972 307300 157984
rect 307352 157972 307358 158024
rect 265710 157428 265716 157480
rect 265768 157468 265774 157480
rect 307478 157468 307484 157480
rect 265768 157440 307484 157468
rect 265768 157428 265774 157440
rect 307478 157428 307484 157440
rect 307536 157428 307542 157480
rect 258810 157360 258816 157412
rect 258868 157400 258874 157412
rect 307662 157400 307668 157412
rect 258868 157372 307668 157400
rect 258868 157360 258874 157372
rect 307662 157360 307668 157372
rect 307720 157360 307726 157412
rect 171778 157292 171784 157344
rect 171836 157332 171842 157344
rect 214006 157332 214012 157344
rect 171836 157304 214012 157332
rect 171836 157292 171842 157304
rect 214006 157292 214012 157304
rect 214064 157292 214070 157344
rect 324314 157292 324320 157344
rect 324372 157332 324378 157344
rect 385034 157332 385040 157344
rect 324372 157304 385040 157332
rect 324372 157292 324378 157304
rect 385034 157292 385040 157304
rect 385092 157292 385098 157344
rect 192478 157224 192484 157276
rect 192536 157264 192542 157276
rect 213914 157264 213920 157276
rect 192536 157236 213920 157264
rect 192536 157224 192542 157236
rect 213914 157224 213920 157236
rect 213972 157224 213978 157276
rect 324406 157224 324412 157276
rect 324464 157264 324470 157276
rect 345290 157264 345296 157276
rect 324464 157236 345296 157264
rect 324464 157224 324470 157236
rect 345290 157224 345296 157236
rect 345348 157264 345354 157276
rect 346302 157264 346308 157276
rect 345348 157236 346308 157264
rect 345348 157224 345354 157236
rect 346302 157224 346308 157236
rect 346360 157224 346366 157276
rect 251174 157088 251180 157140
rect 251232 157128 251238 157140
rect 254026 157128 254032 157140
rect 251232 157100 254032 157128
rect 251232 157088 251238 157100
rect 254026 157088 254032 157100
rect 254084 157088 254090 157140
rect 251358 157020 251364 157072
rect 251416 157060 251422 157072
rect 254118 157060 254124 157072
rect 251416 157032 254124 157060
rect 251416 157020 251422 157032
rect 254118 157020 254124 157032
rect 254176 157020 254182 157072
rect 290642 156612 290648 156664
rect 290700 156652 290706 156664
rect 307570 156652 307576 156664
rect 290700 156624 307576 156652
rect 290700 156612 290706 156624
rect 307570 156612 307576 156624
rect 307628 156612 307634 156664
rect 346302 156612 346308 156664
rect 346360 156652 346366 156664
rect 377490 156652 377496 156664
rect 346360 156624 377496 156652
rect 346360 156612 346366 156624
rect 377490 156612 377496 156624
rect 377548 156612 377554 156664
rect 266998 156000 267004 156052
rect 267056 156040 267062 156052
rect 307662 156040 307668 156052
rect 267056 156012 307668 156040
rect 267056 156000 267062 156012
rect 307662 156000 307668 156012
rect 307720 156000 307726 156052
rect 257614 155932 257620 155984
rect 257672 155972 257678 155984
rect 306742 155972 306748 155984
rect 257672 155944 306748 155972
rect 257672 155932 257678 155944
rect 306742 155932 306748 155944
rect 306800 155932 306806 155984
rect 170398 155864 170404 155916
rect 170456 155904 170462 155916
rect 213914 155904 213920 155916
rect 170456 155876 213920 155904
rect 170456 155864 170462 155876
rect 213914 155864 213920 155876
rect 213972 155864 213978 155916
rect 251818 155864 251824 155916
rect 251876 155904 251882 155916
rect 277394 155904 277400 155916
rect 251876 155876 277400 155904
rect 251876 155864 251882 155876
rect 277394 155864 277400 155876
rect 277452 155864 277458 155916
rect 324314 155864 324320 155916
rect 324372 155904 324378 155916
rect 342438 155904 342444 155916
rect 324372 155876 342444 155904
rect 324372 155864 324378 155876
rect 342438 155864 342444 155876
rect 342496 155864 342502 155916
rect 252462 155796 252468 155848
rect 252520 155836 252526 155848
rect 267734 155836 267740 155848
rect 252520 155808 267740 155836
rect 252520 155796 252526 155808
rect 267734 155796 267740 155808
rect 267792 155796 267798 155848
rect 252370 155728 252376 155780
rect 252428 155768 252434 155780
rect 263594 155768 263600 155780
rect 252428 155740 263600 155768
rect 252428 155728 252434 155740
rect 263594 155728 263600 155740
rect 263652 155728 263658 155780
rect 252278 155252 252284 155304
rect 252336 155292 252342 155304
rect 266538 155292 266544 155304
rect 252336 155264 266544 155292
rect 252336 155252 252342 155264
rect 266538 155252 266544 155264
rect 266596 155252 266602 155304
rect 287882 155252 287888 155304
rect 287940 155292 287946 155304
rect 306926 155292 306932 155304
rect 287940 155264 306932 155292
rect 287940 155252 287946 155264
rect 306926 155252 306932 155264
rect 306984 155252 306990 155304
rect 264974 155184 264980 155236
rect 265032 155224 265038 155236
rect 293126 155224 293132 155236
rect 265032 155196 293132 155224
rect 265032 155184 265038 155196
rect 293126 155184 293132 155196
rect 293184 155184 293190 155236
rect 342438 155184 342444 155236
rect 342496 155224 342502 155236
rect 384390 155224 384396 155236
rect 342496 155196 384396 155224
rect 342496 155184 342502 155196
rect 384390 155184 384396 155196
rect 384448 155184 384454 155236
rect 574738 155184 574744 155236
rect 574796 155224 574802 155236
rect 580350 155224 580356 155236
rect 574796 155196 580356 155224
rect 574796 155184 574802 155196
rect 580350 155184 580356 155196
rect 580408 155184 580414 155236
rect 300210 154640 300216 154692
rect 300268 154680 300274 154692
rect 307662 154680 307668 154692
rect 300268 154652 307668 154680
rect 300268 154640 300274 154652
rect 307662 154640 307668 154652
rect 307720 154640 307726 154692
rect 260282 154572 260288 154624
rect 260340 154612 260346 154624
rect 307478 154612 307484 154624
rect 260340 154584 307484 154612
rect 260340 154572 260346 154584
rect 307478 154572 307484 154584
rect 307536 154572 307542 154624
rect 252462 154504 252468 154556
rect 252520 154544 252526 154556
rect 269298 154544 269304 154556
rect 252520 154516 269304 154544
rect 252520 154504 252526 154516
rect 269298 154504 269304 154516
rect 269356 154504 269362 154556
rect 324314 154504 324320 154556
rect 324372 154544 324378 154556
rect 346486 154544 346492 154556
rect 324372 154516 346492 154544
rect 324372 154504 324378 154516
rect 346486 154504 346492 154516
rect 346544 154544 346550 154556
rect 347682 154544 347688 154556
rect 346544 154516 347688 154544
rect 346544 154504 346550 154516
rect 347682 154504 347688 154516
rect 347740 154504 347746 154556
rect 324406 154436 324412 154488
rect 324464 154476 324470 154488
rect 334250 154476 334256 154488
rect 324464 154448 334256 154476
rect 324464 154436 324470 154448
rect 334250 154436 334256 154448
rect 334308 154476 334314 154488
rect 334618 154476 334624 154488
rect 334308 154448 334624 154476
rect 334308 154436 334314 154448
rect 334618 154436 334624 154448
rect 334676 154436 334682 154488
rect 252094 154300 252100 154352
rect 252152 154340 252158 154352
rect 257338 154340 257344 154352
rect 252152 154312 257344 154340
rect 252152 154300 252158 154312
rect 257338 154300 257344 154312
rect 257396 154300 257402 154352
rect 347682 153892 347688 153944
rect 347740 153932 347746 153944
rect 360930 153932 360936 153944
rect 347740 153904 360936 153932
rect 347740 153892 347746 153904
rect 360930 153892 360936 153904
rect 360988 153892 360994 153944
rect 276014 153824 276020 153876
rect 276072 153864 276078 153876
rect 291930 153864 291936 153876
rect 276072 153836 291936 153864
rect 276072 153824 276078 153836
rect 291930 153824 291936 153836
rect 291988 153824 291994 153876
rect 334618 153824 334624 153876
rect 334676 153864 334682 153876
rect 385770 153864 385776 153876
rect 334676 153836 385776 153864
rect 334676 153824 334682 153836
rect 385770 153824 385776 153836
rect 385828 153824 385834 153876
rect 575382 153824 575388 153876
rect 575440 153864 575446 153876
rect 580994 153864 581000 153876
rect 575440 153836 581000 153864
rect 575440 153824 575446 153836
rect 580994 153824 581000 153836
rect 581052 153824 581058 153876
rect 296254 153348 296260 153400
rect 296312 153388 296318 153400
rect 307662 153388 307668 153400
rect 296312 153360 307668 153388
rect 296312 153348 296318 153360
rect 307662 153348 307668 153360
rect 307720 153348 307726 153400
rect 192478 153280 192484 153332
rect 192536 153320 192542 153332
rect 213914 153320 213920 153332
rect 192536 153292 213920 153320
rect 192536 153280 192542 153292
rect 213914 153280 213920 153292
rect 213972 153280 213978 153332
rect 264330 153280 264336 153332
rect 264388 153320 264394 153332
rect 307570 153320 307576 153332
rect 264388 153292 307576 153320
rect 264388 153280 264394 153292
rect 307570 153280 307576 153292
rect 307628 153280 307634 153332
rect 177298 153212 177304 153264
rect 177356 153252 177362 153264
rect 214006 153252 214012 153264
rect 177356 153224 214012 153252
rect 177356 153212 177362 153224
rect 214006 153212 214012 153224
rect 214064 153212 214070 153264
rect 258718 153212 258724 153264
rect 258776 153252 258782 153264
rect 306558 153252 306564 153264
rect 258776 153224 306564 153252
rect 258776 153212 258782 153224
rect 306558 153212 306564 153224
rect 306616 153212 306622 153264
rect 324958 153212 324964 153264
rect 325016 153252 325022 153264
rect 376018 153252 376024 153264
rect 325016 153224 376024 153252
rect 325016 153212 325022 153224
rect 376018 153212 376024 153224
rect 376076 153212 376082 153264
rect 572622 153212 572628 153264
rect 572680 153252 572686 153264
rect 575382 153252 575388 153264
rect 572680 153224 575388 153252
rect 572680 153212 572686 153224
rect 575382 153212 575388 153224
rect 575440 153212 575446 153264
rect 252370 153144 252376 153196
rect 252428 153184 252434 153196
rect 272058 153184 272064 153196
rect 252428 153156 272064 153184
rect 252428 153144 252434 153156
rect 272058 153144 272064 153156
rect 272116 153144 272122 153196
rect 349798 153144 349804 153196
rect 349856 153184 349862 153196
rect 386874 153184 386880 153196
rect 349856 153156 386880 153184
rect 349856 153144 349862 153156
rect 386874 153144 386880 153156
rect 386932 153144 386938 153196
rect 252462 153076 252468 153128
rect 252520 153116 252526 153128
rect 270494 153116 270500 153128
rect 252520 153088 270500 153116
rect 252520 153076 252526 153088
rect 270494 153076 270500 153088
rect 270552 153076 270558 153128
rect 254578 153008 254584 153060
rect 254636 153048 254642 153060
rect 255406 153048 255412 153060
rect 254636 153020 255412 153048
rect 254636 153008 254642 153020
rect 255406 153008 255412 153020
rect 255464 153008 255470 153060
rect 256234 152464 256240 152516
rect 256292 152504 256298 152516
rect 304994 152504 305000 152516
rect 256292 152476 305000 152504
rect 256292 152464 256298 152476
rect 304994 152464 305000 152476
rect 305052 152464 305058 152516
rect 273990 151920 273996 151972
rect 274048 151960 274054 151972
rect 307662 151960 307668 151972
rect 274048 151932 307668 151960
rect 274048 151920 274054 151932
rect 307662 151920 307668 151932
rect 307720 151920 307726 151972
rect 202230 151852 202236 151904
rect 202288 151892 202294 151904
rect 213914 151892 213920 151904
rect 202288 151864 213920 151892
rect 202288 151852 202294 151864
rect 213914 151852 213920 151864
rect 213972 151852 213978 151904
rect 257338 151852 257344 151904
rect 257396 151892 257402 151904
rect 306558 151892 306564 151904
rect 257396 151864 306564 151892
rect 257396 151852 257402 151864
rect 306558 151852 306564 151864
rect 306616 151852 306622 151904
rect 171778 151784 171784 151836
rect 171836 151824 171842 151836
rect 214006 151824 214012 151836
rect 171836 151796 214012 151824
rect 171836 151784 171842 151796
rect 214006 151784 214012 151796
rect 214064 151784 214070 151836
rect 254118 151784 254124 151836
rect 254176 151824 254182 151836
rect 307570 151824 307576 151836
rect 254176 151796 307576 151824
rect 254176 151784 254182 151796
rect 307570 151784 307576 151796
rect 307628 151784 307634 151836
rect 252462 151716 252468 151768
rect 252520 151756 252526 151768
rect 273254 151756 273260 151768
rect 252520 151728 273260 151756
rect 252520 151716 252526 151728
rect 273254 151716 273260 151728
rect 273312 151716 273318 151768
rect 324314 151716 324320 151768
rect 324372 151756 324378 151768
rect 337470 151756 337476 151768
rect 324372 151728 337476 151756
rect 324372 151716 324378 151728
rect 337470 151716 337476 151728
rect 337528 151716 337534 151768
rect 251910 151648 251916 151700
rect 251968 151688 251974 151700
rect 266446 151688 266452 151700
rect 251968 151660 266452 151688
rect 251968 151648 251974 151660
rect 266446 151648 266452 151660
rect 266504 151648 266510 151700
rect 167638 151036 167644 151088
rect 167696 151076 167702 151088
rect 205634 151076 205640 151088
rect 167696 151048 205640 151076
rect 167696 151036 167702 151048
rect 205634 151036 205640 151048
rect 205692 151036 205698 151088
rect 250622 151036 250628 151088
rect 250680 151076 250686 151088
rect 259454 151076 259460 151088
rect 250680 151048 259460 151076
rect 250680 151036 250686 151048
rect 259454 151036 259460 151048
rect 259512 151036 259518 151088
rect 572622 151036 572628 151088
rect 572680 151076 572686 151088
rect 579614 151076 579620 151088
rect 572680 151048 579620 151076
rect 572680 151036 572686 151048
rect 579614 151036 579620 151048
rect 579672 151036 579678 151088
rect 304350 150560 304356 150612
rect 304408 150600 304414 150612
rect 307662 150600 307668 150612
rect 304408 150572 307668 150600
rect 304408 150560 304414 150572
rect 307662 150560 307668 150572
rect 307720 150560 307726 150612
rect 211890 150492 211896 150544
rect 211948 150532 211954 150544
rect 214006 150532 214012 150544
rect 211948 150504 214012 150532
rect 211948 150492 211954 150504
rect 214006 150492 214012 150504
rect 214064 150492 214070 150544
rect 289354 150492 289360 150544
rect 289412 150532 289418 150544
rect 307478 150532 307484 150544
rect 289412 150504 307484 150532
rect 289412 150492 289418 150504
rect 307478 150492 307484 150504
rect 307536 150492 307542 150544
rect 203610 150424 203616 150476
rect 203668 150464 203674 150476
rect 213914 150464 213920 150476
rect 203668 150436 213920 150464
rect 203668 150424 203674 150436
rect 213914 150424 213920 150436
rect 213972 150424 213978 150476
rect 256050 150424 256056 150476
rect 256108 150464 256114 150476
rect 307570 150464 307576 150476
rect 256108 150436 307576 150464
rect 256108 150424 256114 150436
rect 307570 150424 307576 150436
rect 307628 150424 307634 150476
rect 324406 150424 324412 150476
rect 324464 150464 324470 150476
rect 333882 150464 333888 150476
rect 324464 150436 333888 150464
rect 324464 150424 324470 150436
rect 333882 150424 333888 150436
rect 333940 150464 333946 150476
rect 335538 150464 335544 150476
rect 333940 150436 335544 150464
rect 333940 150424 333946 150436
rect 335538 150424 335544 150436
rect 335596 150424 335602 150476
rect 579614 150424 579620 150476
rect 579672 150464 579678 150476
rect 580258 150464 580264 150476
rect 579672 150436 580264 150464
rect 579672 150424 579678 150436
rect 580258 150424 580264 150436
rect 580316 150424 580322 150476
rect 166442 150356 166448 150408
rect 166500 150396 166506 150408
rect 214006 150396 214012 150408
rect 166500 150368 214012 150396
rect 166500 150356 166506 150368
rect 214006 150356 214012 150368
rect 214064 150356 214070 150408
rect 324314 150356 324320 150408
rect 324372 150396 324378 150408
rect 331306 150396 331312 150408
rect 324372 150368 331312 150396
rect 324372 150356 324378 150368
rect 331306 150356 331312 150368
rect 331364 150356 331370 150408
rect 334158 150356 334164 150408
rect 334216 150396 334222 150408
rect 386598 150396 386604 150408
rect 334216 150368 386604 150396
rect 334216 150356 334222 150368
rect 386598 150356 386604 150368
rect 386656 150356 386662 150408
rect 205634 150288 205640 150340
rect 205692 150328 205698 150340
rect 213914 150328 213920 150340
rect 205692 150300 213920 150328
rect 205692 150288 205698 150300
rect 213914 150288 213920 150300
rect 213972 150288 213978 150340
rect 324406 150288 324412 150340
rect 324464 150328 324470 150340
rect 338206 150328 338212 150340
rect 324464 150300 338212 150328
rect 324464 150288 324470 150300
rect 338206 150288 338212 150300
rect 338264 150288 338270 150340
rect 251174 150152 251180 150204
rect 251232 150192 251238 150204
rect 253934 150192 253940 150204
rect 251232 150164 253940 150192
rect 251232 150152 251238 150164
rect 253934 150152 253940 150164
rect 253992 150152 253998 150204
rect 295978 149676 295984 149728
rect 296036 149716 296042 149728
rect 307202 149716 307208 149728
rect 296036 149688 307208 149716
rect 296036 149676 296042 149688
rect 307202 149676 307208 149688
rect 307260 149676 307266 149728
rect 338206 149676 338212 149728
rect 338264 149716 338270 149728
rect 388438 149716 388444 149728
rect 338264 149688 388444 149716
rect 338264 149676 338270 149688
rect 388438 149676 388444 149688
rect 388496 149676 388502 149728
rect 260190 149064 260196 149116
rect 260248 149104 260254 149116
rect 307478 149104 307484 149116
rect 260248 149076 307484 149104
rect 260248 149064 260254 149076
rect 307478 149064 307484 149076
rect 307536 149064 307542 149116
rect 329190 149064 329196 149116
rect 329248 149104 329254 149116
rect 334158 149104 334164 149116
rect 329248 149076 334164 149104
rect 329248 149064 329254 149076
rect 334158 149064 334164 149076
rect 334216 149064 334222 149116
rect 166258 148996 166264 149048
rect 166316 149036 166322 149048
rect 213914 149036 213920 149048
rect 166316 149008 213920 149036
rect 166316 148996 166322 149008
rect 213914 148996 213920 149008
rect 213972 148996 213978 149048
rect 252462 148996 252468 149048
rect 252520 149036 252526 149048
rect 278774 149036 278780 149048
rect 252520 149008 278780 149036
rect 252520 148996 252526 149008
rect 278774 148996 278780 149008
rect 278832 148996 278838 149048
rect 177850 148316 177856 148368
rect 177908 148356 177914 148368
rect 216122 148356 216128 148368
rect 177908 148328 216128 148356
rect 177908 148316 177914 148328
rect 216122 148316 216128 148328
rect 216180 148316 216186 148368
rect 272610 147772 272616 147824
rect 272668 147812 272674 147824
rect 307570 147812 307576 147824
rect 272668 147784 307576 147812
rect 272668 147772 272674 147784
rect 307570 147772 307576 147784
rect 307628 147772 307634 147824
rect 269850 147704 269856 147756
rect 269908 147744 269914 147756
rect 307662 147744 307668 147756
rect 269908 147716 307668 147744
rect 269908 147704 269914 147716
rect 307662 147704 307668 147716
rect 307720 147704 307726 147756
rect 254670 147636 254676 147688
rect 254728 147676 254734 147688
rect 307478 147676 307484 147688
rect 254728 147648 307484 147676
rect 254728 147636 254734 147648
rect 307478 147636 307484 147648
rect 307536 147636 307542 147688
rect 322842 147636 322848 147688
rect 322900 147676 322906 147688
rect 382918 147676 382924 147688
rect 322900 147648 382924 147676
rect 322900 147636 322906 147648
rect 382918 147636 382924 147648
rect 382976 147636 382982 147688
rect 252370 147568 252376 147620
rect 252428 147608 252434 147620
rect 281534 147608 281540 147620
rect 252428 147580 281540 147608
rect 252428 147568 252434 147580
rect 281534 147568 281540 147580
rect 281592 147568 281598 147620
rect 324314 147568 324320 147620
rect 324372 147608 324378 147620
rect 335630 147608 335636 147620
rect 324372 147580 335636 147608
rect 324372 147568 324378 147580
rect 335630 147568 335636 147580
rect 335688 147608 335694 147620
rect 380158 147608 380164 147620
rect 335688 147580 380164 147608
rect 335688 147568 335694 147580
rect 380158 147568 380164 147580
rect 380216 147568 380222 147620
rect 252462 147500 252468 147552
rect 252520 147540 252526 147552
rect 277486 147540 277492 147552
rect 252520 147512 277492 147540
rect 252520 147500 252526 147512
rect 277486 147500 277492 147512
rect 277544 147500 277550 147552
rect 251726 147432 251732 147484
rect 251784 147472 251790 147484
rect 255498 147472 255504 147484
rect 251784 147444 255504 147472
rect 251784 147432 251790 147444
rect 255498 147432 255504 147444
rect 255556 147432 255562 147484
rect 571702 147296 571708 147348
rect 571760 147336 571766 147348
rect 574738 147336 574744 147348
rect 571760 147308 574744 147336
rect 571760 147296 571766 147308
rect 574738 147296 574744 147308
rect 574796 147296 574802 147348
rect 251542 146956 251548 147008
rect 251600 146996 251606 147008
rect 265066 146996 265072 147008
rect 251600 146968 265072 146996
rect 251600 146956 251606 146968
rect 265066 146956 265072 146968
rect 265124 146956 265130 147008
rect 256142 146888 256148 146940
rect 256200 146928 256206 146940
rect 306926 146928 306932 146940
rect 256200 146900 306932 146928
rect 256200 146888 256206 146900
rect 306926 146888 306932 146900
rect 306984 146888 306990 146940
rect 301590 146412 301596 146464
rect 301648 146452 301654 146464
rect 307662 146452 307668 146464
rect 301648 146424 307668 146452
rect 301648 146412 301654 146424
rect 307662 146412 307668 146424
rect 307720 146412 307726 146464
rect 185578 146344 185584 146396
rect 185636 146384 185642 146396
rect 213914 146384 213920 146396
rect 185636 146356 213920 146384
rect 185636 146344 185642 146356
rect 213914 146344 213920 146356
rect 213972 146344 213978 146396
rect 283834 146344 283840 146396
rect 283892 146384 283898 146396
rect 307570 146384 307576 146396
rect 283892 146356 307576 146384
rect 283892 146344 283898 146356
rect 307570 146344 307576 146356
rect 307628 146344 307634 146396
rect 166258 146276 166264 146328
rect 166316 146316 166322 146328
rect 214006 146316 214012 146328
rect 166316 146288 214012 146316
rect 166316 146276 166322 146288
rect 214006 146276 214012 146288
rect 214064 146276 214070 146328
rect 263042 146276 263048 146328
rect 263100 146316 263106 146328
rect 307478 146316 307484 146328
rect 263100 146288 307484 146316
rect 263100 146276 263106 146288
rect 307478 146276 307484 146288
rect 307536 146276 307542 146328
rect 252094 146208 252100 146260
rect 252152 146248 252158 146260
rect 274634 146248 274640 146260
rect 252152 146220 274640 146248
rect 252152 146208 252158 146220
rect 274634 146208 274640 146220
rect 274692 146208 274698 146260
rect 342438 146208 342444 146260
rect 342496 146248 342502 146260
rect 387058 146248 387064 146260
rect 342496 146220 387064 146248
rect 342496 146208 342502 146220
rect 387058 146208 387064 146220
rect 387116 146208 387122 146260
rect 252278 146140 252284 146192
rect 252336 146180 252342 146192
rect 258350 146180 258356 146192
rect 252336 146152 258356 146180
rect 252336 146140 252342 146152
rect 258350 146140 258356 146152
rect 258408 146140 258414 146192
rect 330570 145596 330576 145648
rect 330628 145636 330634 145648
rect 342438 145636 342444 145648
rect 330628 145608 342444 145636
rect 330628 145596 330634 145608
rect 342438 145596 342444 145608
rect 342496 145596 342502 145648
rect 193858 145528 193864 145580
rect 193916 145568 193922 145580
rect 214098 145568 214104 145580
rect 193916 145540 214104 145568
rect 193916 145528 193922 145540
rect 214098 145528 214104 145540
rect 214156 145528 214162 145580
rect 324314 145528 324320 145580
rect 324372 145568 324378 145580
rect 336826 145568 336832 145580
rect 324372 145540 336832 145568
rect 324372 145528 324378 145540
rect 336826 145528 336832 145540
rect 336884 145568 336890 145580
rect 337470 145568 337476 145580
rect 336884 145540 337476 145568
rect 336884 145528 336890 145540
rect 337470 145528 337476 145540
rect 337528 145528 337534 145580
rect 254854 145052 254860 145104
rect 254912 145092 254918 145104
rect 306926 145092 306932 145104
rect 254912 145064 306932 145092
rect 254912 145052 254918 145064
rect 306926 145052 306932 145064
rect 306984 145052 306990 145104
rect 204898 144984 204904 145036
rect 204956 145024 204962 145036
rect 214006 145024 214012 145036
rect 204956 144996 214012 145024
rect 204956 144984 204962 144996
rect 214006 144984 214012 144996
rect 214064 144984 214070 145036
rect 255958 144984 255964 145036
rect 256016 145024 256022 145036
rect 306558 145024 306564 145036
rect 256016 144996 306564 145024
rect 256016 144984 256022 144996
rect 306558 144984 306564 144996
rect 306616 144984 306622 145036
rect 167638 144916 167644 144968
rect 167696 144956 167702 144968
rect 213914 144956 213920 144968
rect 167696 144928 213920 144956
rect 167696 144916 167702 144928
rect 213914 144916 213920 144928
rect 213972 144916 213978 144968
rect 373258 144916 373264 144968
rect 373316 144956 373322 144968
rect 386598 144956 386604 144968
rect 373316 144928 386604 144956
rect 373316 144916 373322 144928
rect 386598 144916 386604 144928
rect 386656 144916 386662 144968
rect 251910 144848 251916 144900
rect 251968 144888 251974 144900
rect 270586 144888 270592 144900
rect 251968 144860 270592 144888
rect 251968 144848 251974 144860
rect 270586 144848 270592 144860
rect 270644 144848 270650 144900
rect 324406 144848 324412 144900
rect 324464 144888 324470 144900
rect 330478 144888 330484 144900
rect 324464 144860 330484 144888
rect 324464 144848 324470 144860
rect 330478 144848 330484 144860
rect 330536 144848 330542 144900
rect 252462 144780 252468 144832
rect 252520 144820 252526 144832
rect 262214 144820 262220 144832
rect 252520 144792 262220 144820
rect 252520 144780 252526 144792
rect 262214 144780 262220 144792
rect 262272 144780 262278 144832
rect 324314 144780 324320 144832
rect 324372 144820 324378 144832
rect 327166 144820 327172 144832
rect 324372 144792 327172 144820
rect 324372 144780 324378 144792
rect 327166 144780 327172 144792
rect 327224 144780 327230 144832
rect 274634 144236 274640 144288
rect 274692 144276 274698 144288
rect 295334 144276 295340 144288
rect 274692 144248 295340 144276
rect 274692 144236 274698 144248
rect 295334 144236 295340 144248
rect 295392 144236 295398 144288
rect 254762 144168 254768 144220
rect 254820 144208 254826 144220
rect 307386 144208 307392 144220
rect 254820 144180 307392 144208
rect 254820 144168 254826 144180
rect 307386 144168 307392 144180
rect 307444 144168 307450 144220
rect 328362 144168 328368 144220
rect 328420 144208 328426 144220
rect 339494 144208 339500 144220
rect 328420 144180 339500 144208
rect 328420 144168 328426 144180
rect 339494 144168 339500 144180
rect 339552 144168 339558 144220
rect 212074 143624 212080 143676
rect 212132 143664 212138 143676
rect 214650 143664 214656 143676
rect 212132 143636 214656 143664
rect 212132 143624 212138 143636
rect 214650 143624 214656 143636
rect 214708 143624 214714 143676
rect 298738 143624 298744 143676
rect 298796 143664 298802 143676
rect 306926 143664 306932 143676
rect 298796 143636 306932 143664
rect 298796 143624 298802 143636
rect 306926 143624 306932 143636
rect 306984 143624 306990 143676
rect 189810 143556 189816 143608
rect 189868 143596 189874 143608
rect 213914 143596 213920 143608
rect 189868 143568 213920 143596
rect 189868 143556 189874 143568
rect 213914 143556 213920 143568
rect 213972 143556 213978 143608
rect 293402 143556 293408 143608
rect 293460 143596 293466 143608
rect 307662 143596 307668 143608
rect 293460 143568 307668 143596
rect 293460 143556 293466 143568
rect 307662 143556 307668 143568
rect 307720 143556 307726 143608
rect 572622 143556 572628 143608
rect 572680 143596 572686 143608
rect 575566 143596 575572 143608
rect 572680 143568 575572 143596
rect 572680 143556 572686 143568
rect 575566 143556 575572 143568
rect 575624 143556 575630 143608
rect 252370 143488 252376 143540
rect 252428 143528 252434 143540
rect 274726 143528 274732 143540
rect 252428 143500 274732 143528
rect 252428 143488 252434 143500
rect 274726 143488 274732 143500
rect 274784 143488 274790 143540
rect 324406 143488 324412 143540
rect 324464 143528 324470 143540
rect 332686 143528 332692 143540
rect 324464 143500 332692 143528
rect 324464 143488 324470 143500
rect 332686 143488 332692 143500
rect 332744 143488 332750 143540
rect 338850 143488 338856 143540
rect 338908 143528 338914 143540
rect 385678 143528 385684 143540
rect 338908 143500 385684 143528
rect 338908 143488 338914 143500
rect 385678 143488 385684 143500
rect 385736 143488 385742 143540
rect 252462 143420 252468 143472
rect 252520 143460 252526 143472
rect 269206 143460 269212 143472
rect 252520 143432 269212 143460
rect 252520 143420 252526 143432
rect 269206 143420 269212 143432
rect 269264 143420 269270 143472
rect 324314 143352 324320 143404
rect 324372 143392 324378 143404
rect 326338 143392 326344 143404
rect 324372 143364 326344 143392
rect 324372 143352 324378 143364
rect 326338 143352 326344 143364
rect 326396 143352 326402 143404
rect 251818 142808 251824 142860
rect 251876 142848 251882 142860
rect 265710 142848 265716 142860
rect 251876 142820 265716 142848
rect 251876 142808 251882 142820
rect 265710 142808 265716 142820
rect 265768 142808 265774 142860
rect 210510 142672 210516 142724
rect 210568 142712 210574 142724
rect 213914 142712 213920 142724
rect 210568 142684 213920 142712
rect 210568 142672 210574 142684
rect 213914 142672 213920 142684
rect 213972 142672 213978 142724
rect 301498 142264 301504 142316
rect 301556 142304 301562 142316
rect 306742 142304 306748 142316
rect 301556 142276 306748 142304
rect 301556 142264 301562 142276
rect 306742 142264 306748 142276
rect 306800 142264 306806 142316
rect 278314 142196 278320 142248
rect 278372 142236 278378 142248
rect 307478 142236 307484 142248
rect 278372 142208 307484 142236
rect 278372 142196 278378 142208
rect 307478 142196 307484 142208
rect 307536 142196 307542 142248
rect 267090 142128 267096 142180
rect 267148 142168 267154 142180
rect 307662 142168 307668 142180
rect 267148 142140 307668 142168
rect 267148 142128 267154 142140
rect 307662 142128 307668 142140
rect 307720 142128 307726 142180
rect 360102 142128 360108 142180
rect 360160 142168 360166 142180
rect 380158 142168 380164 142180
rect 360160 142140 380164 142168
rect 360160 142128 360166 142140
rect 380158 142128 380164 142140
rect 380216 142128 380222 142180
rect 252462 142060 252468 142112
rect 252520 142100 252526 142112
rect 260926 142100 260932 142112
rect 252520 142072 260932 142100
rect 252520 142060 252526 142072
rect 260926 142060 260932 142072
rect 260984 142060 260990 142112
rect 324406 142060 324412 142112
rect 324464 142100 324470 142112
rect 345198 142100 345204 142112
rect 324464 142072 345204 142100
rect 324464 142060 324470 142072
rect 345198 142060 345204 142072
rect 345256 142100 345262 142112
rect 384298 142100 384304 142112
rect 345256 142072 384304 142100
rect 345256 142060 345262 142072
rect 384298 142060 384304 142072
rect 384356 142060 384362 142112
rect 324314 141992 324320 142044
rect 324372 142032 324378 142044
rect 359550 142032 359556 142044
rect 324372 142004 359556 142032
rect 324372 141992 324378 142004
rect 359550 141992 359556 142004
rect 359608 142032 359614 142044
rect 360102 142032 360108 142044
rect 359608 142004 360108 142032
rect 359608 141992 359614 142004
rect 360102 141992 360108 142004
rect 360160 141992 360166 142044
rect 275462 141448 275468 141500
rect 275520 141488 275526 141500
rect 298094 141488 298100 141500
rect 275520 141460 298100 141488
rect 275520 141448 275526 141460
rect 298094 141448 298100 141460
rect 298152 141448 298158 141500
rect 253474 141380 253480 141432
rect 253532 141420 253538 141432
rect 307110 141420 307116 141432
rect 253532 141392 307116 141420
rect 253532 141380 253538 141392
rect 307110 141380 307116 141392
rect 307168 141380 307174 141432
rect 186958 140836 186964 140888
rect 187016 140876 187022 140888
rect 214006 140876 214012 140888
rect 187016 140848 214012 140876
rect 187016 140836 187022 140848
rect 214006 140836 214012 140848
rect 214064 140836 214070 140888
rect 173342 140768 173348 140820
rect 173400 140808 173406 140820
rect 213914 140808 213920 140820
rect 173400 140780 213920 140808
rect 173400 140768 173406 140780
rect 213914 140768 213920 140780
rect 213972 140768 213978 140820
rect 299106 140768 299112 140820
rect 299164 140808 299170 140820
rect 307662 140808 307668 140820
rect 299164 140780 307668 140808
rect 299164 140768 299170 140780
rect 307662 140768 307668 140780
rect 307720 140768 307726 140820
rect 252094 140700 252100 140752
rect 252152 140740 252158 140752
rect 280154 140740 280160 140752
rect 252152 140712 280160 140740
rect 252152 140700 252158 140712
rect 280154 140700 280160 140712
rect 280212 140700 280218 140752
rect 324314 140700 324320 140752
rect 324372 140740 324378 140752
rect 358170 140740 358176 140752
rect 324372 140712 358176 140740
rect 324372 140700 324378 140712
rect 358170 140700 358176 140712
rect 358228 140700 358234 140752
rect 251726 140632 251732 140684
rect 251784 140672 251790 140684
rect 273346 140672 273352 140684
rect 251784 140644 273352 140672
rect 251784 140632 251790 140644
rect 273346 140632 273352 140644
rect 273404 140632 273410 140684
rect 167822 140020 167828 140072
rect 167880 140060 167886 140072
rect 211890 140060 211896 140072
rect 167880 140032 211896 140060
rect 167880 140020 167886 140032
rect 211890 140020 211896 140032
rect 211948 140020 211954 140072
rect 252186 140020 252192 140072
rect 252244 140060 252250 140072
rect 279418 140060 279424 140072
rect 252244 140032 279424 140060
rect 252244 140020 252250 140032
rect 279418 140020 279424 140032
rect 279476 140020 279482 140072
rect 373442 140020 373448 140072
rect 373500 140060 373506 140072
rect 387610 140060 387616 140072
rect 373500 140032 387616 140060
rect 373500 140020 373506 140032
rect 387610 140020 387616 140032
rect 387668 140020 387674 140072
rect 251726 139748 251732 139800
rect 251784 139788 251790 139800
rect 255590 139788 255596 139800
rect 251784 139760 255596 139788
rect 251784 139748 251790 139760
rect 255590 139748 255596 139760
rect 255648 139748 255654 139800
rect 211982 139476 211988 139528
rect 212040 139516 212046 139528
rect 214650 139516 214656 139528
rect 212040 139488 214656 139516
rect 212040 139476 212046 139488
rect 214650 139476 214656 139488
rect 214708 139476 214714 139528
rect 282362 139476 282368 139528
rect 282420 139516 282426 139528
rect 307570 139516 307576 139528
rect 282420 139488 307576 139516
rect 282420 139476 282426 139488
rect 307570 139476 307576 139488
rect 307628 139476 307634 139528
rect 202138 139408 202144 139460
rect 202196 139448 202202 139460
rect 213914 139448 213920 139460
rect 202196 139420 213920 139448
rect 202196 139408 202202 139420
rect 213914 139408 213920 139420
rect 213972 139408 213978 139460
rect 253382 139408 253388 139460
rect 253440 139448 253446 139460
rect 307662 139448 307668 139460
rect 253440 139420 307668 139448
rect 253440 139408 253446 139420
rect 307662 139408 307668 139420
rect 307720 139408 307726 139460
rect 572622 139408 572628 139460
rect 572680 139448 572686 139460
rect 582650 139448 582656 139460
rect 572680 139420 582656 139448
rect 572680 139408 572686 139420
rect 582650 139408 582656 139420
rect 582708 139408 582714 139460
rect 251358 138728 251364 138780
rect 251416 138768 251422 138780
rect 254578 138768 254584 138780
rect 251416 138740 254584 138768
rect 251416 138728 251422 138740
rect 254578 138728 254584 138740
rect 254636 138728 254642 138780
rect 271414 138660 271420 138712
rect 271472 138700 271478 138712
rect 307294 138700 307300 138712
rect 271472 138672 307300 138700
rect 271472 138660 271478 138672
rect 307294 138660 307300 138672
rect 307352 138660 307358 138712
rect 188430 138048 188436 138100
rect 188488 138088 188494 138100
rect 213914 138088 213920 138100
rect 188488 138060 213920 138088
rect 188488 138048 188494 138060
rect 213914 138048 213920 138060
rect 213972 138048 213978 138100
rect 171870 137980 171876 138032
rect 171928 138020 171934 138032
rect 214006 138020 214012 138032
rect 171928 137992 214012 138020
rect 171928 137980 171934 137992
rect 214006 137980 214012 137992
rect 214064 137980 214070 138032
rect 250530 137980 250536 138032
rect 250588 138020 250594 138032
rect 306926 138020 306932 138032
rect 250588 137992 306932 138020
rect 250588 137980 250594 137992
rect 306926 137980 306932 137992
rect 306984 137980 306990 138032
rect 322842 137980 322848 138032
rect 322900 138020 322906 138032
rect 384298 138020 384304 138032
rect 322900 137992 384304 138020
rect 322900 137980 322906 137992
rect 384298 137980 384304 137992
rect 384356 137980 384362 138032
rect 574738 137980 574744 138032
rect 574796 138020 574802 138032
rect 580166 138020 580172 138032
rect 574796 137992 580172 138020
rect 574796 137980 574802 137992
rect 580166 137980 580172 137992
rect 580224 137980 580230 138032
rect 252462 137912 252468 137964
rect 252520 137952 252526 137964
rect 276106 137952 276112 137964
rect 252520 137924 276112 137952
rect 252520 137912 252526 137924
rect 276106 137912 276112 137924
rect 276164 137912 276170 137964
rect 324314 137912 324320 137964
rect 324372 137952 324378 137964
rect 328546 137952 328552 137964
rect 324372 137924 328552 137952
rect 324372 137912 324378 137924
rect 328546 137912 328552 137924
rect 328604 137952 328610 137964
rect 373258 137952 373264 137964
rect 328604 137924 373264 137952
rect 328604 137912 328610 137924
rect 373258 137912 373264 137924
rect 373316 137912 373322 137964
rect 572622 137912 572628 137964
rect 572680 137952 572686 137964
rect 583018 137952 583024 137964
rect 572680 137924 583024 137952
rect 572680 137912 572686 137924
rect 583018 137912 583024 137924
rect 583076 137912 583082 137964
rect 252094 137844 252100 137896
rect 252152 137884 252158 137896
rect 271966 137884 271972 137896
rect 252152 137856 271972 137884
rect 252152 137844 252158 137856
rect 271966 137844 271972 137856
rect 272024 137844 272030 137896
rect 324406 137844 324412 137896
rect 324464 137884 324470 137896
rect 329834 137884 329840 137896
rect 324464 137856 329840 137884
rect 324464 137844 324470 137856
rect 329834 137844 329840 137856
rect 329892 137884 329898 137896
rect 330294 137884 330300 137896
rect 329892 137856 330300 137884
rect 329892 137844 329898 137856
rect 330294 137844 330300 137856
rect 330352 137844 330358 137896
rect 252002 137300 252008 137352
rect 252060 137340 252066 137352
rect 266998 137340 267004 137352
rect 252060 137312 267004 137340
rect 252060 137300 252066 137312
rect 266998 137300 267004 137312
rect 267056 137300 267062 137352
rect 177482 137232 177488 137284
rect 177540 137272 177546 137284
rect 214742 137272 214748 137284
rect 177540 137244 214748 137272
rect 177540 137232 177546 137244
rect 214742 137232 214748 137244
rect 214800 137232 214806 137284
rect 264514 137232 264520 137284
rect 264572 137272 264578 137284
rect 306558 137272 306564 137284
rect 264572 137244 306564 137272
rect 264572 137232 264578 137244
rect 306558 137232 306564 137244
rect 306616 137232 306622 137284
rect 330294 137232 330300 137284
rect 330352 137272 330358 137284
rect 388622 137272 388628 137284
rect 330352 137244 388628 137272
rect 330352 137232 330358 137244
rect 388622 137232 388628 137244
rect 388680 137232 388686 137284
rect 279418 136688 279424 136740
rect 279476 136728 279482 136740
rect 306926 136728 306932 136740
rect 279476 136700 306932 136728
rect 279476 136688 279482 136700
rect 306926 136688 306932 136700
rect 306984 136688 306990 136740
rect 250438 136620 250444 136672
rect 250496 136660 250502 136672
rect 307662 136660 307668 136672
rect 250496 136632 307668 136660
rect 250496 136620 250502 136632
rect 307662 136620 307668 136632
rect 307720 136620 307726 136672
rect 252370 136552 252376 136604
rect 252428 136592 252434 136604
rect 283742 136592 283748 136604
rect 252428 136564 283748 136592
rect 252428 136552 252434 136564
rect 283742 136552 283748 136564
rect 283800 136552 283806 136604
rect 324314 136552 324320 136604
rect 324372 136592 324378 136604
rect 343818 136592 343824 136604
rect 324372 136564 343824 136592
rect 324372 136552 324378 136564
rect 343818 136552 343824 136564
rect 343876 136592 343882 136604
rect 344462 136592 344468 136604
rect 343876 136564 344468 136592
rect 343876 136552 343882 136564
rect 344462 136552 344468 136564
rect 344520 136552 344526 136604
rect 252094 136484 252100 136536
rect 252152 136524 252158 136536
rect 274082 136524 274088 136536
rect 252152 136496 274088 136524
rect 252152 136484 252158 136496
rect 274082 136484 274088 136496
rect 274140 136484 274146 136536
rect 324406 136484 324412 136536
rect 324464 136524 324470 136536
rect 338850 136524 338856 136536
rect 324464 136496 338856 136524
rect 324464 136484 324470 136496
rect 338850 136484 338856 136496
rect 338908 136484 338914 136536
rect 251726 136416 251732 136468
rect 251784 136456 251790 136468
rect 264238 136456 264244 136468
rect 251784 136428 264244 136456
rect 251784 136416 251790 136428
rect 264238 136416 264244 136428
rect 264296 136416 264302 136468
rect 369118 135940 369124 135992
rect 369176 135980 369182 135992
rect 386414 135980 386420 135992
rect 369176 135952 386420 135980
rect 369176 135940 369182 135952
rect 386414 135940 386420 135952
rect 386472 135980 386478 135992
rect 386690 135980 386696 135992
rect 386472 135952 386696 135980
rect 386472 135940 386478 135952
rect 386690 135940 386696 135952
rect 386748 135940 386754 135992
rect 344462 135872 344468 135924
rect 344520 135912 344526 135924
rect 385678 135912 385684 135924
rect 344520 135884 385684 135912
rect 344520 135872 344526 135884
rect 385678 135872 385684 135884
rect 385736 135872 385742 135924
rect 273898 135464 273904 135516
rect 273956 135504 273962 135516
rect 306926 135504 306932 135516
rect 273956 135476 306932 135504
rect 273956 135464 273962 135476
rect 306926 135464 306932 135476
rect 306984 135464 306990 135516
rect 285030 135396 285036 135448
rect 285088 135436 285094 135448
rect 307478 135436 307484 135448
rect 285088 135408 307484 135436
rect 285088 135396 285094 135408
rect 307478 135396 307484 135408
rect 307536 135396 307542 135448
rect 170398 135328 170404 135380
rect 170456 135368 170462 135380
rect 213914 135368 213920 135380
rect 170456 135340 213920 135368
rect 170456 135328 170462 135340
rect 213914 135328 213920 135340
rect 213972 135328 213978 135380
rect 283558 135328 283564 135380
rect 283616 135368 283622 135380
rect 307570 135368 307576 135380
rect 283616 135340 307576 135368
rect 283616 135328 283622 135340
rect 307570 135328 307576 135340
rect 307628 135328 307634 135380
rect 169110 135260 169116 135312
rect 169168 135300 169174 135312
rect 214006 135300 214012 135312
rect 169168 135272 214012 135300
rect 169168 135260 169174 135272
rect 214006 135260 214012 135272
rect 214064 135260 214070 135312
rect 304258 135260 304264 135312
rect 304316 135300 304322 135312
rect 307662 135300 307668 135312
rect 304316 135272 307668 135300
rect 304316 135260 304322 135272
rect 307662 135260 307668 135272
rect 307720 135260 307726 135312
rect 252462 135192 252468 135244
rect 252520 135232 252526 135244
rect 283650 135232 283656 135244
rect 252520 135204 283656 135232
rect 252520 135192 252526 135204
rect 283650 135192 283656 135204
rect 283708 135192 283714 135244
rect 324314 135192 324320 135244
rect 324372 135232 324378 135244
rect 347958 135232 347964 135244
rect 324372 135204 347964 135232
rect 324372 135192 324378 135204
rect 347958 135192 347964 135204
rect 348016 135232 348022 135244
rect 388530 135232 388536 135244
rect 348016 135204 388536 135232
rect 348016 135192 348022 135204
rect 388530 135192 388536 135204
rect 388588 135192 388594 135244
rect 252278 135124 252284 135176
rect 252336 135164 252342 135176
rect 269758 135164 269764 135176
rect 252336 135136 269764 135164
rect 252336 135124 252342 135136
rect 269758 135124 269764 135136
rect 269816 135124 269822 135176
rect 324406 135124 324412 135176
rect 324464 135164 324470 135176
rect 353294 135164 353300 135176
rect 324464 135136 353300 135164
rect 324464 135124 324470 135136
rect 353294 135124 353300 135136
rect 353352 135164 353358 135176
rect 364978 135164 364984 135176
rect 353352 135136 364984 135164
rect 353352 135124 353358 135136
rect 364978 135124 364984 135136
rect 365036 135124 365042 135176
rect 325510 134512 325516 134564
rect 325568 134552 325574 134564
rect 366358 134552 366364 134564
rect 325568 134524 366364 134552
rect 325568 134512 325574 134524
rect 366358 134512 366364 134524
rect 366416 134512 366422 134564
rect 282178 133968 282184 134020
rect 282236 134008 282242 134020
rect 306742 134008 306748 134020
rect 282236 133980 306748 134008
rect 282236 133968 282242 133980
rect 306742 133968 306748 133980
rect 306800 133968 306806 134020
rect 207750 133900 207756 133952
rect 207808 133940 207814 133952
rect 213914 133940 213920 133952
rect 207808 133912 213920 133940
rect 207808 133900 207814 133912
rect 213914 133900 213920 133912
rect 213972 133900 213978 133952
rect 271322 133900 271328 133952
rect 271380 133940 271386 133952
rect 307662 133940 307668 133952
rect 271380 133912 307668 133940
rect 271380 133900 271386 133912
rect 307662 133900 307668 133912
rect 307720 133900 307726 133952
rect 252370 133832 252376 133884
rect 252428 133872 252434 133884
rect 289446 133872 289452 133884
rect 252428 133844 289452 133872
rect 252428 133832 252434 133844
rect 289446 133832 289452 133844
rect 289504 133832 289510 133884
rect 324314 133832 324320 133884
rect 324372 133872 324378 133884
rect 341058 133872 341064 133884
rect 324372 133844 341064 133872
rect 324372 133832 324378 133844
rect 341058 133832 341064 133844
rect 341116 133872 341122 133884
rect 341242 133872 341248 133884
rect 341116 133844 341248 133872
rect 341116 133832 341122 133844
rect 341242 133832 341248 133844
rect 341300 133832 341306 133884
rect 251726 133764 251732 133816
rect 251784 133804 251790 133816
rect 262858 133804 262864 133816
rect 251784 133776 262864 133804
rect 251784 133764 251790 133776
rect 262858 133764 262864 133776
rect 262916 133764 262922 133816
rect 252462 133696 252468 133748
rect 252520 133736 252526 133748
rect 261662 133736 261668 133748
rect 252520 133708 261668 133736
rect 252520 133696 252526 133708
rect 261662 133696 261668 133708
rect 261720 133696 261726 133748
rect 341242 133220 341248 133272
rect 341300 133260 341306 133272
rect 359550 133260 359556 133272
rect 341300 133232 359556 133260
rect 341300 133220 341306 133232
rect 359550 133220 359556 133232
rect 359608 133220 359614 133272
rect 261754 133152 261760 133204
rect 261812 133192 261818 133204
rect 307386 133192 307392 133204
rect 261812 133164 307392 133192
rect 261812 133152 261818 133164
rect 307386 133152 307392 133164
rect 307444 133152 307450 133204
rect 337470 133152 337476 133204
rect 337528 133192 337534 133204
rect 387610 133192 387616 133204
rect 337528 133164 387616 133192
rect 337528 133152 337534 133164
rect 387610 133152 387616 133164
rect 387668 133152 387674 133204
rect 289170 132540 289176 132592
rect 289228 132580 289234 132592
rect 307478 132580 307484 132592
rect 289228 132552 307484 132580
rect 289228 132540 289234 132552
rect 307478 132540 307484 132552
rect 307536 132540 307542 132592
rect 173250 132472 173256 132524
rect 173308 132512 173314 132524
rect 213914 132512 213920 132524
rect 173308 132484 213920 132512
rect 173308 132472 173314 132484
rect 213914 132472 213920 132484
rect 213972 132472 213978 132524
rect 280982 132472 280988 132524
rect 281040 132512 281046 132524
rect 306926 132512 306932 132524
rect 281040 132484 306932 132512
rect 281040 132472 281046 132484
rect 306926 132472 306932 132484
rect 306984 132472 306990 132524
rect 252462 132404 252468 132456
rect 252520 132444 252526 132456
rect 268470 132444 268476 132456
rect 252520 132416 268476 132444
rect 252520 132404 252526 132416
rect 268470 132404 268476 132416
rect 268528 132404 268534 132456
rect 324314 132404 324320 132456
rect 324372 132444 324378 132456
rect 358814 132444 358820 132456
rect 324372 132416 358820 132444
rect 324372 132404 324378 132416
rect 358814 132404 358820 132416
rect 358872 132444 358878 132456
rect 373442 132444 373448 132456
rect 358872 132416 373448 132444
rect 358872 132404 358878 132416
rect 373442 132404 373448 132416
rect 373500 132404 373506 132456
rect 324406 132336 324412 132388
rect 324464 132376 324470 132388
rect 347130 132376 347136 132388
rect 324464 132348 347136 132376
rect 324464 132336 324470 132348
rect 347130 132336 347136 132348
rect 347188 132336 347194 132388
rect 278774 131724 278780 131776
rect 278832 131764 278838 131776
rect 293034 131764 293040 131776
rect 278832 131736 293040 131764
rect 278832 131724 278838 131736
rect 293034 131724 293040 131736
rect 293092 131724 293098 131776
rect 373258 131724 373264 131776
rect 373316 131764 373322 131776
rect 386414 131764 386420 131776
rect 373316 131736 386420 131764
rect 373316 131724 373322 131736
rect 386414 131724 386420 131736
rect 386472 131724 386478 131776
rect 252462 131588 252468 131640
rect 252520 131628 252526 131640
rect 260374 131628 260380 131640
rect 252520 131600 260380 131628
rect 252520 131588 252526 131600
rect 260374 131588 260380 131600
rect 260432 131588 260438 131640
rect 290550 131248 290556 131300
rect 290608 131288 290614 131300
rect 307478 131288 307484 131300
rect 290608 131260 307484 131288
rect 290608 131248 290614 131260
rect 307478 131248 307484 131260
rect 307536 131248 307542 131300
rect 286410 131180 286416 131232
rect 286468 131220 286474 131232
rect 307570 131220 307576 131232
rect 286468 131192 307576 131220
rect 286468 131180 286474 131192
rect 307570 131180 307576 131192
rect 307628 131180 307634 131232
rect 192570 131112 192576 131164
rect 192628 131152 192634 131164
rect 213914 131152 213920 131164
rect 192628 131124 213920 131152
rect 192628 131112 192634 131124
rect 213914 131112 213920 131124
rect 213972 131112 213978 131164
rect 262858 131112 262864 131164
rect 262916 131152 262922 131164
rect 307662 131152 307668 131164
rect 262916 131124 307668 131152
rect 262916 131112 262922 131124
rect 307662 131112 307668 131124
rect 307720 131112 307726 131164
rect 328362 131112 328368 131164
rect 328420 131152 328426 131164
rect 378870 131152 378876 131164
rect 328420 131124 378876 131152
rect 328420 131112 328426 131124
rect 378870 131112 378876 131124
rect 378928 131112 378934 131164
rect 252462 131044 252468 131096
rect 252520 131084 252526 131096
rect 282270 131084 282276 131096
rect 252520 131056 282276 131084
rect 252520 131044 252526 131056
rect 282270 131044 282276 131056
rect 282328 131044 282334 131096
rect 324406 131044 324412 131096
rect 324464 131084 324470 131096
rect 332778 131084 332784 131096
rect 324464 131056 332784 131084
rect 324464 131044 324470 131056
rect 332778 131044 332784 131056
rect 332836 131044 332842 131096
rect 252370 130976 252376 131028
rect 252428 131016 252434 131028
rect 265618 131016 265624 131028
rect 252428 130988 265624 131016
rect 252428 130976 252434 130988
rect 265618 130976 265624 130988
rect 265676 130976 265682 131028
rect 324314 130976 324320 131028
rect 324372 131016 324378 131028
rect 328362 131016 328368 131028
rect 324372 130988 328368 131016
rect 324372 130976 324378 130988
rect 328362 130976 328368 130988
rect 328420 130976 328426 131028
rect 332778 130364 332784 130416
rect 332836 130404 332842 130416
rect 381722 130404 381728 130416
rect 332836 130376 381728 130404
rect 332836 130364 332842 130376
rect 381722 130364 381728 130376
rect 381780 130364 381786 130416
rect 572622 130160 572628 130212
rect 572680 130200 572686 130212
rect 577590 130200 577596 130212
rect 572680 130172 577596 130200
rect 572680 130160 572686 130172
rect 577590 130160 577596 130172
rect 577648 130160 577654 130212
rect 303154 129956 303160 130008
rect 303212 129996 303218 130008
rect 306742 129996 306748 130008
rect 303212 129968 306748 129996
rect 303212 129956 303218 129968
rect 306742 129956 306748 129968
rect 306800 129956 306806 130008
rect 298922 129888 298928 129940
rect 298980 129928 298986 129940
rect 307662 129928 307668 129940
rect 298980 129900 307668 129928
rect 298980 129888 298986 129900
rect 307662 129888 307668 129900
rect 307720 129888 307726 129940
rect 286318 129820 286324 129872
rect 286376 129860 286382 129872
rect 307110 129860 307116 129872
rect 286376 129832 307116 129860
rect 286376 129820 286382 129832
rect 307110 129820 307116 129832
rect 307168 129820 307174 129872
rect 265710 129752 265716 129804
rect 265768 129792 265774 129804
rect 307570 129792 307576 129804
rect 265768 129764 307576 129792
rect 265768 129752 265774 129764
rect 307570 129752 307576 129764
rect 307628 129752 307634 129804
rect 252462 129684 252468 129736
rect 252520 129724 252526 129736
rect 271230 129724 271236 129736
rect 252520 129696 271236 129724
rect 252520 129684 252526 129696
rect 271230 129684 271236 129696
rect 271288 129684 271294 129736
rect 373350 129684 373356 129736
rect 373408 129724 373414 129736
rect 386598 129724 386604 129736
rect 373408 129696 386604 129724
rect 373408 129684 373414 129696
rect 386598 129684 386604 129696
rect 386656 129684 386662 129736
rect 252370 129616 252376 129668
rect 252428 129656 252434 129668
rect 264422 129656 264428 129668
rect 252428 129628 264428 129656
rect 252428 129616 252434 129628
rect 264422 129616 264428 129628
rect 264480 129616 264486 129668
rect 324314 129004 324320 129056
rect 324372 129044 324378 129056
rect 340782 129044 340788 129056
rect 324372 129016 340788 129044
rect 324372 129004 324378 129016
rect 340782 129004 340788 129016
rect 340840 129004 340846 129056
rect 356698 129004 356704 129056
rect 356756 129044 356762 129056
rect 387058 129044 387064 129056
rect 356756 129016 387064 129044
rect 356756 129004 356762 129016
rect 387058 129004 387064 129016
rect 387116 129004 387122 129056
rect 251726 128460 251732 128512
rect 251784 128500 251790 128512
rect 258902 128500 258908 128512
rect 251784 128472 258908 128500
rect 251784 128460 251790 128472
rect 258902 128460 258908 128472
rect 258960 128460 258966 128512
rect 196710 128392 196716 128444
rect 196768 128432 196774 128444
rect 214006 128432 214012 128444
rect 196768 128404 214012 128432
rect 196768 128392 196774 128404
rect 214006 128392 214012 128404
rect 214064 128392 214070 128444
rect 278130 128392 278136 128444
rect 278188 128432 278194 128444
rect 307478 128432 307484 128444
rect 278188 128404 307484 128432
rect 278188 128392 278194 128404
rect 307478 128392 307484 128404
rect 307536 128392 307542 128444
rect 169018 128324 169024 128376
rect 169076 128364 169082 128376
rect 213914 128364 213920 128376
rect 169076 128336 213920 128364
rect 169076 128324 169082 128336
rect 213914 128324 213920 128336
rect 213972 128324 213978 128376
rect 265618 128324 265624 128376
rect 265676 128364 265682 128376
rect 307662 128364 307668 128376
rect 265676 128336 307668 128364
rect 265676 128324 265682 128336
rect 307662 128324 307668 128336
rect 307720 128324 307726 128376
rect 252462 128256 252468 128308
rect 252520 128296 252526 128308
rect 279602 128296 279608 128308
rect 252520 128268 279608 128296
rect 252520 128256 252526 128268
rect 279602 128256 279608 128268
rect 279660 128256 279666 128308
rect 324314 128256 324320 128308
rect 324372 128296 324378 128308
rect 354766 128296 354772 128308
rect 324372 128268 354772 128296
rect 324372 128256 324378 128268
rect 354766 128256 354772 128268
rect 354824 128296 354830 128308
rect 355962 128296 355968 128308
rect 354824 128268 355968 128296
rect 354824 128256 354830 128268
rect 355962 128256 355968 128268
rect 356020 128256 356026 128308
rect 252370 128188 252376 128240
rect 252428 128228 252434 128240
rect 268562 128228 268568 128240
rect 252428 128200 268568 128228
rect 252428 128188 252434 128200
rect 268562 128188 268568 128200
rect 268620 128188 268626 128240
rect 172330 127576 172336 127628
rect 172388 127616 172394 127628
rect 198090 127616 198096 127628
rect 172388 127588 198096 127616
rect 172388 127576 172394 127588
rect 198090 127576 198096 127588
rect 198148 127576 198154 127628
rect 355962 127576 355968 127628
rect 356020 127616 356026 127628
rect 374730 127616 374736 127628
rect 356020 127588 374736 127616
rect 356020 127576 356026 127588
rect 374730 127576 374736 127588
rect 374788 127576 374794 127628
rect 252094 127168 252100 127220
rect 252152 127208 252158 127220
rect 253290 127208 253296 127220
rect 252152 127180 253296 127208
rect 252152 127168 252158 127180
rect 253290 127168 253296 127180
rect 253348 127168 253354 127220
rect 280798 127100 280804 127152
rect 280856 127140 280862 127152
rect 307662 127140 307668 127152
rect 280856 127112 307668 127140
rect 280856 127100 280862 127112
rect 307662 127100 307668 127112
rect 307720 127100 307726 127152
rect 279510 127032 279516 127084
rect 279568 127072 279574 127084
rect 307478 127072 307484 127084
rect 279568 127044 307484 127072
rect 279568 127032 279574 127044
rect 307478 127032 307484 127044
rect 307536 127032 307542 127084
rect 206462 126964 206468 127016
rect 206520 127004 206526 127016
rect 213914 127004 213920 127016
rect 206520 126976 213920 127004
rect 206520 126964 206526 126976
rect 213914 126964 213920 126976
rect 213972 126964 213978 127016
rect 269758 126964 269764 127016
rect 269816 127004 269822 127016
rect 307570 127004 307576 127016
rect 269816 126976 307576 127004
rect 269816 126964 269822 126976
rect 307570 126964 307576 126976
rect 307628 126964 307634 127016
rect 252370 126896 252376 126948
rect 252428 126936 252434 126948
rect 292022 126936 292028 126948
rect 252428 126908 292028 126936
rect 252428 126896 252434 126908
rect 292022 126896 292028 126908
rect 292080 126896 292086 126948
rect 324314 126896 324320 126948
rect 324372 126936 324378 126948
rect 378134 126936 378140 126948
rect 324372 126908 378140 126936
rect 324372 126896 324378 126908
rect 378134 126896 378140 126908
rect 378192 126896 378198 126948
rect 252462 126828 252468 126880
rect 252520 126868 252526 126880
rect 278222 126868 278228 126880
rect 252520 126840 278228 126868
rect 252520 126828 252526 126840
rect 278222 126828 278228 126840
rect 278280 126828 278286 126880
rect 252462 126556 252468 126608
rect 252520 126596 252526 126608
rect 257522 126596 257528 126608
rect 252520 126568 257528 126596
rect 252520 126556 252526 126568
rect 257522 126556 257528 126568
rect 257580 126556 257586 126608
rect 257706 126216 257712 126268
rect 257764 126256 257770 126268
rect 280890 126256 280896 126268
rect 257764 126228 280896 126256
rect 257764 126216 257770 126228
rect 280890 126216 280896 126228
rect 280948 126216 280954 126268
rect 569218 126216 569224 126268
rect 569276 126256 569282 126268
rect 578326 126256 578332 126268
rect 569276 126228 578332 126256
rect 569276 126216 569282 126228
rect 578326 126216 578332 126228
rect 578384 126256 578390 126268
rect 579614 126256 579620 126268
rect 578384 126228 579620 126256
rect 578384 126216 578390 126228
rect 579614 126216 579620 126228
rect 579672 126216 579678 126268
rect 196802 125672 196808 125724
rect 196860 125712 196866 125724
rect 214006 125712 214012 125724
rect 196860 125684 214012 125712
rect 196860 125672 196866 125684
rect 214006 125672 214012 125684
rect 214064 125672 214070 125724
rect 291930 125672 291936 125724
rect 291988 125712 291994 125724
rect 307570 125712 307576 125724
rect 291988 125684 307576 125712
rect 291988 125672 291994 125684
rect 307570 125672 307576 125684
rect 307628 125672 307634 125724
rect 173434 125604 173440 125656
rect 173492 125644 173498 125656
rect 213914 125644 213920 125656
rect 173492 125616 213920 125644
rect 173492 125604 173498 125616
rect 213914 125604 213920 125616
rect 213972 125604 213978 125656
rect 268470 125604 268476 125656
rect 268528 125644 268534 125656
rect 307662 125644 307668 125656
rect 268528 125616 307668 125644
rect 268528 125604 268534 125616
rect 307662 125604 307668 125616
rect 307720 125604 307726 125656
rect 324314 125536 324320 125588
rect 324372 125576 324378 125588
rect 349246 125576 349252 125588
rect 324372 125548 349252 125576
rect 324372 125536 324378 125548
rect 349246 125536 349252 125548
rect 349304 125576 349310 125588
rect 349614 125576 349620 125588
rect 349304 125548 349620 125576
rect 349304 125536 349310 125548
rect 349614 125536 349620 125548
rect 349672 125536 349678 125588
rect 252462 125468 252468 125520
rect 252520 125508 252526 125520
rect 275278 125508 275284 125520
rect 252520 125480 275284 125508
rect 252520 125468 252526 125480
rect 275278 125468 275284 125480
rect 275336 125468 275342 125520
rect 324406 125468 324412 125520
rect 324464 125508 324470 125520
rect 347866 125508 347872 125520
rect 324464 125480 347872 125508
rect 324464 125468 324470 125480
rect 347866 125468 347872 125480
rect 347924 125508 347930 125520
rect 367830 125508 367836 125520
rect 347924 125480 367836 125508
rect 347924 125468 347930 125480
rect 367830 125468 367836 125480
rect 367888 125468 367894 125520
rect 252370 125400 252376 125452
rect 252428 125440 252434 125452
rect 279694 125440 279700 125452
rect 252428 125412 279700 125440
rect 252428 125400 252434 125412
rect 279694 125400 279700 125412
rect 279752 125400 279758 125452
rect 251174 125332 251180 125384
rect 251232 125372 251238 125384
rect 253474 125372 253480 125384
rect 251232 125344 253480 125372
rect 251232 125332 251238 125344
rect 253474 125332 253480 125344
rect 253532 125332 253538 125384
rect 280154 124924 280160 124976
rect 280212 124964 280218 124976
rect 291838 124964 291844 124976
rect 280212 124936 291844 124964
rect 280212 124924 280218 124936
rect 291838 124924 291844 124936
rect 291896 124924 291902 124976
rect 275370 124856 275376 124908
rect 275428 124896 275434 124908
rect 307018 124896 307024 124908
rect 275428 124868 307024 124896
rect 275428 124856 275434 124868
rect 307018 124856 307024 124868
rect 307076 124856 307082 124908
rect 349614 124856 349620 124908
rect 349672 124896 349678 124908
rect 389818 124896 389824 124908
rect 349672 124868 389824 124896
rect 349672 124856 349678 124868
rect 389818 124856 389824 124868
rect 389876 124856 389882 124908
rect 260374 124380 260380 124432
rect 260432 124420 260438 124432
rect 306742 124420 306748 124432
rect 260432 124392 306748 124420
rect 260432 124380 260438 124392
rect 306742 124380 306748 124392
rect 306800 124380 306806 124432
rect 296070 124312 296076 124364
rect 296128 124352 296134 124364
rect 307478 124352 307484 124364
rect 296128 124324 307484 124352
rect 296128 124312 296134 124324
rect 307478 124312 307484 124324
rect 307536 124312 307542 124364
rect 170490 124244 170496 124296
rect 170548 124284 170554 124296
rect 213914 124284 213920 124296
rect 170548 124256 213920 124284
rect 170548 124244 170554 124256
rect 213914 124244 213920 124256
rect 213972 124244 213978 124296
rect 278222 124244 278228 124296
rect 278280 124284 278286 124296
rect 307662 124284 307668 124296
rect 278280 124256 307668 124284
rect 278280 124244 278286 124256
rect 307662 124244 307668 124256
rect 307720 124244 307726 124296
rect 166350 124176 166356 124228
rect 166408 124216 166414 124228
rect 214006 124216 214012 124228
rect 166408 124188 214012 124216
rect 166408 124176 166414 124188
rect 214006 124176 214012 124188
rect 214064 124176 214070 124228
rect 252278 124108 252284 124160
rect 252336 124148 252342 124160
rect 295978 124148 295984 124160
rect 252336 124120 295984 124148
rect 252336 124108 252342 124120
rect 295978 124108 295984 124120
rect 296036 124108 296042 124160
rect 324498 124108 324504 124160
rect 324556 124148 324562 124160
rect 350626 124148 350632 124160
rect 324556 124120 350632 124148
rect 324556 124108 324562 124120
rect 350626 124108 350632 124120
rect 350684 124108 350690 124160
rect 572622 124108 572628 124160
rect 572680 124148 572686 124160
rect 583294 124148 583300 124160
rect 572680 124120 583300 124148
rect 572680 124108 572686 124120
rect 583294 124108 583300 124120
rect 583352 124108 583358 124160
rect 252462 124040 252468 124092
rect 252520 124080 252526 124092
rect 289262 124080 289268 124092
rect 252520 124052 289268 124080
rect 252520 124040 252526 124052
rect 289262 124040 289268 124052
rect 289320 124040 289326 124092
rect 324314 124040 324320 124092
rect 324372 124080 324378 124092
rect 334066 124080 334072 124092
rect 324372 124052 334072 124080
rect 324372 124040 324378 124052
rect 334066 124040 334072 124052
rect 334124 124040 334130 124092
rect 252370 123972 252376 124024
rect 252428 124012 252434 124024
rect 261478 124012 261484 124024
rect 252428 123984 261484 124012
rect 252428 123972 252434 123984
rect 261478 123972 261484 123984
rect 261536 123972 261542 124024
rect 324406 123972 324412 124024
rect 324464 124012 324470 124024
rect 329190 124012 329196 124024
rect 324464 123984 329196 124012
rect 324464 123972 324470 123984
rect 329190 123972 329196 123984
rect 329248 123972 329254 124024
rect 350626 123428 350632 123480
rect 350684 123468 350690 123480
rect 385862 123468 385868 123480
rect 350684 123440 385868 123468
rect 350684 123428 350690 123440
rect 385862 123428 385868 123440
rect 385920 123428 385926 123480
rect 294598 122952 294604 123004
rect 294656 122992 294662 123004
rect 307110 122992 307116 123004
rect 294656 122964 307116 122992
rect 294656 122952 294662 122964
rect 307110 122952 307116 122964
rect 307168 122952 307174 123004
rect 170582 122884 170588 122936
rect 170640 122924 170646 122936
rect 213914 122924 213920 122936
rect 170640 122896 213920 122924
rect 170640 122884 170646 122896
rect 213914 122884 213920 122896
rect 213972 122884 213978 122936
rect 293218 122884 293224 122936
rect 293276 122924 293282 122936
rect 307662 122924 307668 122936
rect 293276 122896 307668 122924
rect 293276 122884 293282 122896
rect 307662 122884 307668 122896
rect 307720 122884 307726 122936
rect 167730 122816 167736 122868
rect 167788 122856 167794 122868
rect 214006 122856 214012 122868
rect 167788 122828 214012 122856
rect 167788 122816 167794 122828
rect 214006 122816 214012 122828
rect 214064 122816 214070 122868
rect 287790 122816 287796 122868
rect 287848 122856 287854 122868
rect 307478 122856 307484 122868
rect 287848 122828 307484 122856
rect 287848 122816 287854 122828
rect 307478 122816 307484 122828
rect 307536 122816 307542 122868
rect 252462 122748 252468 122800
rect 252520 122788 252526 122800
rect 287698 122788 287704 122800
rect 252520 122760 287704 122788
rect 252520 122748 252526 122760
rect 287698 122748 287704 122760
rect 287756 122748 287762 122800
rect 321646 122748 321652 122800
rect 321704 122788 321710 122800
rect 341518 122788 341524 122800
rect 321704 122760 341524 122788
rect 321704 122748 321710 122760
rect 341518 122748 341524 122760
rect 341576 122748 341582 122800
rect 377398 122748 377404 122800
rect 377456 122788 377462 122800
rect 386782 122788 386788 122800
rect 377456 122760 386788 122788
rect 377456 122748 377462 122760
rect 386782 122748 386788 122760
rect 386840 122748 386846 122800
rect 252370 122680 252376 122732
rect 252428 122720 252434 122732
rect 281074 122720 281080 122732
rect 252428 122692 281080 122720
rect 252428 122680 252434 122692
rect 281074 122680 281080 122692
rect 281132 122680 281138 122732
rect 324314 122476 324320 122528
rect 324372 122516 324378 122528
rect 327074 122516 327080 122528
rect 324372 122488 327080 122516
rect 324372 122476 324378 122488
rect 327074 122476 327080 122488
rect 327132 122476 327138 122528
rect 167914 122068 167920 122120
rect 167972 122108 167978 122120
rect 203610 122108 203616 122120
rect 167972 122080 203616 122108
rect 167972 122068 167978 122080
rect 203610 122068 203616 122080
rect 203668 122068 203674 122120
rect 337470 122068 337476 122120
rect 337528 122108 337534 122120
rect 387150 122108 387156 122120
rect 337528 122080 387156 122108
rect 337528 122068 337534 122080
rect 387150 122068 387156 122080
rect 387208 122068 387214 122120
rect 252462 121864 252468 121916
rect 252520 121904 252526 121916
rect 260098 121904 260104 121916
rect 252520 121876 260104 121904
rect 252520 121864 252526 121876
rect 260098 121864 260104 121876
rect 260156 121864 260162 121916
rect 290458 121592 290464 121644
rect 290516 121632 290522 121644
rect 307662 121632 307668 121644
rect 290516 121604 307668 121632
rect 290516 121592 290522 121604
rect 307662 121592 307668 121604
rect 307720 121592 307726 121644
rect 206554 121524 206560 121576
rect 206612 121564 206618 121576
rect 214006 121564 214012 121576
rect 206612 121536 214012 121564
rect 206612 121524 206618 121536
rect 214006 121524 214012 121536
rect 214064 121524 214070 121576
rect 283742 121524 283748 121576
rect 283800 121564 283806 121576
rect 307570 121564 307576 121576
rect 283800 121536 307576 121564
rect 283800 121524 283806 121536
rect 307570 121524 307576 121536
rect 307628 121524 307634 121576
rect 184290 121456 184296 121508
rect 184348 121496 184354 121508
rect 213914 121496 213920 121508
rect 184348 121468 213920 121496
rect 184348 121456 184354 121468
rect 213914 121456 213920 121468
rect 213972 121456 213978 121508
rect 266998 121456 267004 121508
rect 267056 121496 267062 121508
rect 307478 121496 307484 121508
rect 267056 121468 307484 121496
rect 267056 121456 267062 121468
rect 307478 121456 307484 121468
rect 307536 121456 307542 121508
rect 252370 121388 252376 121440
rect 252428 121428 252434 121440
rect 297542 121428 297548 121440
rect 252428 121400 297548 121428
rect 252428 121388 252434 121400
rect 297542 121388 297548 121400
rect 297600 121388 297606 121440
rect 324314 121388 324320 121440
rect 324372 121428 324378 121440
rect 343726 121428 343732 121440
rect 324372 121400 343732 121428
rect 324372 121388 324378 121400
rect 343726 121388 343732 121400
rect 343784 121388 343790 121440
rect 252462 121320 252468 121372
rect 252520 121360 252526 121372
rect 263134 121360 263140 121372
rect 252520 121332 263140 121360
rect 252520 121320 252526 121332
rect 263134 121320 263140 121332
rect 263192 121320 263198 121372
rect 324406 121320 324412 121372
rect 324464 121360 324470 121372
rect 327534 121360 327540 121372
rect 324464 121332 327540 121360
rect 324464 121320 324470 121332
rect 327534 121320 327540 121332
rect 327592 121320 327598 121372
rect 251542 121252 251548 121304
rect 251600 121292 251606 121304
rect 257430 121292 257436 121304
rect 251600 121264 257436 121292
rect 251600 121252 251606 121264
rect 257430 121252 257436 121264
rect 257488 121252 257494 121304
rect 343726 120708 343732 120760
rect 343784 120748 343790 120760
rect 383102 120748 383108 120760
rect 343784 120720 383108 120748
rect 343784 120708 343790 120720
rect 383102 120708 383108 120720
rect 383160 120708 383166 120760
rect 297634 120232 297640 120284
rect 297692 120272 297698 120284
rect 307570 120272 307576 120284
rect 297692 120244 307576 120272
rect 297692 120232 297698 120244
rect 307570 120232 307576 120244
rect 307628 120232 307634 120284
rect 187050 120164 187056 120216
rect 187108 120204 187114 120216
rect 213914 120204 213920 120216
rect 187108 120176 213920 120204
rect 187108 120164 187114 120176
rect 213914 120164 213920 120176
rect 213972 120164 213978 120216
rect 291838 120164 291844 120216
rect 291896 120204 291902 120216
rect 307662 120204 307668 120216
rect 291896 120176 307668 120204
rect 291896 120164 291902 120176
rect 307662 120164 307668 120176
rect 307720 120164 307726 120216
rect 182910 120096 182916 120148
rect 182968 120136 182974 120148
rect 214006 120136 214012 120148
rect 182968 120108 214012 120136
rect 182968 120096 182974 120108
rect 214006 120096 214012 120108
rect 214064 120096 214070 120148
rect 262950 120096 262956 120148
rect 263008 120136 263014 120148
rect 306742 120136 306748 120148
rect 263008 120108 306748 120136
rect 263008 120096 263014 120108
rect 306742 120096 306748 120108
rect 306800 120096 306806 120148
rect 252370 120028 252376 120080
rect 252428 120068 252434 120080
rect 289078 120068 289084 120080
rect 252428 120040 289084 120068
rect 252428 120028 252434 120040
rect 289078 120028 289084 120040
rect 289136 120028 289142 120080
rect 324314 120028 324320 120080
rect 324372 120068 324378 120080
rect 349338 120068 349344 120080
rect 324372 120040 349344 120068
rect 324372 120028 324378 120040
rect 349338 120028 349344 120040
rect 349396 120028 349402 120080
rect 370590 120028 370596 120080
rect 370648 120068 370654 120080
rect 386874 120068 386880 120080
rect 370648 120040 386880 120068
rect 370648 120028 370654 120040
rect 386874 120028 386880 120040
rect 386932 120028 386938 120080
rect 252462 119960 252468 120012
rect 252520 120000 252526 120012
rect 261570 120000 261576 120012
rect 252520 119972 261576 120000
rect 252520 119960 252526 119972
rect 261570 119960 261576 119972
rect 261628 119960 261634 120012
rect 340230 119960 340236 120012
rect 340288 120000 340294 120012
rect 363598 120000 363604 120012
rect 340288 119972 363604 120000
rect 340288 119960 340294 119972
rect 363598 119960 363604 119972
rect 363656 119960 363662 120012
rect 251726 119348 251732 119400
rect 251784 119388 251790 119400
rect 298738 119388 298744 119400
rect 251784 119360 298744 119388
rect 251784 119348 251790 119360
rect 298738 119348 298744 119360
rect 298796 119348 298802 119400
rect 349338 119348 349344 119400
rect 349396 119388 349402 119400
rect 378962 119388 378968 119400
rect 349396 119360 378968 119388
rect 349396 119348 349402 119360
rect 378962 119348 378968 119360
rect 379020 119348 379026 119400
rect 210602 118804 210608 118856
rect 210660 118844 210666 118856
rect 214098 118844 214104 118856
rect 210660 118816 214104 118844
rect 210660 118804 210666 118816
rect 214098 118804 214104 118816
rect 214156 118804 214162 118856
rect 302970 118804 302976 118856
rect 303028 118844 303034 118856
rect 307662 118844 307668 118856
rect 303028 118816 307668 118844
rect 303028 118804 303034 118816
rect 307662 118804 307668 118816
rect 307720 118804 307726 118856
rect 212166 118736 212172 118788
rect 212224 118776 212230 118788
rect 214006 118776 214012 118788
rect 212224 118748 214012 118776
rect 212224 118736 212230 118748
rect 214006 118736 214012 118748
rect 214064 118736 214070 118788
rect 296162 118736 296168 118788
rect 296220 118776 296226 118788
rect 307110 118776 307116 118788
rect 296220 118748 307116 118776
rect 296220 118736 296226 118748
rect 307110 118736 307116 118748
rect 307168 118736 307174 118788
rect 166442 118668 166448 118720
rect 166500 118708 166506 118720
rect 213914 118708 213920 118720
rect 166500 118680 213920 118708
rect 166500 118668 166506 118680
rect 213914 118668 213920 118680
rect 213972 118668 213978 118720
rect 287698 118668 287704 118720
rect 287756 118708 287762 118720
rect 306558 118708 306564 118720
rect 287756 118680 306564 118708
rect 287756 118668 287762 118680
rect 306558 118668 306564 118680
rect 306616 118668 306622 118720
rect 252370 118600 252376 118652
rect 252428 118640 252434 118652
rect 290642 118640 290648 118652
rect 252428 118612 290648 118640
rect 252428 118600 252434 118612
rect 290642 118600 290648 118612
rect 290700 118600 290706 118652
rect 324406 118600 324412 118652
rect 324464 118640 324470 118652
rect 340230 118640 340236 118652
rect 324464 118612 340236 118640
rect 324464 118600 324470 118612
rect 340230 118600 340236 118612
rect 340288 118600 340294 118652
rect 252462 118532 252468 118584
rect 252520 118572 252526 118584
rect 258810 118572 258816 118584
rect 252520 118544 258816 118572
rect 252520 118532 252526 118544
rect 258810 118532 258816 118544
rect 258868 118532 258874 118584
rect 324314 118532 324320 118584
rect 324372 118572 324378 118584
rect 330570 118572 330576 118584
rect 324372 118544 330576 118572
rect 324372 118532 324378 118544
rect 330570 118532 330576 118544
rect 330628 118532 330634 118584
rect 252094 117920 252100 117972
rect 252152 117960 252158 117972
rect 301590 117960 301596 117972
rect 252152 117932 301596 117960
rect 252152 117920 252158 117932
rect 301590 117920 301596 117932
rect 301648 117920 301654 117972
rect 324498 117920 324504 117972
rect 324556 117960 324562 117972
rect 354674 117960 354680 117972
rect 324556 117932 354680 117960
rect 324556 117920 324562 117932
rect 354674 117920 354680 117932
rect 354732 117920 354738 117972
rect 300118 117444 300124 117496
rect 300176 117484 300182 117496
rect 306558 117484 306564 117496
rect 300176 117456 306564 117484
rect 300176 117444 300182 117456
rect 306558 117444 306564 117456
rect 306616 117444 306622 117496
rect 203610 117376 203616 117428
rect 203668 117416 203674 117428
rect 213914 117416 213920 117428
rect 203668 117388 213920 117416
rect 203668 117376 203674 117388
rect 213914 117376 213920 117388
rect 213972 117376 213978 117428
rect 301774 117376 301780 117428
rect 301832 117416 301838 117428
rect 307662 117416 307668 117428
rect 301832 117388 307668 117416
rect 301832 117376 301838 117388
rect 307662 117376 307668 117388
rect 307720 117376 307726 117428
rect 195330 117308 195336 117360
rect 195388 117348 195394 117360
rect 214006 117348 214012 117360
rect 195388 117320 214012 117348
rect 195388 117308 195394 117320
rect 214006 117308 214012 117320
rect 214064 117308 214070 117360
rect 289262 117308 289268 117360
rect 289320 117348 289326 117360
rect 306926 117348 306932 117360
rect 289320 117320 306932 117348
rect 289320 117308 289326 117320
rect 306926 117308 306932 117320
rect 306984 117308 306990 117360
rect 252462 117240 252468 117292
rect 252520 117280 252526 117292
rect 287974 117280 287980 117292
rect 252520 117252 287980 117280
rect 252520 117240 252526 117252
rect 287974 117240 287980 117252
rect 288032 117240 288038 117292
rect 324314 117240 324320 117292
rect 324372 117280 324378 117292
rect 356054 117280 356060 117292
rect 324372 117252 356060 117280
rect 324372 117240 324378 117252
rect 356054 117240 356060 117252
rect 356112 117280 356118 117292
rect 357342 117280 357348 117292
rect 356112 117252 357348 117280
rect 356112 117240 356118 117252
rect 357342 117240 357348 117252
rect 357400 117240 357406 117292
rect 572622 117240 572628 117292
rect 572680 117280 572686 117292
rect 583202 117280 583208 117292
rect 572680 117252 583208 117280
rect 572680 117240 572686 117252
rect 583202 117240 583208 117252
rect 583260 117240 583266 117292
rect 251818 116560 251824 116612
rect 251876 116600 251882 116612
rect 264330 116600 264336 116612
rect 251876 116572 264336 116600
rect 251876 116560 251882 116572
rect 264330 116560 264336 116572
rect 264388 116560 264394 116612
rect 252002 116356 252008 116408
rect 252060 116396 252066 116408
rect 257614 116396 257620 116408
rect 252060 116368 257620 116396
rect 252060 116356 252066 116368
rect 257614 116356 257620 116368
rect 257672 116356 257678 116408
rect 298738 116084 298744 116136
rect 298796 116124 298802 116136
rect 307570 116124 307576 116136
rect 298796 116096 307576 116124
rect 298796 116084 298802 116096
rect 307570 116084 307576 116096
rect 307628 116084 307634 116136
rect 282270 116016 282276 116068
rect 282328 116056 282334 116068
rect 307662 116056 307668 116068
rect 282328 116028 307668 116056
rect 282328 116016 282334 116028
rect 307662 116016 307668 116028
rect 307720 116016 307726 116068
rect 193950 115948 193956 116000
rect 194008 115988 194014 116000
rect 213914 115988 213920 116000
rect 194008 115960 213920 115988
rect 194008 115948 194014 115960
rect 213914 115948 213920 115960
rect 213972 115948 213978 116000
rect 261570 115948 261576 116000
rect 261628 115988 261634 116000
rect 307478 115988 307484 116000
rect 261628 115960 307484 115988
rect 261628 115948 261634 115960
rect 307478 115948 307484 115960
rect 307536 115948 307542 116000
rect 252002 115880 252008 115932
rect 252060 115920 252066 115932
rect 300210 115920 300216 115932
rect 252060 115892 300216 115920
rect 252060 115880 252066 115892
rect 300210 115880 300216 115892
rect 300268 115880 300274 115932
rect 324406 115880 324412 115932
rect 324464 115920 324470 115932
rect 345106 115920 345112 115932
rect 324464 115892 345112 115920
rect 324464 115880 324470 115892
rect 345106 115880 345112 115892
rect 345164 115920 345170 115932
rect 346302 115920 346308 115932
rect 345164 115892 346308 115920
rect 345164 115880 345170 115892
rect 346302 115880 346308 115892
rect 346360 115880 346366 115932
rect 252278 115812 252284 115864
rect 252336 115852 252342 115864
rect 287882 115852 287888 115864
rect 252336 115824 287888 115852
rect 252336 115812 252342 115824
rect 287882 115812 287888 115824
rect 287940 115812 287946 115864
rect 324774 115200 324780 115252
rect 324832 115240 324838 115252
rect 340138 115240 340144 115252
rect 324832 115212 340144 115240
rect 324832 115200 324838 115212
rect 340138 115200 340144 115212
rect 340196 115200 340202 115252
rect 324314 115064 324320 115116
rect 324372 115104 324378 115116
rect 327718 115104 327724 115116
rect 324372 115076 327724 115104
rect 324372 115064 324378 115076
rect 327718 115064 327724 115076
rect 327776 115064 327782 115116
rect 210418 114588 210424 114640
rect 210476 114628 210482 114640
rect 214006 114628 214012 114640
rect 210476 114600 214012 114628
rect 210476 114588 210482 114600
rect 214006 114588 214012 114600
rect 214064 114588 214070 114640
rect 293310 114588 293316 114640
rect 293368 114628 293374 114640
rect 307478 114628 307484 114640
rect 293368 114600 307484 114628
rect 293368 114588 293374 114600
rect 307478 114588 307484 114600
rect 307536 114588 307542 114640
rect 177390 114520 177396 114572
rect 177448 114560 177454 114572
rect 213914 114560 213920 114572
rect 177448 114532 213920 114560
rect 177448 114520 177454 114532
rect 213914 114520 213920 114532
rect 213972 114520 213978 114572
rect 249150 114520 249156 114572
rect 249208 114560 249214 114572
rect 307110 114560 307116 114572
rect 249208 114532 307116 114560
rect 249208 114520 249214 114532
rect 307110 114520 307116 114532
rect 307168 114520 307174 114572
rect 352558 114520 352564 114572
rect 352616 114560 352622 114572
rect 354674 114560 354680 114572
rect 352616 114532 354680 114560
rect 352616 114520 352622 114532
rect 354674 114520 354680 114532
rect 354732 114560 354738 114572
rect 386874 114560 386880 114572
rect 354732 114532 386880 114560
rect 354732 114520 354738 114532
rect 386874 114520 386880 114532
rect 386932 114520 386938 114572
rect 251542 114452 251548 114504
rect 251600 114492 251606 114504
rect 271414 114492 271420 114504
rect 251600 114464 271420 114492
rect 251600 114452 251606 114464
rect 271414 114452 271420 114464
rect 271472 114452 271478 114504
rect 324406 114452 324412 114504
rect 324464 114492 324470 114504
rect 373994 114492 374000 114504
rect 324464 114464 374000 114492
rect 324464 114452 324470 114464
rect 373994 114452 374000 114464
rect 374052 114452 374058 114504
rect 252462 114384 252468 114436
rect 252520 114424 252526 114436
rect 260282 114424 260288 114436
rect 252520 114396 260288 114424
rect 252520 114384 252526 114396
rect 260282 114384 260288 114396
rect 260340 114384 260346 114436
rect 324314 114384 324320 114436
rect 324372 114424 324378 114436
rect 336734 114424 336740 114436
rect 324372 114396 336740 114424
rect 324372 114384 324378 114396
rect 336734 114384 336740 114396
rect 336792 114424 336798 114436
rect 338022 114424 338028 114436
rect 336792 114396 338028 114424
rect 336792 114384 336798 114396
rect 338022 114384 338028 114396
rect 338080 114384 338086 114436
rect 252186 114316 252192 114368
rect 252244 114356 252250 114368
rect 254854 114356 254860 114368
rect 252244 114328 254860 114356
rect 252244 114316 252250 114328
rect 254854 114316 254860 114328
rect 254912 114316 254918 114368
rect 260098 113772 260104 113824
rect 260156 113812 260162 113824
rect 284294 113812 284300 113824
rect 260156 113784 284300 113812
rect 260156 113772 260162 113784
rect 284294 113772 284300 113784
rect 284352 113772 284358 113824
rect 338022 113772 338028 113824
rect 338080 113812 338086 113824
rect 388530 113812 388536 113824
rect 338080 113784 388536 113812
rect 338080 113772 338086 113784
rect 388530 113772 388536 113784
rect 388588 113772 388594 113824
rect 289078 113296 289084 113348
rect 289136 113336 289142 113348
rect 307662 113336 307668 113348
rect 289136 113308 307668 113336
rect 289136 113296 289142 113308
rect 307662 113296 307668 113308
rect 307720 113296 307726 113348
rect 184382 113228 184388 113280
rect 184440 113268 184446 113280
rect 213914 113268 213920 113280
rect 184440 113240 213920 113268
rect 184440 113228 184446 113240
rect 213914 113228 213920 113240
rect 213972 113228 213978 113280
rect 254578 113228 254584 113280
rect 254636 113268 254642 113280
rect 254636 113240 258074 113268
rect 254636 113228 254642 113240
rect 171962 113160 171968 113212
rect 172020 113200 172026 113212
rect 214006 113200 214012 113212
rect 172020 113172 214012 113200
rect 172020 113160 172026 113172
rect 214006 113160 214012 113172
rect 214064 113160 214070 113212
rect 258046 113200 258074 113240
rect 272518 113228 272524 113280
rect 272576 113268 272582 113280
rect 307570 113268 307576 113280
rect 272576 113240 307576 113268
rect 272576 113228 272582 113240
rect 307570 113228 307576 113240
rect 307628 113228 307634 113280
rect 306558 113200 306564 113212
rect 258046 113172 306564 113200
rect 306558 113160 306564 113172
rect 306616 113160 306622 113212
rect 251542 113092 251548 113144
rect 251600 113132 251606 113144
rect 296254 113132 296260 113144
rect 251600 113104 296260 113132
rect 251600 113092 251606 113104
rect 296254 113092 296260 113104
rect 296312 113092 296318 113144
rect 324314 113092 324320 113144
rect 324372 113132 324378 113144
rect 338114 113132 338120 113144
rect 324372 113104 338120 113132
rect 324372 113092 324378 113104
rect 338114 113092 338120 113104
rect 338172 113092 338178 113144
rect 252462 113024 252468 113076
rect 252520 113064 252526 113076
rect 275370 113064 275376 113076
rect 252520 113036 275376 113064
rect 252520 113024 252526 113036
rect 275370 113024 275376 113036
rect 275428 113024 275434 113076
rect 338114 112480 338120 112532
rect 338172 112520 338178 112532
rect 376110 112520 376116 112532
rect 338172 112492 376116 112520
rect 338172 112480 338178 112492
rect 376110 112480 376116 112492
rect 376168 112480 376174 112532
rect 325050 112412 325056 112464
rect 325108 112452 325114 112464
rect 387150 112452 387156 112464
rect 325108 112424 387156 112452
rect 325108 112412 325114 112424
rect 387150 112412 387156 112424
rect 387208 112412 387214 112464
rect 252370 112208 252376 112260
rect 252428 112248 252434 112260
rect 258718 112248 258724 112260
rect 252428 112220 258724 112248
rect 252428 112208 252434 112220
rect 258718 112208 258724 112220
rect 258776 112208 258782 112260
rect 199378 111868 199384 111920
rect 199436 111908 199442 111920
rect 213914 111908 213920 111920
rect 199436 111880 213920 111908
rect 199436 111868 199442 111880
rect 213914 111868 213920 111880
rect 213972 111868 213978 111920
rect 299014 111868 299020 111920
rect 299072 111908 299078 111920
rect 307570 111908 307576 111920
rect 299072 111880 307576 111908
rect 299072 111868 299078 111880
rect 307570 111868 307576 111880
rect 307628 111868 307634 111920
rect 192662 111800 192668 111852
rect 192720 111840 192726 111852
rect 214006 111840 214012 111852
rect 192720 111812 214012 111840
rect 192720 111800 192726 111812
rect 214006 111800 214012 111812
rect 214064 111800 214070 111852
rect 295978 111800 295984 111852
rect 296036 111840 296042 111852
rect 307662 111840 307668 111852
rect 296036 111812 307668 111840
rect 296036 111800 296042 111812
rect 307662 111800 307668 111812
rect 307720 111800 307726 111852
rect 570598 111800 570604 111852
rect 570656 111840 570662 111852
rect 579890 111840 579896 111852
rect 570656 111812 579896 111840
rect 570656 111800 570662 111812
rect 579890 111800 579896 111812
rect 579948 111800 579954 111852
rect 252462 111732 252468 111784
rect 252520 111772 252526 111784
rect 273990 111772 273996 111784
rect 252520 111744 273996 111772
rect 252520 111732 252526 111744
rect 273990 111732 273996 111744
rect 274048 111732 274054 111784
rect 324314 111732 324320 111784
rect 324372 111772 324378 111784
rect 347774 111772 347780 111784
rect 324372 111744 347780 111772
rect 324372 111732 324378 111744
rect 347774 111732 347780 111744
rect 347832 111732 347838 111784
rect 252370 111664 252376 111716
rect 252428 111704 252434 111716
rect 257338 111704 257344 111716
rect 252428 111676 257344 111704
rect 252428 111664 252434 111676
rect 257338 111664 257344 111676
rect 257396 111664 257402 111716
rect 347774 111052 347780 111104
rect 347832 111092 347838 111104
rect 388714 111092 388720 111104
rect 347832 111064 388720 111092
rect 347832 111052 347838 111064
rect 388714 111052 388720 111064
rect 388772 111052 388778 111104
rect 324406 110712 324412 110764
rect 324464 110752 324470 110764
rect 327074 110752 327080 110764
rect 324464 110724 327080 110752
rect 324464 110712 324470 110724
rect 327074 110712 327080 110724
rect 327132 110712 327138 110764
rect 300210 110576 300216 110628
rect 300268 110616 300274 110628
rect 307662 110616 307668 110628
rect 300268 110588 307668 110616
rect 300268 110576 300274 110588
rect 307662 110576 307668 110588
rect 307720 110576 307726 110628
rect 189902 110508 189908 110560
rect 189960 110548 189966 110560
rect 213914 110548 213920 110560
rect 189960 110520 213920 110548
rect 189960 110508 189966 110520
rect 213914 110508 213920 110520
rect 213972 110508 213978 110560
rect 274082 110508 274088 110560
rect 274140 110548 274146 110560
rect 307478 110548 307484 110560
rect 274140 110520 307484 110548
rect 274140 110508 274146 110520
rect 307478 110508 307484 110520
rect 307536 110508 307542 110560
rect 169202 110440 169208 110492
rect 169260 110480 169266 110492
rect 214006 110480 214012 110492
rect 169260 110452 214012 110480
rect 169260 110440 169266 110452
rect 214006 110440 214012 110452
rect 214064 110440 214070 110492
rect 258718 110440 258724 110492
rect 258776 110480 258782 110492
rect 307570 110480 307576 110492
rect 258776 110452 307576 110480
rect 258776 110440 258782 110452
rect 307570 110440 307576 110452
rect 307628 110440 307634 110492
rect 252370 110372 252376 110424
rect 252428 110412 252434 110424
rect 304350 110412 304356 110424
rect 252428 110384 304356 110412
rect 252428 110372 252434 110384
rect 304350 110372 304356 110384
rect 304408 110372 304414 110424
rect 324314 110372 324320 110424
rect 324372 110412 324378 110424
rect 329926 110412 329932 110424
rect 324372 110384 329932 110412
rect 324372 110372 324378 110384
rect 329926 110372 329932 110384
rect 329984 110372 329990 110424
rect 252462 110304 252468 110356
rect 252520 110344 252526 110356
rect 289354 110344 289360 110356
rect 252520 110316 289360 110344
rect 252520 110304 252526 110316
rect 289354 110304 289360 110316
rect 289412 110304 289418 110356
rect 252094 109964 252100 110016
rect 252152 110004 252158 110016
rect 256050 110004 256056 110016
rect 252152 109976 256056 110004
rect 252152 109964 252158 109976
rect 256050 109964 256056 109976
rect 256108 109964 256114 110016
rect 301590 109148 301596 109200
rect 301648 109188 301654 109200
rect 307662 109188 307668 109200
rect 301648 109160 307668 109188
rect 301648 109148 301654 109160
rect 307662 109148 307668 109160
rect 307720 109148 307726 109200
rect 209038 109080 209044 109132
rect 209096 109120 209102 109132
rect 214006 109120 214012 109132
rect 209096 109092 214012 109120
rect 209096 109080 209102 109092
rect 214006 109080 214012 109092
rect 214064 109080 214070 109132
rect 304534 109080 304540 109132
rect 304592 109120 304598 109132
rect 306926 109120 306932 109132
rect 304592 109092 306932 109120
rect 304592 109080 304598 109092
rect 306926 109080 306932 109092
rect 306984 109080 306990 109132
rect 167914 109012 167920 109064
rect 167972 109052 167978 109064
rect 213914 109052 213920 109064
rect 167972 109024 213920 109052
rect 167972 109012 167978 109024
rect 213914 109012 213920 109024
rect 213972 109012 213978 109064
rect 273990 109012 273996 109064
rect 274048 109052 274054 109064
rect 307570 109052 307576 109064
rect 274048 109024 307576 109052
rect 274048 109012 274054 109024
rect 307570 109012 307576 109024
rect 307628 109012 307634 109064
rect 168098 108944 168104 108996
rect 168156 108984 168162 108996
rect 177482 108984 177488 108996
rect 168156 108956 177488 108984
rect 168156 108944 168162 108956
rect 177482 108944 177488 108956
rect 177540 108944 177546 108996
rect 252462 108944 252468 108996
rect 252520 108984 252526 108996
rect 283926 108984 283932 108996
rect 252520 108956 283932 108984
rect 252520 108944 252526 108956
rect 283926 108944 283932 108956
rect 283984 108944 283990 108996
rect 353938 108944 353944 108996
rect 353996 108984 354002 108996
rect 386598 108984 386604 108996
rect 353996 108956 386604 108984
rect 353996 108944 354002 108956
rect 386598 108944 386604 108956
rect 386656 108944 386662 108996
rect 252370 108876 252376 108928
rect 252428 108916 252434 108928
rect 260190 108916 260196 108928
rect 252428 108888 260196 108916
rect 252428 108876 252434 108888
rect 260190 108876 260196 108888
rect 260248 108876 260254 108928
rect 252094 108672 252100 108724
rect 252152 108712 252158 108724
rect 256142 108712 256148 108724
rect 252152 108684 256148 108712
rect 252152 108672 252158 108684
rect 256142 108672 256148 108684
rect 256200 108672 256206 108724
rect 214742 108400 214748 108452
rect 214800 108400 214806 108452
rect 214650 108196 214656 108248
rect 214708 108236 214714 108248
rect 214760 108236 214788 108400
rect 324314 108332 324320 108384
rect 324372 108372 324378 108384
rect 325786 108372 325792 108384
rect 324372 108344 325792 108372
rect 324372 108332 324378 108344
rect 325786 108332 325792 108344
rect 325844 108372 325850 108384
rect 329190 108372 329196 108384
rect 325844 108344 329196 108372
rect 325844 108332 325850 108344
rect 329190 108332 329196 108344
rect 329248 108332 329254 108384
rect 324406 108264 324412 108316
rect 324464 108304 324470 108316
rect 351270 108304 351276 108316
rect 324464 108276 351276 108304
rect 324464 108264 324470 108276
rect 351270 108264 351276 108276
rect 351328 108264 351334 108316
rect 214708 108208 214788 108236
rect 214708 108196 214714 108208
rect 258810 107856 258816 107908
rect 258868 107896 258874 107908
rect 307662 107896 307668 107908
rect 258868 107868 307668 107896
rect 258868 107856 258874 107868
rect 307662 107856 307668 107868
rect 307720 107856 307726 107908
rect 300302 107788 300308 107840
rect 300360 107828 300366 107840
rect 307570 107828 307576 107840
rect 300360 107800 307576 107828
rect 300360 107788 300366 107800
rect 307570 107788 307576 107800
rect 307628 107788 307634 107840
rect 207842 107720 207848 107772
rect 207900 107760 207906 107772
rect 213914 107760 213920 107772
rect 207900 107732 213920 107760
rect 207900 107720 207906 107732
rect 213914 107720 213920 107732
rect 213972 107720 213978 107772
rect 264238 107720 264244 107772
rect 264296 107760 264302 107772
rect 307386 107760 307392 107772
rect 264296 107732 307392 107760
rect 264296 107720 264302 107732
rect 307386 107720 307392 107732
rect 307444 107720 307450 107772
rect 188522 107652 188528 107704
rect 188580 107692 188586 107704
rect 214006 107692 214012 107704
rect 188580 107664 214012 107692
rect 188580 107652 188586 107664
rect 214006 107652 214012 107664
rect 214064 107652 214070 107704
rect 304442 107652 304448 107704
rect 304500 107692 304506 107704
rect 307478 107692 307484 107704
rect 304500 107664 307484 107692
rect 304500 107652 304506 107664
rect 307478 107652 307484 107664
rect 307536 107652 307542 107704
rect 252462 107584 252468 107636
rect 252520 107624 252526 107636
rect 272610 107624 272616 107636
rect 252520 107596 272616 107624
rect 252520 107584 252526 107596
rect 272610 107584 272616 107596
rect 272668 107584 272674 107636
rect 252370 107516 252376 107568
rect 252428 107556 252434 107568
rect 269850 107556 269856 107568
rect 252428 107528 269856 107556
rect 252428 107516 252434 107528
rect 269850 107516 269856 107528
rect 269908 107516 269914 107568
rect 251542 107040 251548 107092
rect 251600 107080 251606 107092
rect 254670 107080 254676 107092
rect 251600 107052 254676 107080
rect 251600 107040 251606 107052
rect 254670 107040 254676 107052
rect 254728 107040 254734 107092
rect 252462 106904 252468 106956
rect 252520 106944 252526 106956
rect 263042 106944 263048 106956
rect 252520 106916 263048 106944
rect 252520 106904 252526 106916
rect 263042 106904 263048 106916
rect 263100 106904 263106 106956
rect 575382 106904 575388 106956
rect 575440 106944 575446 106956
rect 580350 106944 580356 106956
rect 575440 106916 580356 106944
rect 575440 106904 575446 106916
rect 580350 106904 580356 106916
rect 580408 106904 580414 106956
rect 256050 106428 256056 106480
rect 256108 106468 256114 106480
rect 307662 106468 307668 106480
rect 256108 106440 307668 106468
rect 256108 106428 256114 106440
rect 307662 106428 307668 106440
rect 307720 106428 307726 106480
rect 185670 106360 185676 106412
rect 185728 106400 185734 106412
rect 213914 106400 213920 106412
rect 185728 106372 213920 106400
rect 185728 106360 185734 106372
rect 213914 106360 213920 106372
rect 213972 106360 213978 106412
rect 271414 106360 271420 106412
rect 271472 106400 271478 106412
rect 307570 106400 307576 106412
rect 271472 106372 307576 106400
rect 271472 106360 271478 106372
rect 307570 106360 307576 106372
rect 307628 106360 307634 106412
rect 170674 106292 170680 106344
rect 170732 106332 170738 106344
rect 214006 106332 214012 106344
rect 170732 106304 214012 106332
rect 170732 106292 170738 106304
rect 214006 106292 214012 106304
rect 214064 106292 214070 106344
rect 321554 106292 321560 106344
rect 321612 106332 321618 106344
rect 387242 106332 387248 106344
rect 321612 106304 387248 106332
rect 321612 106292 321618 106304
rect 387242 106292 387248 106304
rect 387300 106292 387306 106344
rect 571242 106292 571248 106344
rect 571300 106332 571306 106344
rect 574830 106332 574836 106344
rect 571300 106304 574836 106332
rect 571300 106292 571306 106304
rect 574830 106292 574836 106304
rect 574888 106292 574894 106344
rect 252094 106224 252100 106276
rect 252152 106264 252158 106276
rect 283834 106264 283840 106276
rect 252152 106236 283840 106264
rect 252152 106224 252158 106236
rect 283834 106224 283840 106236
rect 283892 106224 283898 106276
rect 324314 106224 324320 106276
rect 324372 106264 324378 106276
rect 354674 106264 354680 106276
rect 324372 106236 354680 106264
rect 324372 106224 324378 106236
rect 354674 106224 354680 106236
rect 354732 106224 354738 106276
rect 251634 106156 251640 106208
rect 251692 106196 251698 106208
rect 254762 106196 254768 106208
rect 251692 106168 254768 106196
rect 251692 106156 251698 106168
rect 254762 106156 254768 106168
rect 254820 106156 254826 106208
rect 252002 105544 252008 105596
rect 252060 105584 252066 105596
rect 301498 105584 301504 105596
rect 252060 105556 301504 105584
rect 252060 105544 252066 105556
rect 301498 105544 301504 105556
rect 301556 105544 301562 105596
rect 337378 105544 337384 105596
rect 337436 105584 337442 105596
rect 389726 105584 389732 105596
rect 337436 105556 389732 105584
rect 337436 105544 337442 105556
rect 389726 105544 389732 105556
rect 389784 105544 389790 105596
rect 205082 105000 205088 105052
rect 205140 105040 205146 105052
rect 213914 105040 213920 105052
rect 205140 105012 213920 105040
rect 205140 105000 205146 105012
rect 213914 105000 213920 105012
rect 213972 105000 213978 105052
rect 203702 104932 203708 104984
rect 203760 104972 203766 104984
rect 214006 104972 214012 104984
rect 203760 104944 214012 104972
rect 203760 104932 203766 104944
rect 214006 104932 214012 104944
rect 214064 104932 214070 104984
rect 301682 104932 301688 104984
rect 301740 104972 301746 104984
rect 307570 104972 307576 104984
rect 301740 104944 307576 104972
rect 301740 104932 301746 104944
rect 307570 104932 307576 104944
rect 307628 104932 307634 104984
rect 191190 104864 191196 104916
rect 191248 104904 191254 104916
rect 214098 104904 214104 104916
rect 191248 104876 214104 104904
rect 191248 104864 191254 104876
rect 214098 104864 214104 104876
rect 214156 104864 214162 104916
rect 283650 104864 283656 104916
rect 283708 104904 283714 104916
rect 307662 104904 307668 104916
rect 283708 104876 307668 104904
rect 283708 104864 283714 104876
rect 307662 104864 307668 104876
rect 307720 104864 307726 104916
rect 252094 104796 252100 104848
rect 252152 104836 252158 104848
rect 305730 104836 305736 104848
rect 252152 104808 305736 104836
rect 252152 104796 252158 104808
rect 305730 104796 305736 104808
rect 305788 104796 305794 104848
rect 252278 104388 252284 104440
rect 252336 104428 252342 104440
rect 255958 104428 255964 104440
rect 252336 104400 255964 104428
rect 252336 104388 252342 104400
rect 255958 104388 255964 104400
rect 256016 104388 256022 104440
rect 285122 103640 285128 103692
rect 285180 103680 285186 103692
rect 307478 103680 307484 103692
rect 285180 103652 307484 103680
rect 285180 103640 285186 103652
rect 307478 103640 307484 103652
rect 307536 103640 307542 103692
rect 198274 103572 198280 103624
rect 198332 103612 198338 103624
rect 213914 103612 213920 103624
rect 198332 103584 213920 103612
rect 198332 103572 198338 103584
rect 213914 103572 213920 103584
rect 213972 103572 213978 103624
rect 296254 103572 296260 103624
rect 296312 103612 296318 103624
rect 307662 103612 307668 103624
rect 296312 103584 307668 103612
rect 296312 103572 296318 103584
rect 307662 103572 307668 103584
rect 307720 103572 307726 103624
rect 194042 103504 194048 103556
rect 194100 103544 194106 103556
rect 214006 103544 214012 103556
rect 194100 103516 214012 103544
rect 194100 103504 194106 103516
rect 214006 103504 214012 103516
rect 214064 103504 214070 103556
rect 322934 103504 322940 103556
rect 322992 103544 322998 103556
rect 385954 103544 385960 103556
rect 322992 103516 385960 103544
rect 322992 103504 322998 103516
rect 385954 103504 385960 103516
rect 386012 103504 386018 103556
rect 252462 103436 252468 103488
rect 252520 103476 252526 103488
rect 264514 103476 264520 103488
rect 252520 103448 264520 103476
rect 252520 103436 252526 103448
rect 264514 103436 264520 103448
rect 264572 103436 264578 103488
rect 324406 103436 324412 103488
rect 324464 103476 324470 103488
rect 346394 103476 346400 103488
rect 324464 103448 346400 103476
rect 324464 103436 324470 103448
rect 346394 103436 346400 103448
rect 346452 103436 346458 103488
rect 252370 102756 252376 102808
rect 252428 102796 252434 102808
rect 293402 102796 293408 102808
rect 252428 102768 293408 102796
rect 252428 102756 252434 102768
rect 293402 102756 293408 102768
rect 293460 102756 293466 102808
rect 304350 102280 304356 102332
rect 304408 102320 304414 102332
rect 306742 102320 306748 102332
rect 304408 102292 306748 102320
rect 304408 102280 304414 102292
rect 306742 102280 306748 102292
rect 306800 102280 306806 102332
rect 200758 102212 200764 102264
rect 200816 102252 200822 102264
rect 214006 102252 214012 102264
rect 200816 102224 214012 102252
rect 200816 102212 200822 102224
rect 214006 102212 214012 102224
rect 214064 102212 214070 102264
rect 292022 102212 292028 102264
rect 292080 102252 292086 102264
rect 307478 102252 307484 102264
rect 292080 102224 307484 102252
rect 292080 102212 292086 102224
rect 307478 102212 307484 102224
rect 307536 102212 307542 102264
rect 198182 102144 198188 102196
rect 198240 102184 198246 102196
rect 213914 102184 213920 102196
rect 198240 102156 213920 102184
rect 198240 102144 198246 102156
rect 213914 102144 213920 102156
rect 213972 102144 213978 102196
rect 269850 102144 269856 102196
rect 269908 102184 269914 102196
rect 307662 102184 307668 102196
rect 269908 102156 307668 102184
rect 269908 102144 269914 102156
rect 307662 102144 307668 102156
rect 307720 102144 307726 102196
rect 572622 102144 572628 102196
rect 572680 102184 572686 102196
rect 574186 102184 574192 102196
rect 572680 102156 574192 102184
rect 572680 102144 572686 102156
rect 574186 102144 574192 102156
rect 574244 102144 574250 102196
rect 252094 102076 252100 102128
rect 252152 102116 252158 102128
rect 278314 102116 278320 102128
rect 252152 102088 278320 102116
rect 252152 102076 252158 102088
rect 278314 102076 278320 102088
rect 278372 102076 278378 102128
rect 251818 102008 251824 102060
rect 251876 102048 251882 102060
rect 267090 102048 267096 102060
rect 251876 102020 267096 102048
rect 251876 102008 251882 102020
rect 267090 102008 267096 102020
rect 267148 102008 267154 102060
rect 292666 101396 292672 101448
rect 292724 101436 292730 101448
rect 302234 101436 302240 101448
rect 292724 101408 302240 101436
rect 292724 101396 292730 101408
rect 302234 101396 302240 101408
rect 302292 101396 302298 101448
rect 324590 101396 324596 101448
rect 324648 101436 324654 101448
rect 337470 101436 337476 101448
rect 324648 101408 337476 101436
rect 324648 101396 324654 101408
rect 337470 101396 337476 101408
rect 337528 101396 337534 101448
rect 303062 100920 303068 100972
rect 303120 100960 303126 100972
rect 306742 100960 306748 100972
rect 303120 100932 306748 100960
rect 303120 100920 303126 100932
rect 306742 100920 306748 100932
rect 306800 100920 306806 100972
rect 287882 100852 287888 100904
rect 287940 100892 287946 100904
rect 307478 100892 307484 100904
rect 287940 100864 307484 100892
rect 287940 100852 287946 100864
rect 307478 100852 307484 100864
rect 307536 100852 307542 100904
rect 275370 100784 275376 100836
rect 275428 100824 275434 100836
rect 307662 100824 307668 100836
rect 275428 100796 307668 100824
rect 275428 100784 275434 100796
rect 307662 100784 307668 100796
rect 307720 100784 307726 100836
rect 204990 100716 204996 100768
rect 205048 100756 205054 100768
rect 213914 100756 213920 100768
rect 205048 100728 213920 100756
rect 205048 100716 205054 100728
rect 213914 100716 213920 100728
rect 213972 100716 213978 100768
rect 271230 100716 271236 100768
rect 271288 100756 271294 100768
rect 307570 100756 307576 100768
rect 271288 100728 307576 100756
rect 271288 100716 271294 100728
rect 307570 100716 307576 100728
rect 307628 100716 307634 100768
rect 251910 100648 251916 100700
rect 251968 100688 251974 100700
rect 297726 100688 297732 100700
rect 251968 100660 297732 100688
rect 251968 100648 251974 100660
rect 297726 100648 297732 100660
rect 297784 100648 297790 100700
rect 252094 100580 252100 100632
rect 252152 100620 252158 100632
rect 261754 100620 261760 100632
rect 252152 100592 261760 100620
rect 252152 100580 252158 100592
rect 261754 100580 261760 100592
rect 261812 100580 261818 100632
rect 169294 100036 169300 100088
rect 169352 100076 169358 100088
rect 214650 100076 214656 100088
rect 169352 100048 214656 100076
rect 169352 100036 169358 100048
rect 214650 100036 214656 100048
rect 214708 100036 214714 100088
rect 166534 99968 166540 100020
rect 166592 100008 166598 100020
rect 214374 100008 214380 100020
rect 166592 99980 214380 100008
rect 166592 99968 166598 99980
rect 214374 99968 214380 99980
rect 214432 99968 214438 100020
rect 252278 99968 252284 100020
rect 252336 100008 252342 100020
rect 306006 100008 306012 100020
rect 252336 99980 306012 100008
rect 252336 99968 252342 99980
rect 306006 99968 306012 99980
rect 306064 99968 306070 100020
rect 297542 99356 297548 99408
rect 297600 99396 297606 99408
rect 307478 99396 307484 99408
rect 297600 99368 307484 99396
rect 297600 99356 297606 99368
rect 307478 99356 307484 99368
rect 307536 99356 307542 99408
rect 172422 99288 172428 99340
rect 172480 99328 172486 99340
rect 217962 99328 217968 99340
rect 172480 99300 217968 99328
rect 172480 99288 172486 99300
rect 217962 99288 217968 99300
rect 218020 99288 218026 99340
rect 324314 99288 324320 99340
rect 324372 99328 324378 99340
rect 368474 99328 368480 99340
rect 324372 99300 368480 99328
rect 324372 99288 324378 99300
rect 368474 99288 368480 99300
rect 368532 99288 368538 99340
rect 381630 99288 381636 99340
rect 381688 99328 381694 99340
rect 386874 99328 386880 99340
rect 381688 99300 386880 99328
rect 381688 99288 381694 99300
rect 386874 99288 386880 99300
rect 386932 99288 386938 99340
rect 252370 99220 252376 99272
rect 252428 99260 252434 99272
rect 299106 99260 299112 99272
rect 252428 99232 299112 99260
rect 252428 99220 252434 99232
rect 299106 99220 299112 99232
rect 299164 99220 299170 99272
rect 324406 99220 324412 99272
rect 324464 99260 324470 99272
rect 345014 99260 345020 99272
rect 324464 99232 345020 99260
rect 324464 99220 324470 99232
rect 345014 99220 345020 99232
rect 345072 99220 345078 99272
rect 251174 98948 251180 99000
rect 251232 98988 251238 99000
rect 253198 98988 253204 99000
rect 251232 98960 253204 98988
rect 251232 98948 251238 98960
rect 253198 98948 253204 98960
rect 253256 98948 253262 99000
rect 191098 98676 191104 98728
rect 191156 98716 191162 98728
rect 217318 98716 217324 98728
rect 191156 98688 217324 98716
rect 191156 98676 191162 98688
rect 217318 98676 217324 98688
rect 217376 98676 217382 98728
rect 188338 98608 188344 98660
rect 188396 98648 188402 98660
rect 217410 98648 217416 98660
rect 188396 98620 217416 98648
rect 188396 98608 188402 98620
rect 217410 98608 217416 98620
rect 217468 98608 217474 98660
rect 251910 98608 251916 98660
rect 251968 98648 251974 98660
rect 282362 98648 282368 98660
rect 251968 98620 282368 98648
rect 251968 98608 251974 98620
rect 282362 98608 282368 98620
rect 282420 98608 282426 98660
rect 301498 98132 301504 98184
rect 301556 98172 301562 98184
rect 306558 98172 306564 98184
rect 301556 98144 306564 98172
rect 301556 98132 301562 98144
rect 306558 98132 306564 98144
rect 306616 98132 306622 98184
rect 298830 98064 298836 98116
rect 298888 98104 298894 98116
rect 307570 98104 307576 98116
rect 298888 98076 307576 98104
rect 298888 98064 298894 98076
rect 307570 98064 307576 98076
rect 307628 98064 307634 98116
rect 167822 97996 167828 98048
rect 167880 98036 167886 98048
rect 213914 98036 213920 98048
rect 167880 98008 213920 98036
rect 167880 97996 167886 98008
rect 213914 97996 213920 98008
rect 213972 97996 213978 98048
rect 255958 97996 255964 98048
rect 256016 98036 256022 98048
rect 307662 98036 307668 98048
rect 256016 98008 307668 98036
rect 256016 97996 256022 98008
rect 307662 97996 307668 98008
rect 307720 97996 307726 98048
rect 389634 96772 389640 96824
rect 389692 96812 389698 96824
rect 389818 96812 389824 96824
rect 389692 96784 389824 96812
rect 389692 96772 389698 96784
rect 389818 96772 389824 96784
rect 389876 96772 389882 96824
rect 275278 96704 275284 96756
rect 275336 96744 275342 96756
rect 307662 96744 307668 96756
rect 275336 96716 307668 96744
rect 275336 96704 275342 96716
rect 307662 96704 307668 96716
rect 307720 96704 307726 96756
rect 207934 96636 207940 96688
rect 207992 96676 207998 96688
rect 213914 96676 213920 96688
rect 207992 96648 213920 96676
rect 207992 96636 207998 96648
rect 213914 96636 213920 96648
rect 213972 96636 213978 96688
rect 253290 96636 253296 96688
rect 253348 96676 253354 96688
rect 307478 96676 307484 96688
rect 253348 96648 307484 96676
rect 253348 96636 253354 96648
rect 307478 96636 307484 96648
rect 307536 96636 307542 96688
rect 198090 96568 198096 96620
rect 198148 96608 198154 96620
rect 321738 96608 321744 96620
rect 198148 96580 321744 96608
rect 198148 96568 198154 96580
rect 321738 96568 321744 96580
rect 321796 96568 321802 96620
rect 324314 96568 324320 96620
rect 324372 96608 324378 96620
rect 342346 96608 342352 96620
rect 324372 96580 342352 96608
rect 324372 96568 324378 96580
rect 342346 96568 342352 96580
rect 342404 96568 342410 96620
rect 378870 96568 378876 96620
rect 378928 96608 378934 96620
rect 575566 96608 575572 96620
rect 378928 96580 575572 96608
rect 378928 96568 378934 96580
rect 575566 96568 575572 96580
rect 575624 96568 575630 96620
rect 383010 96500 383016 96552
rect 383068 96540 383074 96552
rect 568574 96540 568580 96552
rect 383068 96512 568580 96540
rect 383068 96500 383074 96512
rect 568574 96500 568580 96512
rect 568632 96500 568638 96552
rect 165522 95888 165528 95940
rect 165580 95928 165586 95940
rect 214006 95928 214012 95940
rect 165580 95900 214012 95928
rect 165580 95888 165586 95900
rect 214006 95888 214012 95900
rect 214064 95888 214070 95940
rect 261478 95888 261484 95940
rect 261536 95928 261542 95940
rect 292574 95928 292580 95940
rect 261536 95900 292580 95928
rect 261536 95888 261542 95900
rect 292574 95888 292580 95900
rect 292632 95888 292638 95940
rect 367922 95412 367928 95464
rect 367980 95452 367986 95464
rect 392578 95452 392584 95464
rect 367980 95424 392584 95452
rect 367980 95412 367986 95424
rect 392578 95412 392584 95424
rect 392636 95412 392642 95464
rect 385770 95344 385776 95396
rect 385828 95384 385834 95396
rect 427998 95384 428004 95396
rect 385828 95356 428004 95384
rect 385828 95344 385834 95356
rect 427998 95344 428004 95356
rect 428056 95344 428062 95396
rect 380250 95276 380256 95328
rect 380308 95316 380314 95328
rect 500770 95316 500776 95328
rect 380308 95288 500776 95316
rect 380308 95276 380314 95288
rect 500770 95276 500776 95288
rect 500828 95276 500834 95328
rect 172054 95208 172060 95260
rect 172112 95248 172118 95260
rect 213914 95248 213920 95260
rect 172112 95220 213920 95248
rect 172112 95208 172118 95220
rect 213914 95208 213920 95220
rect 213972 95208 213978 95260
rect 249058 95208 249064 95260
rect 249116 95248 249122 95260
rect 307662 95248 307668 95260
rect 249116 95220 307668 95248
rect 249116 95208 249122 95220
rect 307662 95208 307668 95220
rect 307720 95208 307726 95260
rect 355318 95208 355324 95260
rect 355376 95248 355382 95260
rect 507210 95248 507216 95260
rect 355376 95220 507216 95248
rect 355376 95208 355382 95220
rect 507210 95208 507216 95220
rect 507268 95208 507274 95260
rect 523310 95208 523316 95260
rect 523368 95248 523374 95260
rect 578234 95248 578240 95260
rect 523368 95220 578240 95248
rect 523368 95208 523374 95220
rect 578234 95208 578240 95220
rect 578292 95208 578298 95260
rect 174538 95140 174544 95192
rect 174596 95180 174602 95192
rect 324682 95180 324688 95192
rect 174596 95152 324688 95180
rect 174596 95140 174602 95152
rect 324682 95140 324688 95152
rect 324740 95140 324746 95192
rect 388714 95140 388720 95192
rect 388772 95180 388778 95192
rect 399018 95180 399024 95192
rect 388772 95152 399024 95180
rect 388772 95140 388778 95152
rect 399018 95140 399024 95152
rect 399076 95140 399082 95192
rect 548426 95140 548432 95192
rect 548484 95180 548490 95192
rect 576118 95180 576124 95192
rect 548484 95152 576124 95180
rect 548484 95140 548490 95152
rect 576118 95140 576124 95152
rect 576176 95140 576182 95192
rect 207658 95072 207664 95124
rect 207716 95112 207722 95124
rect 325694 95112 325700 95124
rect 207716 95084 325700 95112
rect 207716 95072 207722 95084
rect 325694 95072 325700 95084
rect 325752 95072 325758 95124
rect 385678 95072 385684 95124
rect 385736 95112 385742 95124
rect 395798 95112 395804 95124
rect 385736 95084 395804 95112
rect 385736 95072 385742 95084
rect 395798 95072 395804 95084
rect 395856 95072 395862 95124
rect 418338 95072 418344 95124
rect 418396 95112 418402 95124
rect 574738 95112 574744 95124
rect 418396 95084 574744 95112
rect 418396 95072 418402 95084
rect 574738 95072 574744 95084
rect 574796 95072 574802 95124
rect 331950 95004 331956 95056
rect 332008 95044 332014 95056
rect 424778 95044 424784 95056
rect 332008 95016 424784 95044
rect 332008 95004 332014 95016
rect 424778 95004 424784 95016
rect 424836 95004 424842 95056
rect 541986 95004 541992 95056
rect 542044 95044 542050 95056
rect 569218 95044 569224 95056
rect 542044 95016 569224 95044
rect 542044 95004 542050 95016
rect 569218 95004 569224 95016
rect 569276 95004 569282 95056
rect 382918 94936 382924 94988
rect 382976 94976 382982 94988
rect 437014 94976 437020 94988
rect 382976 94948 437020 94976
rect 382976 94936 382982 94948
rect 437014 94936 437020 94948
rect 437072 94936 437078 94988
rect 322934 94868 322940 94920
rect 322992 94908 322998 94920
rect 513650 94908 513656 94920
rect 322992 94880 513656 94908
rect 322992 94868 322998 94880
rect 513650 94868 513656 94880
rect 513708 94868 513714 94920
rect 388622 94800 388628 94852
rect 388680 94840 388686 94852
rect 421558 94840 421564 94852
rect 388680 94812 421564 94840
rect 388680 94800 388686 94812
rect 421558 94800 421564 94812
rect 421616 94800 421622 94852
rect 126882 94460 126888 94512
rect 126940 94500 126946 94512
rect 214098 94500 214104 94512
rect 126940 94472 214104 94500
rect 126940 94460 126946 94472
rect 214098 94460 214104 94472
rect 214156 94460 214162 94512
rect 246298 94460 246304 94512
rect 246356 94500 246362 94512
rect 257706 94500 257712 94512
rect 246356 94472 257712 94500
rect 246356 94460 246362 94472
rect 257706 94460 257712 94472
rect 257764 94460 257770 94512
rect 151906 94052 151912 94104
rect 151964 94092 151970 94104
rect 171778 94092 171784 94104
rect 151964 94064 171784 94092
rect 151964 94052 151970 94064
rect 171778 94052 171784 94064
rect 171836 94052 171842 94104
rect 123202 93984 123208 94036
rect 123260 94024 123266 94036
rect 173342 94024 173348 94036
rect 123260 93996 173348 94024
rect 123260 93984 123266 93996
rect 173342 93984 173348 93996
rect 173400 93984 173406 94036
rect 112346 93916 112352 93968
rect 112404 93956 112410 93968
rect 166442 93956 166448 93968
rect 112404 93928 166448 93956
rect 112404 93916 112410 93928
rect 166442 93916 166448 93928
rect 166500 93916 166506 93968
rect 113174 93848 113180 93900
rect 113232 93888 113238 93900
rect 169110 93888 169116 93900
rect 113232 93860 169116 93888
rect 113232 93848 113238 93860
rect 169110 93848 169116 93860
rect 169168 93848 169174 93900
rect 322934 93888 322940 93900
rect 322860 93860 322940 93888
rect 67634 93780 67640 93832
rect 67692 93820 67698 93832
rect 205082 93820 205088 93832
rect 67692 93792 205088 93820
rect 67692 93780 67698 93792
rect 205082 93780 205088 93792
rect 205140 93780 205146 93832
rect 217410 93780 217416 93832
rect 217468 93820 217474 93832
rect 322860 93820 322888 93860
rect 322934 93848 322940 93860
rect 322992 93848 322998 93900
rect 325694 93848 325700 93900
rect 325752 93888 325758 93900
rect 325752 93860 328454 93888
rect 325752 93848 325758 93860
rect 217468 93792 322888 93820
rect 217468 93780 217474 93792
rect 328426 93752 328454 93860
rect 564526 93780 564532 93832
rect 564584 93820 564590 93832
rect 582926 93820 582932 93832
rect 564584 93792 582932 93820
rect 564584 93780 564590 93792
rect 582926 93780 582932 93792
rect 582984 93780 582990 93832
rect 443454 93752 443460 93764
rect 328426 93724 443460 93752
rect 443454 93712 443460 93724
rect 443512 93712 443518 93764
rect 456334 93712 456340 93764
rect 456392 93752 456398 93764
rect 582374 93752 582380 93764
rect 456392 93724 582380 93752
rect 456392 93712 456398 93724
rect 582374 93712 582380 93724
rect 582432 93712 582438 93764
rect 384298 93644 384304 93696
rect 384356 93684 384362 93696
rect 475654 93684 475660 93696
rect 384356 93656 475660 93684
rect 384356 93644 384362 93656
rect 475654 93644 475660 93656
rect 475712 93644 475718 93696
rect 487798 93644 487804 93696
rect 487856 93684 487862 93696
rect 573358 93684 573364 93696
rect 487856 93656 573364 93684
rect 487856 93644 487862 93656
rect 573358 93644 573364 93656
rect 573416 93644 573422 93696
rect 356790 93576 356796 93628
rect 356848 93616 356854 93628
rect 402238 93616 402244 93628
rect 356848 93588 402244 93616
rect 356848 93576 356854 93588
rect 402238 93576 402244 93588
rect 402296 93576 402302 93628
rect 529750 93576 529756 93628
rect 529808 93616 529814 93628
rect 569310 93616 569316 93628
rect 529808 93588 569316 93616
rect 529808 93576 529814 93588
rect 569310 93576 569316 93588
rect 569368 93576 569374 93628
rect 387150 93508 387156 93560
rect 387208 93548 387214 93560
rect 415118 93548 415124 93560
rect 387208 93520 415124 93548
rect 387208 93508 387214 93520
rect 415118 93508 415124 93520
rect 415176 93508 415182 93560
rect 567746 93508 567752 93560
rect 567804 93548 567810 93560
rect 582834 93548 582840 93560
rect 567804 93520 582840 93548
rect 567804 93508 567810 93520
rect 582834 93508 582840 93520
rect 582892 93508 582898 93560
rect 385862 93440 385868 93492
rect 385920 93480 385926 93492
rect 411898 93480 411904 93492
rect 385920 93452 411904 93480
rect 385920 93440 385926 93452
rect 411898 93440 411904 93452
rect 411956 93440 411962 93492
rect 376018 93372 376024 93424
rect 376076 93412 376082 93424
rect 572714 93412 572720 93424
rect 376076 93384 572720 93412
rect 376076 93372 376082 93384
rect 572714 93372 572720 93384
rect 572772 93372 572778 93424
rect 121730 93304 121736 93356
rect 121788 93344 121794 93356
rect 167730 93344 167736 93356
rect 121788 93316 167736 93344
rect 121788 93304 121794 93316
rect 167730 93304 167736 93316
rect 167788 93304 167794 93356
rect 151538 93236 151544 93288
rect 151596 93276 151602 93288
rect 202230 93276 202236 93288
rect 151596 93248 202236 93276
rect 151596 93236 151602 93248
rect 202230 93236 202236 93248
rect 202288 93236 202294 93288
rect 93946 93168 93952 93220
rect 94004 93208 94010 93220
rect 207842 93208 207848 93220
rect 94004 93180 207848 93208
rect 94004 93168 94010 93180
rect 207842 93168 207848 93180
rect 207900 93168 207906 93220
rect 107746 93100 107752 93152
rect 107804 93140 107810 93152
rect 193950 93140 193956 93152
rect 107804 93112 193956 93140
rect 107804 93100 107810 93112
rect 193950 93100 193956 93112
rect 194008 93100 194014 93152
rect 206370 93100 206376 93152
rect 206428 93140 206434 93152
rect 324314 93140 324320 93152
rect 206428 93112 324320 93140
rect 206428 93100 206434 93112
rect 324314 93100 324320 93112
rect 324372 93100 324378 93152
rect 88978 92420 88984 92472
rect 89036 92460 89042 92472
rect 165522 92460 165528 92472
rect 89036 92432 165528 92460
rect 89036 92420 89042 92432
rect 165522 92420 165528 92432
rect 165580 92420 165586 92472
rect 380342 92420 380348 92472
rect 380400 92460 380406 92472
rect 576854 92460 576860 92472
rect 380400 92432 576860 92460
rect 380400 92420 380406 92432
rect 576854 92420 576860 92432
rect 576912 92420 576918 92472
rect 118050 92352 118056 92404
rect 118108 92392 118114 92404
rect 188430 92392 188436 92404
rect 118108 92364 188436 92392
rect 118108 92352 118114 92364
rect 188430 92352 188436 92364
rect 188488 92352 188494 92404
rect 388438 92352 388444 92404
rect 388496 92392 388502 92404
rect 571426 92392 571432 92404
rect 388496 92364 571432 92392
rect 388496 92352 388502 92364
rect 571426 92352 571432 92364
rect 571484 92352 571490 92404
rect 87230 92284 87236 92336
rect 87288 92324 87294 92336
rect 126882 92324 126888 92336
rect 87288 92296 126888 92324
rect 87288 92284 87294 92296
rect 126882 92284 126888 92296
rect 126940 92284 126946 92336
rect 129458 92284 129464 92336
rect 129516 92324 129522 92336
rect 189810 92324 189816 92336
rect 129516 92296 189816 92324
rect 129516 92284 129522 92296
rect 189810 92284 189816 92296
rect 189868 92284 189874 92336
rect 387702 92284 387708 92336
rect 387760 92324 387766 92336
rect 570598 92324 570604 92336
rect 387760 92296 570604 92324
rect 387760 92284 387766 92296
rect 570598 92284 570604 92296
rect 570656 92284 570662 92336
rect 107470 92216 107476 92268
rect 107528 92256 107534 92268
rect 128354 92256 128360 92268
rect 107528 92228 128360 92256
rect 107528 92216 107534 92228
rect 128354 92216 128360 92228
rect 128412 92216 128418 92268
rect 135714 92216 135720 92268
rect 135772 92256 135778 92268
rect 193858 92256 193864 92268
rect 135772 92228 193864 92256
rect 135772 92216 135778 92228
rect 193858 92216 193864 92228
rect 193916 92216 193922 92268
rect 360838 92216 360844 92268
rect 360896 92256 360902 92268
rect 509878 92256 509884 92268
rect 360896 92228 509884 92256
rect 360896 92216 360902 92228
rect 509878 92216 509884 92228
rect 509936 92256 509942 92268
rect 510522 92256 510528 92268
rect 509936 92228 510528 92256
rect 509936 92216 509942 92228
rect 510522 92216 510528 92228
rect 510580 92216 510586 92268
rect 114186 92148 114192 92200
rect 114244 92188 114250 92200
rect 169294 92188 169300 92200
rect 114244 92160 169300 92188
rect 114244 92148 114250 92160
rect 169294 92148 169300 92160
rect 169352 92148 169358 92200
rect 351178 92148 351184 92200
rect 351236 92188 351242 92200
rect 418338 92188 418344 92200
rect 351236 92160 418344 92188
rect 351236 92148 351242 92160
rect 418338 92148 418344 92160
rect 418396 92148 418402 92200
rect 449894 92148 449900 92200
rect 449952 92188 449958 92200
rect 576210 92188 576216 92200
rect 449952 92160 576216 92188
rect 449952 92148 449958 92160
rect 576210 92148 576216 92160
rect 576268 92148 576274 92200
rect 125778 92080 125784 92132
rect 125836 92120 125842 92132
rect 166534 92120 166540 92132
rect 125836 92092 166540 92120
rect 125836 92080 125842 92092
rect 166534 92080 166540 92092
rect 166592 92080 166598 92132
rect 381538 92080 381544 92132
rect 381596 92120 381602 92132
rect 446674 92120 446680 92132
rect 381596 92092 446680 92120
rect 381596 92080 381602 92092
rect 446674 92080 446680 92092
rect 446732 92080 446738 92132
rect 238018 91876 238024 91928
rect 238076 91916 238082 91928
rect 250990 91916 250996 91928
rect 238076 91888 250996 91916
rect 238076 91876 238082 91888
rect 250990 91876 250996 91888
rect 251048 91876 251054 91928
rect 166994 91808 167000 91860
rect 167052 91848 167058 91860
rect 204898 91848 204904 91860
rect 167052 91820 204904 91848
rect 167052 91808 167058 91820
rect 204898 91808 204904 91820
rect 204956 91808 204962 91860
rect 228358 91808 228364 91860
rect 228416 91848 228422 91860
rect 260374 91848 260380 91860
rect 228416 91820 260380 91848
rect 228416 91808 228422 91820
rect 260374 91808 260380 91820
rect 260432 91808 260438 91860
rect 198734 91740 198740 91792
rect 198792 91780 198798 91792
rect 276106 91780 276112 91792
rect 198792 91752 276112 91780
rect 198792 91740 198798 91752
rect 276106 91740 276112 91752
rect 276164 91740 276170 91792
rect 430482 91740 430488 91792
rect 430540 91780 430546 91792
rect 431218 91780 431224 91792
rect 430540 91752 431224 91780
rect 430540 91740 430546 91752
rect 431218 91740 431224 91752
rect 431276 91740 431282 91792
rect 109678 91128 109684 91180
rect 109736 91168 109742 91180
rect 116670 91168 116676 91180
rect 109736 91140 116676 91168
rect 109736 91128 109742 91140
rect 116670 91128 116676 91140
rect 116728 91128 116734 91180
rect 85758 91060 85764 91112
rect 85816 91100 85822 91112
rect 116578 91100 116584 91112
rect 85816 91072 116584 91100
rect 85816 91060 85822 91072
rect 116578 91060 116584 91072
rect 116636 91060 116642 91112
rect 64782 90992 64788 91044
rect 64840 91032 64846 91044
rect 198274 91032 198280 91044
rect 64840 91004 198280 91032
rect 64840 90992 64846 91004
rect 198274 90992 198280 91004
rect 198332 90992 198338 91044
rect 324314 90992 324320 91044
rect 324372 91032 324378 91044
rect 569954 91032 569960 91044
rect 324372 91004 569960 91032
rect 324372 90992 324378 91004
rect 569954 90992 569960 91004
rect 570012 90992 570018 91044
rect 111610 90924 111616 90976
rect 111668 90964 111674 90976
rect 195330 90964 195336 90976
rect 111668 90936 195336 90964
rect 111668 90924 111674 90936
rect 195330 90924 195336 90936
rect 195388 90924 195394 90976
rect 469214 90924 469220 90976
rect 469272 90964 469278 90976
rect 577498 90964 577504 90976
rect 469272 90936 577504 90964
rect 469272 90924 469278 90936
rect 577498 90924 577504 90936
rect 577556 90924 577562 90976
rect 100478 90856 100484 90908
rect 100536 90896 100542 90908
rect 169202 90896 169208 90908
rect 100536 90868 169208 90896
rect 100536 90856 100542 90868
rect 169202 90856 169208 90868
rect 169260 90856 169266 90908
rect 378778 90856 378784 90908
rect 378836 90896 378842 90908
rect 478874 90896 478880 90908
rect 378836 90868 478880 90896
rect 378836 90856 378842 90868
rect 478874 90856 478880 90868
rect 478932 90856 478938 90908
rect 124490 90788 124496 90840
rect 124548 90828 124554 90840
rect 186958 90828 186964 90840
rect 124548 90800 186964 90828
rect 124548 90788 124554 90800
rect 186958 90788 186964 90800
rect 187016 90788 187022 90840
rect 387242 90788 387248 90840
rect 387300 90828 387306 90840
rect 434438 90828 434444 90840
rect 387300 90800 434444 90828
rect 387300 90788 387306 90800
rect 434438 90788 434444 90800
rect 434496 90788 434502 90840
rect 125410 90720 125416 90772
rect 125468 90760 125474 90772
rect 173434 90760 173440 90772
rect 125468 90732 173440 90760
rect 125468 90720 125474 90732
rect 173434 90720 173440 90732
rect 173492 90720 173498 90772
rect 388530 90720 388536 90772
rect 388588 90760 388594 90772
rect 472434 90760 472440 90772
rect 388588 90732 472440 90760
rect 388588 90720 388594 90732
rect 472434 90720 472440 90732
rect 472492 90720 472498 90772
rect 151722 90652 151728 90704
rect 151780 90692 151786 90704
rect 177298 90692 177304 90704
rect 151780 90664 177304 90692
rect 151780 90652 151786 90664
rect 177298 90652 177304 90664
rect 177356 90652 177362 90704
rect 308398 90312 308404 90364
rect 308456 90352 308462 90364
rect 317414 90352 317420 90364
rect 308456 90324 317420 90352
rect 308456 90312 308462 90324
rect 317414 90312 317420 90324
rect 317472 90312 317478 90364
rect 63310 89632 63316 89684
rect 63368 89672 63374 89684
rect 200758 89672 200764 89684
rect 63368 89644 200764 89672
rect 63368 89632 63374 89644
rect 200758 89632 200764 89644
rect 200816 89632 200822 89684
rect 217318 89632 217324 89684
rect 217376 89672 217382 89684
rect 327074 89672 327080 89684
rect 217376 89644 327080 89672
rect 217376 89632 217382 89644
rect 327074 89632 327080 89644
rect 327132 89672 327138 89684
rect 328362 89672 328368 89684
rect 327132 89644 328368 89672
rect 327132 89632 327138 89644
rect 328362 89632 328368 89644
rect 328420 89632 328426 89684
rect 378962 89632 378968 89684
rect 379020 89672 379026 89684
rect 554866 89672 554872 89684
rect 379020 89644 554872 89672
rect 379020 89632 379026 89644
rect 554866 89632 554872 89644
rect 554924 89632 554930 89684
rect 115382 89564 115388 89616
rect 115440 89604 115446 89616
rect 210602 89604 210608 89616
rect 115440 89576 210608 89604
rect 115440 89564 115446 89576
rect 210602 89564 210608 89576
rect 210660 89564 210666 89616
rect 363690 89564 363696 89616
rect 363748 89604 363754 89616
rect 526530 89604 526536 89616
rect 363748 89576 526536 89604
rect 363748 89564 363754 89576
rect 526530 89564 526536 89576
rect 526588 89564 526594 89616
rect 128170 89496 128176 89548
rect 128228 89536 128234 89548
rect 212074 89536 212080 89548
rect 128228 89508 212080 89536
rect 128228 89496 128234 89508
rect 212074 89496 212080 89508
rect 212132 89496 212138 89548
rect 429194 89496 429200 89548
rect 429252 89536 429258 89548
rect 430482 89536 430488 89548
rect 429252 89508 430488 89536
rect 429252 89496 429258 89508
rect 430482 89496 430488 89508
rect 430540 89536 430546 89548
rect 583846 89536 583852 89548
rect 430540 89508 583852 89536
rect 430540 89496 430546 89508
rect 583846 89496 583852 89508
rect 583904 89496 583910 89548
rect 104250 89428 104256 89480
rect 104308 89468 104314 89480
rect 171962 89468 171968 89480
rect 104308 89440 171968 89468
rect 104308 89428 104314 89440
rect 171962 89428 171968 89440
rect 172020 89428 172026 89480
rect 354030 89428 354036 89480
rect 354088 89468 354094 89480
rect 482094 89468 482100 89480
rect 354088 89440 482100 89468
rect 354088 89428 354094 89440
rect 482094 89428 482100 89440
rect 482152 89428 482158 89480
rect 151354 89360 151360 89412
rect 151412 89400 151418 89412
rect 192478 89400 192484 89412
rect 151412 89372 192484 89400
rect 151412 89360 151418 89372
rect 192478 89360 192484 89372
rect 192536 89360 192542 89412
rect 359458 89360 359464 89412
rect 359516 89400 359522 89412
rect 440234 89400 440240 89412
rect 359516 89372 440240 89400
rect 359516 89360 359522 89372
rect 440234 89360 440240 89372
rect 440292 89360 440298 89412
rect 132218 89292 132224 89344
rect 132276 89332 132282 89344
rect 166994 89332 167000 89344
rect 132276 89304 167000 89332
rect 132276 89292 132282 89304
rect 166994 89292 167000 89304
rect 167052 89292 167058 89344
rect 211890 88952 211896 89004
rect 211948 88992 211954 89004
rect 307294 88992 307300 89004
rect 211948 88964 307300 88992
rect 211948 88952 211954 88964
rect 307294 88952 307300 88964
rect 307352 88952 307358 89004
rect 206278 88272 206284 88324
rect 206336 88312 206342 88324
rect 429194 88312 429200 88324
rect 206336 88284 429200 88312
rect 206336 88272 206342 88284
rect 429194 88272 429200 88284
rect 429252 88272 429258 88324
rect 90726 88204 90732 88256
rect 90784 88244 90790 88256
rect 203702 88244 203708 88256
rect 90784 88216 203708 88244
rect 90784 88204 90790 88216
rect 203702 88204 203708 88216
rect 203760 88204 203766 88256
rect 369210 88204 369216 88256
rect 369268 88244 369274 88256
rect 571610 88244 571616 88256
rect 369268 88216 571616 88244
rect 369268 88204 369274 88216
rect 571610 88204 571616 88216
rect 571668 88204 571674 88256
rect 117130 88136 117136 88188
rect 117188 88176 117194 88188
rect 182910 88176 182916 88188
rect 117188 88148 182916 88176
rect 117188 88136 117194 88148
rect 182910 88136 182916 88148
rect 182968 88136 182974 88188
rect 328362 88136 328368 88188
rect 328420 88176 328426 88188
rect 459554 88176 459560 88188
rect 328420 88148 459560 88176
rect 328420 88136 328426 88148
rect 459554 88136 459560 88148
rect 459612 88136 459618 88188
rect 133138 88068 133144 88120
rect 133196 88108 133202 88120
rect 185578 88108 185584 88120
rect 133196 88080 185584 88108
rect 133196 88068 133202 88080
rect 185578 88068 185584 88080
rect 185636 88068 185642 88120
rect 383102 88068 383108 88120
rect 383160 88108 383166 88120
rect 462774 88108 462780 88120
rect 383160 88080 462780 88108
rect 383160 88068 383166 88080
rect 462774 88068 462780 88080
rect 462832 88068 462838 88120
rect 120718 88000 120724 88052
rect 120776 88040 120782 88052
rect 170582 88040 170588 88052
rect 120776 88012 170588 88040
rect 120776 88000 120782 88012
rect 170582 88000 170588 88012
rect 170640 88000 170646 88052
rect 64690 87932 64696 87984
rect 64748 87972 64754 87984
rect 207934 87972 207940 87984
rect 64748 87944 207940 87972
rect 64748 87932 64754 87944
rect 207934 87932 207940 87944
rect 207992 87932 207998 87984
rect 184198 87592 184204 87644
rect 184256 87632 184262 87644
rect 233878 87632 233884 87644
rect 184256 87604 233884 87632
rect 184256 87592 184262 87604
rect 233878 87592 233884 87604
rect 233936 87592 233942 87644
rect 302878 87592 302884 87644
rect 302936 87632 302942 87644
rect 324498 87632 324504 87644
rect 302936 87604 324504 87632
rect 302936 87592 302942 87604
rect 324498 87592 324504 87604
rect 324556 87592 324562 87644
rect 67726 86912 67732 86964
rect 67784 86952 67790 86964
rect 214834 86952 214840 86964
rect 67784 86924 214840 86952
rect 67784 86912 67790 86924
rect 214834 86912 214840 86924
rect 214892 86912 214898 86964
rect 327902 86912 327908 86964
rect 327960 86952 327966 86964
rect 560294 86952 560300 86964
rect 327960 86924 560300 86952
rect 327960 86912 327966 86924
rect 560294 86912 560300 86924
rect 560352 86912 560358 86964
rect 573450 86912 573456 86964
rect 573508 86952 573514 86964
rect 580166 86952 580172 86964
rect 573508 86924 580172 86952
rect 573508 86912 573514 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 63402 86844 63408 86896
rect 63460 86884 63466 86896
rect 198182 86884 198188 86896
rect 63460 86856 198188 86884
rect 63460 86844 63466 86856
rect 198182 86844 198188 86856
rect 198240 86844 198246 86896
rect 384390 86844 384396 86896
rect 384448 86884 384454 86896
rect 489914 86884 489920 86896
rect 384448 86856 489920 86884
rect 384448 86844 384454 86856
rect 489914 86844 489920 86856
rect 489972 86844 489978 86896
rect 110138 86776 110144 86828
rect 110196 86816 110202 86828
rect 203610 86816 203616 86828
rect 110196 86788 203616 86816
rect 110196 86776 110202 86788
rect 203610 86776 203616 86788
rect 203668 86776 203674 86828
rect 381722 86776 381728 86828
rect 381780 86816 381786 86828
rect 465074 86816 465080 86828
rect 381780 86788 465080 86816
rect 381780 86776 381786 86788
rect 465074 86776 465080 86788
rect 465132 86776 465138 86828
rect 118234 86708 118240 86760
rect 118292 86748 118298 86760
rect 184290 86748 184296 86760
rect 118292 86720 184296 86748
rect 118292 86708 118298 86720
rect 184290 86708 184296 86720
rect 184348 86708 184354 86760
rect 130746 86640 130752 86692
rect 130804 86680 130810 86692
rect 167638 86680 167644 86692
rect 130804 86652 167644 86680
rect 130804 86640 130810 86652
rect 167638 86640 167644 86652
rect 167696 86640 167702 86692
rect 253198 86300 253204 86352
rect 253256 86340 253262 86352
rect 266354 86340 266360 86352
rect 253256 86312 266360 86340
rect 253256 86300 253262 86312
rect 266354 86300 266360 86312
rect 266412 86300 266418 86352
rect 242894 86232 242900 86284
rect 242952 86272 242958 86284
rect 293954 86272 293960 86284
rect 242952 86244 293960 86272
rect 242952 86232 242958 86244
rect 293954 86232 293960 86244
rect 294012 86232 294018 86284
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 26878 85524 26884 85536
rect 3200 85496 26884 85524
rect 3200 85484 3206 85496
rect 26878 85484 26884 85496
rect 26936 85484 26942 85536
rect 113910 85484 113916 85536
rect 113968 85524 113974 85536
rect 212166 85524 212172 85536
rect 113968 85496 212172 85524
rect 113968 85484 113974 85496
rect 212166 85484 212172 85496
rect 212224 85484 212230 85536
rect 329190 85484 329196 85536
rect 329248 85524 329254 85536
rect 531314 85524 531320 85536
rect 329248 85496 531320 85524
rect 329248 85484 329254 85496
rect 531314 85484 531320 85496
rect 531372 85484 531378 85536
rect 101858 85416 101864 85468
rect 101916 85456 101922 85468
rect 192662 85456 192668 85468
rect 101916 85428 192668 85456
rect 101916 85416 101922 85428
rect 192662 85416 192668 85428
rect 192720 85416 192726 85468
rect 338758 85416 338764 85468
rect 338816 85456 338822 85468
rect 487798 85456 487804 85468
rect 338816 85428 487804 85456
rect 338816 85416 338822 85428
rect 487798 85416 487804 85428
rect 487856 85416 487862 85468
rect 108482 85348 108488 85400
rect 108540 85388 108546 85400
rect 173250 85388 173256 85400
rect 108540 85360 173256 85388
rect 108540 85348 108546 85360
rect 173250 85348 173256 85360
rect 173308 85348 173314 85400
rect 385954 85348 385960 85400
rect 386012 85388 386018 85400
rect 496814 85388 496820 85400
rect 386012 85360 496820 85388
rect 386012 85348 386018 85360
rect 496814 85348 496820 85360
rect 496872 85348 496878 85400
rect 119890 85280 119896 85332
rect 119948 85320 119954 85332
rect 171870 85320 171876 85332
rect 119948 85292 171876 85320
rect 119948 85280 119954 85292
rect 171870 85280 171876 85292
rect 171928 85280 171934 85332
rect 360930 85280 360936 85332
rect 360988 85320 360994 85332
rect 452654 85320 452660 85332
rect 360988 85292 452660 85320
rect 360988 85280 360994 85292
rect 452654 85280 452660 85292
rect 452712 85280 452718 85332
rect 124030 85212 124036 85264
rect 124088 85252 124094 85264
rect 166350 85252 166356 85264
rect 124088 85224 166356 85252
rect 124088 85212 124094 85224
rect 166350 85212 166356 85224
rect 166408 85212 166414 85264
rect 134702 85144 134708 85196
rect 134760 85184 134766 85196
rect 166258 85184 166264 85196
rect 134760 85156 166264 85184
rect 134760 85144 134766 85156
rect 166258 85144 166264 85156
rect 166316 85144 166322 85196
rect 176378 84804 176384 84856
rect 176436 84844 176442 84856
rect 267734 84844 267740 84856
rect 176436 84816 267740 84844
rect 176436 84804 176442 84816
rect 267734 84804 267740 84816
rect 267792 84804 267798 84856
rect 510522 84804 510528 84856
rect 510580 84844 510586 84856
rect 522298 84844 522304 84856
rect 510580 84816 522304 84844
rect 510580 84804 510586 84816
rect 522298 84804 522304 84816
rect 522356 84804 522362 84856
rect 99098 84124 99104 84176
rect 99156 84164 99162 84176
rect 206462 84164 206468 84176
rect 99156 84136 206468 84164
rect 99156 84124 99162 84136
rect 206462 84124 206468 84136
rect 206520 84124 206526 84176
rect 359550 84124 359556 84176
rect 359608 84164 359614 84176
rect 557534 84164 557540 84176
rect 359608 84136 557540 84164
rect 359608 84124 359614 84136
rect 557534 84124 557540 84136
rect 557592 84124 557598 84176
rect 107562 84056 107568 84108
rect 107620 84096 107626 84108
rect 210418 84096 210424 84108
rect 107620 84068 210424 84096
rect 107620 84056 107626 84068
rect 210418 84056 210424 84068
rect 210476 84056 210482 84108
rect 374730 84056 374736 84108
rect 374788 84096 374794 84108
rect 516134 84096 516140 84108
rect 374788 84068 516140 84096
rect 374788 84056 374794 84068
rect 516134 84056 516140 84068
rect 516192 84056 516198 84108
rect 96522 83988 96528 84040
rect 96580 84028 96586 84040
rect 167914 84028 167920 84040
rect 96580 84000 167920 84028
rect 96580 83988 96586 84000
rect 167914 83988 167920 84000
rect 167972 83988 167978 84040
rect 115842 83920 115848 83972
rect 115900 83960 115906 83972
rect 187050 83960 187056 83972
rect 115900 83932 187056 83960
rect 115900 83920 115906 83932
rect 187050 83920 187056 83932
rect 187108 83920 187114 83972
rect 124122 83852 124128 83904
rect 124180 83892 124186 83904
rect 170490 83892 170496 83904
rect 124180 83864 170496 83892
rect 124180 83852 124186 83864
rect 170490 83852 170496 83864
rect 170548 83852 170554 83904
rect 212534 83444 212540 83496
rect 212592 83484 212598 83496
rect 327074 83484 327080 83496
rect 212592 83456 327080 83484
rect 212592 83444 212598 83456
rect 327074 83444 327080 83456
rect 327132 83444 327138 83496
rect 67266 82764 67272 82816
rect 67324 82804 67330 82816
rect 324406 82804 324412 82816
rect 67324 82776 324412 82804
rect 67324 82764 67330 82776
rect 324406 82764 324412 82776
rect 324464 82764 324470 82816
rect 358078 82764 358084 82816
rect 358136 82804 358142 82816
rect 548518 82804 548524 82816
rect 358136 82776 548524 82804
rect 358136 82764 358142 82776
rect 548518 82764 548524 82776
rect 548576 82764 548582 82816
rect 97902 82696 97908 82748
rect 97960 82736 97966 82748
rect 209038 82736 209044 82748
rect 97960 82708 209044 82736
rect 97960 82696 97966 82708
rect 209038 82696 209044 82708
rect 209096 82696 209102 82748
rect 367738 82696 367744 82748
rect 367796 82736 367802 82748
rect 503714 82736 503720 82748
rect 367796 82708 503720 82736
rect 367796 82696 367802 82708
rect 503714 82696 503720 82708
rect 503772 82696 503778 82748
rect 111702 82628 111708 82680
rect 111760 82668 111766 82680
rect 207750 82668 207756 82680
rect 111760 82640 207756 82668
rect 111760 82628 111766 82640
rect 207750 82628 207756 82640
rect 207808 82628 207814 82680
rect 377490 82628 377496 82680
rect 377548 82668 377554 82680
rect 494054 82668 494060 82680
rect 377548 82640 494060 82668
rect 377548 82628 377554 82640
rect 494054 82628 494060 82640
rect 494112 82628 494118 82680
rect 103330 82560 103336 82612
rect 103388 82600 103394 82612
rect 184382 82600 184388 82612
rect 103388 82572 184388 82600
rect 103388 82560 103394 82572
rect 184382 82560 184388 82572
rect 184440 82560 184446 82612
rect 46842 81336 46848 81388
rect 46900 81376 46906 81388
rect 321554 81376 321560 81388
rect 46900 81348 321560 81376
rect 46900 81336 46906 81348
rect 321554 81336 321560 81348
rect 321612 81376 321618 81388
rect 582742 81376 582748 81388
rect 321612 81348 582748 81376
rect 321612 81336 321618 81348
rect 582742 81336 582748 81348
rect 582800 81336 582806 81388
rect 92382 81268 92388 81320
rect 92440 81308 92446 81320
rect 185670 81308 185676 81320
rect 92440 81280 185676 81308
rect 92440 81268 92446 81280
rect 185670 81268 185676 81280
rect 185728 81268 185734 81320
rect 333882 81268 333888 81320
rect 333940 81308 333946 81320
rect 518894 81308 518900 81320
rect 333940 81280 518900 81308
rect 333940 81268 333946 81280
rect 518894 81268 518900 81280
rect 518952 81268 518958 81320
rect 126882 81200 126888 81252
rect 126940 81240 126946 81252
rect 210510 81240 210516 81252
rect 126940 81212 210516 81240
rect 126940 81200 126946 81212
rect 210510 81200 210516 81212
rect 210568 81200 210574 81252
rect 373442 81200 373448 81252
rect 373500 81240 373506 81252
rect 550634 81240 550640 81252
rect 373500 81212 550640 81240
rect 373500 81200 373506 81212
rect 550634 81200 550640 81212
rect 550692 81200 550698 81252
rect 126790 81132 126796 81184
rect 126848 81172 126854 81184
rect 196802 81172 196808 81184
rect 126848 81144 196808 81172
rect 126848 81132 126854 81144
rect 196802 81132 196808 81144
rect 196860 81132 196866 81184
rect 210418 80656 210424 80708
rect 210476 80696 210482 80708
rect 307202 80696 307208 80708
rect 210476 80668 307208 80696
rect 210476 80656 210482 80668
rect 307202 80656 307208 80668
rect 307260 80656 307266 80708
rect 95142 79976 95148 80028
rect 95200 80016 95206 80028
rect 188522 80016 188528 80028
rect 95200 79988 188528 80016
rect 95200 79976 95206 79988
rect 188522 79976 188528 79988
rect 188580 79976 188586 80028
rect 324958 79976 324964 80028
rect 325016 80016 325022 80028
rect 570138 80016 570144 80028
rect 325016 79988 570144 80016
rect 325016 79976 325022 79988
rect 570138 79976 570144 79988
rect 570196 79976 570202 80028
rect 121362 79908 121368 79960
rect 121420 79948 121426 79960
rect 211982 79948 211988 79960
rect 121420 79920 211988 79948
rect 121420 79908 121426 79920
rect 211982 79908 211988 79920
rect 212040 79908 212046 79960
rect 365070 79908 365076 79960
rect 365128 79948 365134 79960
rect 574186 79948 574192 79960
rect 365128 79920 574192 79948
rect 365128 79908 365134 79920
rect 574186 79908 574192 79920
rect 574244 79908 574250 79960
rect 119982 79840 119988 79892
rect 120040 79880 120046 79892
rect 206554 79880 206560 79892
rect 120040 79852 206560 79880
rect 120040 79840 120046 79852
rect 206554 79840 206560 79852
rect 206612 79840 206618 79892
rect 86862 79772 86868 79824
rect 86920 79812 86926 79824
rect 167822 79812 167828 79824
rect 86920 79784 167828 79812
rect 86920 79772 86926 79784
rect 167822 79772 167828 79784
rect 167880 79772 167886 79824
rect 99190 79704 99196 79756
rect 99248 79744 99254 79756
rect 169018 79744 169024 79756
rect 99248 79716 169024 79744
rect 99248 79704 99254 79716
rect 169018 79704 169024 79716
rect 169076 79704 169082 79756
rect 238754 79364 238760 79416
rect 238812 79404 238818 79416
rect 294046 79404 294052 79416
rect 238812 79376 294052 79404
rect 238812 79364 238818 79376
rect 294046 79364 294052 79376
rect 294104 79364 294110 79416
rect 179322 79296 179328 79348
rect 179380 79336 179386 79348
rect 245654 79336 245660 79348
rect 179380 79308 245660 79336
rect 179380 79296 179386 79308
rect 245654 79296 245660 79308
rect 245712 79296 245718 79348
rect 297450 79296 297456 79348
rect 297508 79336 297514 79348
rect 320174 79336 320180 79348
rect 297508 79308 320180 79336
rect 297508 79296 297514 79308
rect 320174 79296 320180 79308
rect 320232 79296 320238 79348
rect 116670 78616 116676 78668
rect 116728 78656 116734 78668
rect 213178 78656 213184 78668
rect 116728 78628 213184 78656
rect 116728 78616 116734 78628
rect 213178 78616 213184 78628
rect 213236 78616 213242 78668
rect 276658 78616 276664 78668
rect 276716 78656 276722 78668
rect 570046 78656 570052 78668
rect 276716 78628 570052 78656
rect 276716 78616 276722 78628
rect 570046 78616 570052 78628
rect 570104 78616 570110 78668
rect 102042 78548 102048 78600
rect 102100 78588 102106 78600
rect 196710 78588 196716 78600
rect 102100 78560 196716 78588
rect 102100 78548 102106 78560
rect 196710 78548 196716 78560
rect 196768 78548 196774 78600
rect 99282 78480 99288 78532
rect 99340 78520 99346 78532
rect 189902 78520 189908 78532
rect 99340 78492 189908 78520
rect 99340 78480 99346 78492
rect 189902 78480 189908 78492
rect 189960 78480 189966 78532
rect 122742 78412 122748 78464
rect 122800 78452 122806 78464
rect 202138 78452 202144 78464
rect 122800 78424 202144 78452
rect 122800 78412 122806 78424
rect 202138 78412 202144 78424
rect 202196 78412 202202 78464
rect 93762 78344 93768 78396
rect 93820 78384 93826 78396
rect 170674 78384 170680 78396
rect 93820 78356 170680 78384
rect 93820 78344 93826 78356
rect 170674 78344 170680 78356
rect 170732 78344 170738 78396
rect 257982 78004 257988 78056
rect 258040 78044 258046 78056
rect 275462 78044 275468 78056
rect 258040 78016 275468 78044
rect 258040 78004 258046 78016
rect 275462 78004 275468 78016
rect 275520 78004 275526 78056
rect 200114 77936 200120 77988
rect 200172 77976 200178 77988
rect 311894 77976 311900 77988
rect 200172 77948 311900 77976
rect 200172 77936 200178 77948
rect 311894 77936 311900 77948
rect 311952 77936 311958 77988
rect 66898 77188 66904 77240
rect 66956 77228 66962 77240
rect 484394 77228 484400 77240
rect 66956 77200 484400 77228
rect 66956 77188 66962 77200
rect 484394 77188 484400 77200
rect 484452 77188 484458 77240
rect 75822 77120 75828 77172
rect 75880 77160 75886 77172
rect 172054 77160 172060 77172
rect 75880 77132 172060 77160
rect 75880 77120 75886 77132
rect 172054 77120 172060 77132
rect 172112 77120 172118 77172
rect 347038 77120 347044 77172
rect 347096 77160 347102 77172
rect 545114 77160 545120 77172
rect 347096 77132 545120 77160
rect 347096 77120 347102 77132
rect 545114 77120 545120 77132
rect 545172 77120 545178 77172
rect 106182 77052 106188 77104
rect 106240 77092 106246 77104
rect 177390 77092 177396 77104
rect 106240 77064 177396 77092
rect 106240 77052 106246 77064
rect 177390 77052 177396 77064
rect 177448 77052 177454 77104
rect 120074 76508 120080 76560
rect 120132 76548 120138 76560
rect 250530 76548 250536 76560
rect 120132 76520 250536 76548
rect 120132 76508 120138 76520
rect 250530 76508 250536 76520
rect 250588 76508 250594 76560
rect 100570 75828 100576 75880
rect 100628 75868 100634 75880
rect 199378 75868 199384 75880
rect 100628 75840 199384 75868
rect 100628 75828 100634 75840
rect 199378 75828 199384 75840
rect 199436 75828 199442 75880
rect 113082 75760 113088 75812
rect 113140 75800 113146 75812
rect 170398 75800 170404 75812
rect 113140 75772 170404 75800
rect 113140 75760 113146 75772
rect 170398 75760 170404 75772
rect 170456 75760 170462 75812
rect 175090 75216 175096 75268
rect 175148 75256 175154 75268
rect 331306 75256 331312 75268
rect 175148 75228 331312 75256
rect 175148 75216 175154 75228
rect 331306 75216 331312 75228
rect 331364 75216 331370 75268
rect 49694 75148 49700 75200
rect 49752 75188 49758 75200
rect 265710 75188 265716 75200
rect 49752 75160 265716 75188
rect 49752 75148 49758 75160
rect 265710 75148 265716 75160
rect 265768 75148 265774 75200
rect 116578 74468 116584 74520
rect 116636 74508 116642 74520
rect 214558 74508 214564 74520
rect 116636 74480 214564 74508
rect 116636 74468 116642 74480
rect 214558 74468 214564 74480
rect 214616 74468 214622 74520
rect 104802 74400 104808 74452
rect 104860 74440 104866 74452
rect 192570 74440 192576 74452
rect 104860 74412 192576 74440
rect 104860 74400 104866 74412
rect 192570 74400 192576 74412
rect 192628 74400 192634 74452
rect 52454 73856 52460 73908
rect 52512 73896 52518 73908
rect 301774 73896 301780 73908
rect 52512 73868 301780 73896
rect 52512 73856 52518 73868
rect 301774 73856 301780 73868
rect 301832 73856 301838 73908
rect 27614 73788 27620 73840
rect 27672 73828 27678 73840
rect 279510 73828 279516 73840
rect 27672 73800 279516 73828
rect 27672 73788 27678 73800
rect 279510 73788 279516 73800
rect 279568 73788 279574 73840
rect 85482 73108 85488 73160
rect 85540 73148 85546 73160
rect 204990 73148 204996 73160
rect 85540 73120 204996 73148
rect 85540 73108 85546 73120
rect 204990 73108 204996 73120
rect 205048 73108 205054 73160
rect 574830 73108 574836 73160
rect 574888 73148 574894 73160
rect 579982 73148 579988 73160
rect 574888 73120 579988 73148
rect 574888 73108 574894 73120
rect 579982 73108 579988 73120
rect 580040 73108 580046 73160
rect 114554 72496 114560 72548
rect 114612 72536 114618 72548
rect 274082 72536 274088 72548
rect 114612 72508 274088 72536
rect 114612 72496 114618 72508
rect 274082 72496 274088 72508
rect 274140 72496 274146 72548
rect 66254 72428 66260 72480
rect 66312 72468 66318 72480
rect 296162 72468 296168 72480
rect 66312 72440 296168 72468
rect 66312 72428 66318 72440
rect 296162 72428 296168 72440
rect 296220 72428 296226 72480
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 32398 71720 32404 71732
rect 3476 71692 32404 71720
rect 3476 71680 3482 71692
rect 32398 71680 32404 71692
rect 32456 71680 32462 71732
rect 179138 71136 179144 71188
rect 179196 71176 179202 71188
rect 296714 71176 296720 71188
rect 179196 71148 296720 71176
rect 179196 71136 179202 71148
rect 296714 71136 296720 71148
rect 296772 71136 296778 71188
rect 103514 71068 103520 71120
rect 103572 71108 103578 71120
rect 304534 71108 304540 71120
rect 103572 71080 304540 71108
rect 103572 71068 103578 71080
rect 304534 71068 304540 71080
rect 304592 71068 304598 71120
rect 30374 71000 30380 71052
rect 30432 71040 30438 71052
rect 249150 71040 249156 71052
rect 30432 71012 249156 71040
rect 30432 71000 30438 71012
rect 249150 71000 249156 71012
rect 249208 71000 249214 71052
rect 124214 69708 124220 69760
rect 124272 69748 124278 69760
rect 253382 69748 253388 69760
rect 124272 69720 253388 69748
rect 124272 69708 124278 69720
rect 253382 69708 253388 69720
rect 253440 69708 253446 69760
rect 89714 69640 89720 69692
rect 89772 69680 89778 69692
rect 304442 69680 304448 69692
rect 89772 69652 304448 69680
rect 89772 69640 89778 69652
rect 304442 69640 304448 69652
rect 304500 69640 304506 69692
rect 184934 68416 184940 68468
rect 184992 68456 184998 68468
rect 316126 68456 316132 68468
rect 184992 68428 316132 68456
rect 184992 68416 184998 68428
rect 316126 68416 316132 68428
rect 316184 68416 316190 68468
rect 93854 68348 93860 68400
rect 93912 68388 93918 68400
rect 264238 68388 264244 68400
rect 93912 68360 264244 68388
rect 93912 68348 93918 68360
rect 264238 68348 264244 68360
rect 264296 68348 264302 68400
rect 62114 68280 62120 68332
rect 62172 68320 62178 68332
rect 289262 68320 289268 68332
rect 62172 68292 289268 68320
rect 62172 68280 62178 68292
rect 289262 68280 289268 68292
rect 289320 68280 289326 68332
rect 96614 66852 96620 66904
rect 96672 66892 96678 66904
rect 273990 66892 273996 66904
rect 96672 66864 273996 66892
rect 96672 66852 96678 66864
rect 273990 66852 273996 66864
rect 274048 66852 274054 66904
rect 80054 65560 80060 65612
rect 80112 65600 80118 65612
rect 297634 65600 297640 65612
rect 80112 65572 297640 65600
rect 80112 65560 80118 65572
rect 297634 65560 297640 65572
rect 297692 65560 297698 65612
rect 45554 65492 45560 65544
rect 45612 65532 45618 65544
rect 298922 65532 298928 65544
rect 45612 65504 298928 65532
rect 45612 65492 45618 65504
rect 298922 65492 298928 65504
rect 298980 65492 298986 65544
rect 60734 64132 60740 64184
rect 60792 64172 60798 64184
rect 286410 64172 286416 64184
rect 60792 64144 286416 64172
rect 60792 64132 60798 64144
rect 286410 64132 286416 64144
rect 286468 64132 286474 64184
rect 63494 62840 63500 62892
rect 63552 62880 63558 62892
rect 290550 62880 290556 62892
rect 63552 62852 290556 62880
rect 63552 62840 63558 62852
rect 290550 62840 290556 62852
rect 290608 62840 290614 62892
rect 46934 62772 46940 62824
rect 46992 62812 46998 62824
rect 304350 62812 304356 62824
rect 46992 62784 304356 62812
rect 46992 62772 46998 62784
rect 304350 62772 304356 62784
rect 304408 62772 304414 62824
rect 70394 61412 70400 61464
rect 70452 61452 70458 61464
rect 289170 61452 289176 61464
rect 70452 61424 289176 61452
rect 70452 61412 70458 61424
rect 289170 61412 289176 61424
rect 289228 61412 289234 61464
rect 51074 61344 51080 61396
rect 51132 61384 51138 61396
rect 305914 61384 305920 61396
rect 51132 61356 305920 61384
rect 51132 61344 51138 61356
rect 305914 61344 305920 61356
rect 305972 61344 305978 61396
rect 387610 60664 387616 60716
rect 387668 60704 387674 60716
rect 580166 60704 580172 60716
rect 387668 60676 580172 60704
rect 387668 60664 387674 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 53834 59984 53840 60036
rect 53892 60024 53898 60036
rect 296254 60024 296260 60036
rect 53892 59996 296260 60024
rect 53892 59984 53898 59996
rect 296254 59984 296260 59996
rect 296312 59984 296318 60036
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 373258 59344 373264 59356
rect 3108 59316 373264 59344
rect 3108 59304 3114 59316
rect 373258 59304 373264 59316
rect 373316 59304 373322 59356
rect 74534 58624 74540 58676
rect 74592 58664 74598 58676
rect 280982 58664 280988 58676
rect 74592 58636 280988 58664
rect 74592 58624 74598 58636
rect 280982 58624 280988 58636
rect 281040 58624 281046 58676
rect 81434 57264 81440 57316
rect 81492 57304 81498 57316
rect 271322 57304 271328 57316
rect 81492 57276 271328 57304
rect 81492 57264 81498 57276
rect 271322 57264 271328 57276
rect 271380 57264 271386 57316
rect 57974 57196 57980 57248
rect 58032 57236 58038 57248
rect 285122 57236 285128 57248
rect 58032 57208 285128 57236
rect 58032 57196 58038 57208
rect 285122 57196 285128 57208
rect 285180 57196 285186 57248
rect 85574 55904 85580 55956
rect 85632 55944 85638 55956
rect 282178 55944 282184 55956
rect 85632 55916 282184 55944
rect 85632 55904 85638 55916
rect 282178 55904 282184 55916
rect 282236 55904 282242 55956
rect 64874 55836 64880 55888
rect 64932 55876 64938 55888
rect 301682 55876 301688 55888
rect 64932 55848 301688 55876
rect 64932 55836 64938 55848
rect 301682 55836 301688 55848
rect 301740 55836 301746 55888
rect 52546 54476 52552 54528
rect 52604 54516 52610 54528
rect 303154 54516 303160 54528
rect 52604 54488 303160 54516
rect 52604 54476 52610 54488
rect 303154 54476 303160 54488
rect 303212 54476 303218 54528
rect 121454 53116 121460 53168
rect 121512 53156 121518 53168
rect 299014 53156 299020 53168
rect 121512 53128 299020 53156
rect 121512 53116 121518 53128
rect 299014 53116 299020 53128
rect 299072 53116 299078 53168
rect 9674 53048 9680 53100
rect 9732 53088 9738 53100
rect 291930 53088 291936 53100
rect 9732 53060 291936 53088
rect 9732 53048 9738 53060
rect 291930 53048 291936 53060
rect 291988 53048 291994 53100
rect 110414 51756 110420 51808
rect 110472 51796 110478 51808
rect 300210 51796 300216 51808
rect 110472 51768 300216 51796
rect 110472 51756 110478 51768
rect 300210 51756 300216 51768
rect 300268 51756 300274 51808
rect 44174 51688 44180 51740
rect 44232 51728 44238 51740
rect 261570 51728 261576 51740
rect 44232 51700 261576 51728
rect 44232 51688 44238 51700
rect 261570 51688 261576 51700
rect 261628 51688 261634 51740
rect 85666 50396 85672 50448
rect 85724 50436 85730 50448
rect 258810 50436 258816 50448
rect 85724 50408 258816 50436
rect 85724 50396 85730 50408
rect 258810 50396 258816 50408
rect 258868 50396 258874 50448
rect 34514 50328 34520 50380
rect 34572 50368 34578 50380
rect 293310 50368 293316 50380
rect 34572 50340 293316 50368
rect 34572 50328 34578 50340
rect 293310 50328 293316 50340
rect 293368 50328 293374 50380
rect 82814 49036 82820 49088
rect 82872 49076 82878 49088
rect 300302 49076 300308 49088
rect 82872 49048 300308 49076
rect 82872 49036 82878 49048
rect 300302 49036 300308 49048
rect 300360 49036 300366 49088
rect 37274 48968 37280 49020
rect 37332 49008 37338 49020
rect 307110 49008 307116 49020
rect 37332 48980 307116 49008
rect 37332 48968 37338 48980
rect 307110 48968 307116 48980
rect 307168 48968 307174 49020
rect 49602 48220 49608 48272
rect 49660 48260 49666 48272
rect 249242 48260 249248 48272
rect 49660 48232 249248 48260
rect 49660 48220 49666 48232
rect 249242 48220 249248 48232
rect 249300 48220 249306 48272
rect 48958 47880 48964 47932
rect 49016 47920 49022 47932
rect 49602 47920 49608 47932
rect 49016 47892 49608 47920
rect 49016 47880 49022 47892
rect 49602 47880 49608 47892
rect 49660 47880 49666 47932
rect 179598 47540 179604 47592
rect 179656 47580 179662 47592
rect 306374 47580 306380 47592
rect 179656 47552 306380 47580
rect 179656 47540 179662 47552
rect 306374 47540 306380 47552
rect 306432 47540 306438 47592
rect 88334 46180 88340 46232
rect 88392 46220 88398 46232
rect 304258 46220 304264 46232
rect 88392 46192 304264 46220
rect 88392 46180 88398 46192
rect 304258 46180 304264 46192
rect 304316 46180 304322 46232
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 40678 45540 40684 45552
rect 3476 45512 40684 45540
rect 3476 45500 3482 45512
rect 40678 45500 40684 45512
rect 40736 45500 40742 45552
rect 78674 44888 78680 44940
rect 78732 44928 78738 44940
rect 305822 44928 305828 44940
rect 78732 44900 305828 44928
rect 78732 44888 78738 44900
rect 305822 44888 305828 44900
rect 305880 44888 305886 44940
rect 41414 44820 41420 44872
rect 41472 44860 41478 44872
rect 282270 44860 282276 44872
rect 41472 44832 282276 44860
rect 41472 44820 41478 44832
rect 282270 44820 282276 44832
rect 282328 44820 282334 44872
rect 187694 43596 187700 43648
rect 187752 43636 187758 43648
rect 258810 43636 258816 43648
rect 187752 43608 258816 43636
rect 187752 43596 187758 43608
rect 258810 43596 258816 43608
rect 258868 43596 258874 43648
rect 201494 43528 201500 43580
rect 201552 43568 201558 43580
rect 333238 43568 333244 43580
rect 201552 43540 333244 43568
rect 201552 43528 201558 43540
rect 333238 43528 333244 43540
rect 333296 43528 333302 43580
rect 4154 43460 4160 43512
rect 4212 43500 4218 43512
rect 249058 43500 249064 43512
rect 4212 43472 249064 43500
rect 4212 43460 4218 43472
rect 249058 43460 249064 43472
rect 249116 43460 249122 43512
rect 44266 43392 44272 43444
rect 44324 43432 44330 43444
rect 292022 43432 292028 43444
rect 44324 43404 292028 43432
rect 44324 43392 44330 43404
rect 292022 43392 292028 43404
rect 292080 43392 292086 43444
rect 104894 42100 104900 42152
rect 104952 42140 104958 42152
rect 287790 42140 287796 42152
rect 104952 42112 287796 42140
rect 104952 42100 104958 42112
rect 287790 42100 287796 42112
rect 287848 42100 287854 42152
rect 75914 42032 75920 42084
rect 75972 42072 75978 42084
rect 271414 42072 271420 42084
rect 75972 42044 271420 42072
rect 75972 42032 75978 42044
rect 271414 42032 271420 42044
rect 271472 42032 271478 42084
rect 122834 40672 122840 40724
rect 122892 40712 122898 40724
rect 268470 40712 268476 40724
rect 122892 40684 268476 40712
rect 122892 40672 122898 40684
rect 268470 40672 268476 40684
rect 268528 40672 268534 40724
rect 107654 39380 107660 39432
rect 107712 39420 107718 39432
rect 258718 39420 258724 39432
rect 107712 39392 258724 39420
rect 107712 39380 107718 39392
rect 258718 39380 258724 39392
rect 258776 39380 258782 39432
rect 77294 39312 77300 39364
rect 77352 39352 77358 39364
rect 291838 39352 291844 39364
rect 77352 39324 291844 39352
rect 77352 39312 77358 39324
rect 291838 39312 291844 39324
rect 291896 39312 291902 39364
rect 179506 38020 179512 38072
rect 179564 38060 179570 38072
rect 293954 38060 293960 38072
rect 179564 38032 293960 38060
rect 179564 38020 179570 38032
rect 293954 38020 293960 38032
rect 294012 38020 294018 38072
rect 93946 37952 93952 38004
rect 94004 37992 94010 38004
rect 266998 37992 267004 38004
rect 94004 37964 267004 37992
rect 94004 37952 94010 37964
rect 266998 37952 267004 37964
rect 267056 37952 267062 38004
rect 42794 37884 42800 37936
rect 42852 37924 42858 37936
rect 286318 37924 286324 37936
rect 42852 37896 286324 37924
rect 42852 37884 42858 37896
rect 286318 37884 286324 37896
rect 286376 37884 286382 37936
rect 16574 36524 16580 36576
rect 16632 36564 16638 36576
rect 297542 36564 297548 36576
rect 16632 36536 297548 36564
rect 16632 36524 16638 36536
rect 297542 36524 297548 36536
rect 297600 36524 297606 36576
rect 177942 35300 177948 35352
rect 178000 35340 178006 35352
rect 298922 35340 298928 35352
rect 178000 35312 298928 35340
rect 178000 35300 178006 35312
rect 298922 35300 298928 35312
rect 298980 35300 298986 35352
rect 27706 35232 27712 35284
rect 27764 35272 27770 35284
rect 272518 35272 272524 35284
rect 27764 35244 272524 35272
rect 27764 35232 27770 35244
rect 272518 35232 272524 35244
rect 272576 35232 272582 35284
rect 20714 35164 20720 35216
rect 20772 35204 20778 35216
rect 305730 35204 305736 35216
rect 20772 35176 305736 35204
rect 20772 35164 20778 35176
rect 305730 35164 305736 35176
rect 305788 35164 305794 35216
rect 179414 33872 179420 33924
rect 179472 33912 179478 33924
rect 332686 33912 332692 33924
rect 179472 33884 332692 33912
rect 179472 33872 179478 33884
rect 332686 33872 332692 33884
rect 332744 33872 332750 33924
rect 71774 33804 71780 33856
rect 71832 33844 71838 33856
rect 256050 33844 256056 33856
rect 71832 33816 256056 33844
rect 71832 33804 71838 33816
rect 256050 33804 256056 33816
rect 256108 33804 256114 33856
rect 97994 33736 98000 33788
rect 98052 33776 98058 33788
rect 294598 33776 294604 33788
rect 98052 33748 294604 33776
rect 98052 33736 98058 33748
rect 294598 33736 294604 33748
rect 294656 33736 294662 33788
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 13078 33096 13084 33108
rect 3568 33068 13084 33096
rect 3568 33056 3574 33068
rect 13078 33056 13084 33068
rect 13136 33056 13142 33108
rect 522298 33056 522304 33108
rect 522356 33096 522362 33108
rect 580166 33096 580172 33108
rect 522356 33068 580172 33096
rect 522356 33056 522362 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 208394 32512 208400 32564
rect 208452 32552 208458 32564
rect 323578 32552 323584 32564
rect 208452 32524 323584 32552
rect 208452 32512 208458 32524
rect 323578 32512 323584 32524
rect 323636 32512 323642 32564
rect 106274 32444 106280 32496
rect 106332 32484 106338 32496
rect 250438 32484 250444 32496
rect 106332 32456 250444 32484
rect 106332 32444 106338 32456
rect 250438 32444 250444 32456
rect 250496 32444 250502 32496
rect 48314 32376 48320 32428
rect 48372 32416 48378 32428
rect 298738 32416 298744 32428
rect 48372 32388 298744 32416
rect 48372 32376 48378 32388
rect 298738 32376 298744 32388
rect 298796 32376 298802 32428
rect 73154 31084 73160 31136
rect 73212 31124 73218 31136
rect 302970 31124 302976 31136
rect 73212 31096 302976 31124
rect 73212 31084 73218 31096
rect 302970 31084 302976 31096
rect 303028 31084 303034 31136
rect 33134 31016 33140 31068
rect 33192 31056 33198 31068
rect 287882 31056 287888 31068
rect 33192 31028 287888 31056
rect 33192 31016 33198 31028
rect 287882 31016 287888 31028
rect 287940 31016 287946 31068
rect 176562 29724 176568 29776
rect 176620 29764 176626 29776
rect 262214 29764 262220 29776
rect 176620 29736 262220 29764
rect 176620 29724 176626 29736
rect 262214 29724 262220 29736
rect 262272 29724 262278 29776
rect 118694 29656 118700 29708
rect 118752 29696 118758 29708
rect 228358 29696 228364 29708
rect 118752 29668 228364 29696
rect 118752 29656 118758 29668
rect 228358 29656 228364 29668
rect 228416 29656 228422 29708
rect 12434 29588 12440 29640
rect 12492 29628 12498 29640
rect 289078 29628 289084 29640
rect 12492 29600 289084 29628
rect 12492 29588 12498 29600
rect 289078 29588 289084 29600
rect 289136 29588 289142 29640
rect 102134 28296 102140 28348
rect 102192 28336 102198 28348
rect 293218 28336 293224 28348
rect 102192 28308 293224 28336
rect 102192 28296 102198 28308
rect 293218 28296 293224 28308
rect 293276 28296 293282 28348
rect 26234 28228 26240 28280
rect 26292 28268 26298 28280
rect 275370 28268 275376 28280
rect 26292 28240 275376 28268
rect 26292 28228 26298 28240
rect 275370 28228 275376 28240
rect 275428 28228 275434 28280
rect 100754 26868 100760 26920
rect 100812 26908 100818 26920
rect 301590 26908 301596 26920
rect 100812 26880 301596 26908
rect 100812 26868 100818 26880
rect 301590 26868 301596 26880
rect 301648 26868 301654 26920
rect 91094 25576 91100 25628
rect 91152 25616 91158 25628
rect 283742 25616 283748 25628
rect 91152 25588 283748 25616
rect 91152 25576 91158 25588
rect 283742 25576 283748 25588
rect 283800 25576 283806 25628
rect 24854 25508 24860 25560
rect 24912 25548 24918 25560
rect 298830 25548 298836 25560
rect 24912 25520 298836 25548
rect 24912 25508 24918 25520
rect 298830 25508 298836 25520
rect 298888 25508 298894 25560
rect 193214 24216 193220 24268
rect 193272 24256 193278 24268
rect 242158 24256 242164 24268
rect 193272 24228 242164 24256
rect 193272 24216 193278 24228
rect 242158 24216 242164 24228
rect 242216 24216 242222 24268
rect 56594 24148 56600 24200
rect 56652 24188 56658 24200
rect 262858 24188 262864 24200
rect 56652 24160 262864 24188
rect 56652 24148 56658 24160
rect 262858 24148 262864 24160
rect 262916 24148 262922 24200
rect 2866 24080 2872 24132
rect 2924 24120 2930 24132
rect 275278 24120 275284 24132
rect 2924 24092 275284 24120
rect 2924 24080 2930 24092
rect 275278 24080 275284 24092
rect 275336 24080 275342 24132
rect 86954 22788 86960 22840
rect 87012 22828 87018 22840
rect 290458 22828 290464 22840
rect 87012 22800 290464 22828
rect 87012 22788 87018 22800
rect 290458 22788 290464 22800
rect 290516 22788 290522 22840
rect 19334 22720 19340 22772
rect 19392 22760 19398 22772
rect 255958 22760 255964 22772
rect 19392 22732 255964 22760
rect 19392 22720 19398 22732
rect 255958 22720 255964 22732
rect 256016 22720 256022 22772
rect 179230 21496 179236 21548
rect 179288 21536 179294 21548
rect 284294 21536 284300 21548
rect 179288 21508 284300 21536
rect 179288 21496 179294 21508
rect 284294 21496 284300 21508
rect 284352 21496 284358 21548
rect 40034 21428 40040 21480
rect 40092 21468 40098 21480
rect 269850 21468 269856 21480
rect 40092 21440 269856 21468
rect 40092 21428 40098 21440
rect 269850 21428 269856 21440
rect 269908 21428 269914 21480
rect 15194 21360 15200 21412
rect 15252 21400 15258 21412
rect 307018 21400 307024 21412
rect 15252 21372 307024 21400
rect 15252 21360 15258 21372
rect 307018 21360 307024 21372
rect 307076 21360 307082 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 22830 20652 22836 20664
rect 3476 20624 22836 20652
rect 3476 20612 3482 20624
rect 22830 20612 22836 20624
rect 22888 20612 22894 20664
rect 195238 20068 195244 20120
rect 195296 20108 195302 20120
rect 273254 20108 273260 20120
rect 195296 20080 273260 20108
rect 195296 20068 195302 20080
rect 273254 20068 273260 20080
rect 273312 20068 273318 20120
rect 115934 20000 115940 20052
rect 115992 20040 115998 20052
rect 296070 20040 296076 20052
rect 115992 20012 296076 20040
rect 115992 20000 115998 20012
rect 296070 20000 296076 20012
rect 296128 20000 296134 20052
rect 38654 19932 38660 19984
rect 38712 19972 38718 19984
rect 278130 19972 278136 19984
rect 38712 19944 278136 19972
rect 38712 19932 38718 19944
rect 278130 19932 278136 19944
rect 278188 19932 278194 19984
rect 109034 18640 109040 18692
rect 109092 18680 109098 18692
rect 278222 18680 278228 18692
rect 109092 18652 278228 18680
rect 109092 18640 109098 18652
rect 278222 18640 278228 18652
rect 278280 18640 278286 18692
rect 11146 18572 11152 18624
rect 11204 18612 11210 18624
rect 253290 18612 253296 18624
rect 11204 18584 253296 18612
rect 11204 18572 11210 18584
rect 253290 18572 253296 18584
rect 253348 18572 253354 18624
rect 110506 17280 110512 17332
rect 110564 17320 110570 17332
rect 279418 17320 279424 17332
rect 110564 17292 279424 17320
rect 110564 17280 110570 17292
rect 279418 17280 279424 17292
rect 279476 17280 279482 17332
rect 23474 17212 23480 17264
rect 23532 17252 23538 17264
rect 280798 17252 280804 17264
rect 23532 17224 280804 17252
rect 23532 17212 23538 17224
rect 280798 17212 280804 17224
rect 280856 17212 280862 17264
rect 175182 15920 175188 15972
rect 175240 15960 175246 15972
rect 311434 15960 311440 15972
rect 175240 15932 311440 15960
rect 175240 15920 175246 15932
rect 311434 15920 311440 15932
rect 311492 15920 311498 15972
rect 84194 15852 84200 15904
rect 84252 15892 84258 15904
rect 262950 15892 262956 15904
rect 84252 15864 262956 15892
rect 84252 15852 84258 15864
rect 262950 15852 262956 15864
rect 263008 15852 263014 15904
rect 135254 14492 135260 14544
rect 135312 14532 135318 14544
rect 203518 14532 203524 14544
rect 135312 14504 203524 14532
rect 135312 14492 135318 14504
rect 203518 14492 203524 14504
rect 203576 14492 203582 14544
rect 233878 14492 233884 14544
rect 233936 14532 233942 14544
rect 281534 14532 281540 14544
rect 233936 14504 281540 14532
rect 233936 14492 233942 14504
rect 281534 14492 281540 14504
rect 281592 14492 281598 14544
rect 36722 14424 36728 14476
rect 36780 14464 36786 14476
rect 303062 14464 303068 14476
rect 36780 14436 303068 14464
rect 36780 14424 36786 14436
rect 303062 14424 303068 14436
rect 303120 14424 303126 14476
rect 183554 13200 183560 13252
rect 183612 13240 183618 13252
rect 349246 13240 349252 13252
rect 183612 13212 349252 13240
rect 183612 13200 183618 13212
rect 349246 13200 349252 13212
rect 349304 13200 349310 13252
rect 22554 13132 22560 13184
rect 22612 13172 22618 13184
rect 254578 13172 254584 13184
rect 22612 13144 254584 13172
rect 22612 13132 22618 13144
rect 254578 13132 254584 13144
rect 254636 13132 254642 13184
rect 59354 13064 59360 13116
rect 59412 13104 59418 13116
rect 300118 13104 300124 13116
rect 59412 13076 300124 13104
rect 59412 13064 59418 13076
rect 300118 13064 300124 13076
rect 300176 13064 300182 13116
rect 128906 11840 128912 11892
rect 128964 11880 128970 11892
rect 216674 11880 216680 11892
rect 128964 11852 216680 11880
rect 128964 11840 128970 11852
rect 216674 11840 216680 11852
rect 216732 11840 216738 11892
rect 112346 11772 112352 11824
rect 112404 11812 112410 11824
rect 305638 11812 305644 11824
rect 112404 11784 305644 11812
rect 112404 11772 112410 11784
rect 305638 11772 305644 11784
rect 305696 11772 305702 11824
rect 30098 11704 30104 11756
rect 30156 11744 30162 11756
rect 271230 11744 271236 11756
rect 30156 11716 271236 11744
rect 30156 11704 30162 11716
rect 271230 11704 271236 11716
rect 271288 11704 271294 11756
rect 106 10956 112 11008
rect 164 10996 170 11008
rect 1302 10996 1308 11008
rect 164 10968 1308 10996
rect 164 10956 170 10968
rect 1302 10956 1308 10968
rect 1360 10996 1366 11008
rect 251174 10996 251180 11008
rect 1360 10968 251180 10996
rect 1360 10956 1366 10968
rect 251174 10956 251180 10968
rect 251232 10956 251238 11008
rect 176470 10344 176476 10396
rect 176528 10384 176534 10396
rect 299474 10384 299480 10396
rect 176528 10356 299480 10384
rect 176528 10344 176534 10356
rect 299474 10344 299480 10356
rect 299532 10344 299538 10396
rect 92474 10276 92480 10328
rect 92532 10316 92538 10328
rect 283558 10316 283564 10328
rect 92532 10288 283564 10316
rect 92532 10276 92538 10288
rect 283558 10276 283564 10288
rect 283616 10276 283622 10328
rect 189718 9052 189724 9104
rect 189776 9092 189782 9104
rect 245194 9092 245200 9104
rect 189776 9064 245200 9092
rect 189776 9052 189782 9064
rect 245194 9052 245200 9064
rect 245252 9052 245258 9104
rect 96246 8984 96252 9036
rect 96304 9024 96310 9036
rect 285030 9024 285036 9036
rect 96304 8996 285036 9024
rect 96304 8984 96310 8996
rect 285030 8984 285036 8996
rect 285088 8984 285094 9036
rect 1670 8916 1676 8968
rect 1728 8956 1734 8968
rect 48958 8956 48964 8968
rect 1728 8928 48964 8956
rect 1728 8916 1734 8928
rect 48958 8916 48964 8928
rect 49016 8916 49022 8968
rect 62022 8916 62028 8968
rect 62080 8956 62086 8968
rect 283650 8956 283656 8968
rect 62080 8928 283656 8956
rect 62080 8916 62086 8928
rect 283650 8916 283656 8928
rect 283708 8916 283714 8968
rect 99834 7624 99840 7676
rect 99892 7664 99898 7676
rect 273898 7664 273904 7676
rect 99892 7636 273904 7664
rect 99892 7624 99898 7636
rect 273898 7624 273904 7636
rect 273956 7624 273962 7676
rect 7650 7556 7656 7608
rect 7708 7596 7714 7608
rect 301498 7596 301504 7608
rect 7708 7568 301504 7596
rect 7708 7556 7714 7568
rect 301498 7556 301504 7568
rect 301556 7556 301562 7608
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 35158 6848 35164 6860
rect 3476 6820 35164 6848
rect 3476 6808 3482 6820
rect 35158 6808 35164 6820
rect 35216 6808 35222 6860
rect 180794 6332 180800 6384
rect 180852 6372 180858 6384
rect 268838 6372 268844 6384
rect 180852 6344 268844 6372
rect 180852 6332 180858 6344
rect 268838 6332 268844 6344
rect 268896 6332 268902 6384
rect 211798 6264 211804 6316
rect 211856 6304 211862 6316
rect 305546 6304 305552 6316
rect 211856 6276 305552 6304
rect 211856 6264 211862 6276
rect 305546 6264 305552 6276
rect 305604 6264 305610 6316
rect 309042 6264 309048 6316
rect 309100 6304 309106 6316
rect 335446 6304 335452 6316
rect 309100 6276 335452 6304
rect 309100 6264 309106 6276
rect 335446 6264 335452 6276
rect 335504 6264 335510 6316
rect 182818 6196 182824 6248
rect 182876 6236 182882 6248
rect 348050 6236 348056 6248
rect 182876 6208 348056 6236
rect 182876 6196 182882 6208
rect 348050 6196 348056 6208
rect 348108 6196 348114 6248
rect 70302 6128 70308 6180
rect 70360 6168 70366 6180
rect 287698 6168 287704 6180
rect 70360 6140 287704 6168
rect 70360 6128 70366 6140
rect 287698 6128 287704 6140
rect 287756 6128 287762 6180
rect 303154 6128 303160 6180
rect 303212 6168 303218 6180
rect 332594 6168 332600 6180
rect 303212 6140 332600 6168
rect 303212 6128 303218 6140
rect 332594 6128 332600 6140
rect 332652 6128 332658 6180
rect 197998 4836 198004 4888
rect 198056 4876 198062 4888
rect 260650 4876 260656 4888
rect 198056 4848 260656 4876
rect 198056 4836 198062 4848
rect 260650 4836 260656 4848
rect 260708 4836 260714 4888
rect 35986 4768 35992 4820
rect 36044 4808 36050 4820
rect 265618 4808 265624 4820
rect 36044 4780 265624 4808
rect 36044 4768 36050 4780
rect 265618 4768 265624 4780
rect 265676 4768 265682 4820
rect 216122 3680 216128 3732
rect 216180 3720 216186 3732
rect 240502 3720 240508 3732
rect 216180 3692 240508 3720
rect 216180 3680 216186 3692
rect 240502 3680 240508 3692
rect 240560 3680 240566 3732
rect 242158 3680 242164 3732
rect 242216 3720 242222 3732
rect 247586 3720 247592 3732
rect 242216 3692 247592 3720
rect 242216 3680 242222 3692
rect 247586 3680 247592 3692
rect 247644 3680 247650 3732
rect 253474 3680 253480 3732
rect 253532 3720 253538 3732
rect 261478 3720 261484 3732
rect 253532 3692 261484 3720
rect 253532 3680 253538 3692
rect 261478 3680 261484 3692
rect 261536 3680 261542 3732
rect 114002 3612 114008 3664
rect 114060 3652 114066 3664
rect 114060 3624 122834 3652
rect 114060 3612 114066 3624
rect 110414 3544 110420 3596
rect 110472 3584 110478 3596
rect 111610 3584 111616 3596
rect 110472 3556 111616 3584
rect 110472 3544 110478 3556
rect 111610 3544 111616 3556
rect 111668 3544 111674 3596
rect 118694 3544 118700 3596
rect 118752 3584 118758 3596
rect 119890 3584 119896 3596
rect 118752 3556 119896 3584
rect 118752 3544 118758 3556
rect 119890 3544 119896 3556
rect 119948 3544 119954 3596
rect 122806 3584 122834 3624
rect 211062 3612 211068 3664
rect 211120 3652 211126 3664
rect 248782 3652 248788 3664
rect 211120 3624 248788 3652
rect 211120 3612 211126 3624
rect 248782 3612 248788 3624
rect 248840 3612 248846 3664
rect 254670 3652 254676 3664
rect 251008 3624 254676 3652
rect 210418 3584 210424 3596
rect 122806 3556 210424 3584
rect 210418 3544 210424 3556
rect 210476 3544 210482 3596
rect 216030 3544 216036 3596
rect 216088 3584 216094 3596
rect 251008 3584 251036 3624
rect 254670 3612 254676 3624
rect 254728 3612 254734 3664
rect 268378 3612 268384 3664
rect 268436 3652 268442 3664
rect 268436 3624 277394 3652
rect 268436 3612 268442 3624
rect 216088 3556 251036 3584
rect 216088 3544 216094 3556
rect 251082 3544 251088 3596
rect 251140 3584 251146 3596
rect 252370 3584 252376 3596
rect 251140 3556 252376 3584
rect 251140 3544 251146 3556
rect 252370 3544 252376 3556
rect 252428 3544 252434 3596
rect 257982 3544 257988 3596
rect 258040 3584 258046 3596
rect 264146 3584 264152 3596
rect 258040 3556 264152 3584
rect 258040 3544 258046 3556
rect 264146 3544 264152 3556
rect 264204 3544 264210 3596
rect 276014 3544 276020 3596
rect 276072 3584 276078 3596
rect 276750 3584 276756 3596
rect 276072 3556 276756 3584
rect 276072 3544 276078 3556
rect 276750 3544 276756 3556
rect 276808 3544 276814 3596
rect 277366 3584 277394 3624
rect 284938 3612 284944 3664
rect 284996 3652 285002 3664
rect 298462 3652 298468 3664
rect 284996 3624 298468 3652
rect 284996 3612 285002 3624
rect 298462 3612 298468 3624
rect 298520 3612 298526 3664
rect 288986 3584 288992 3596
rect 277366 3556 288992 3584
rect 288986 3544 288992 3556
rect 289044 3544 289050 3596
rect 299566 3544 299572 3596
rect 299624 3584 299630 3596
rect 300762 3584 300768 3596
rect 299624 3556 300768 3584
rect 299624 3544 299630 3556
rect 300762 3544 300768 3556
rect 300820 3544 300826 3596
rect 319714 3544 319720 3596
rect 319772 3584 319778 3596
rect 331214 3584 331220 3596
rect 319772 3556 331220 3584
rect 319772 3544 319778 3556
rect 331214 3544 331220 3556
rect 331272 3544 331278 3596
rect 331858 3544 331864 3596
rect 331916 3584 331922 3596
rect 333882 3584 333888 3596
rect 331916 3556 333888 3584
rect 331916 3544 331922 3556
rect 333882 3544 333888 3556
rect 333940 3544 333946 3596
rect 11054 3476 11060 3528
rect 11112 3516 11118 3528
rect 11974 3516 11980 3528
rect 11112 3488 11980 3516
rect 11112 3476 11118 3488
rect 11974 3476 11980 3488
rect 12032 3476 12038 3528
rect 27614 3476 27620 3528
rect 27672 3516 27678 3528
rect 28534 3516 28540 3528
rect 27672 3488 28540 3516
rect 27672 3476 27678 3488
rect 28534 3476 28540 3488
rect 28592 3476 28598 3528
rect 44174 3476 44180 3528
rect 44232 3516 44238 3528
rect 45094 3516 45100 3528
rect 44232 3488 45100 3516
rect 44232 3476 44238 3488
rect 45094 3476 45100 3488
rect 45152 3476 45158 3528
rect 103330 3476 103336 3528
rect 103388 3516 103394 3528
rect 211890 3516 211896 3528
rect 103388 3488 211896 3516
rect 103388 3476 103394 3488
rect 211890 3476 211896 3488
rect 211948 3476 211954 3528
rect 215938 3476 215944 3528
rect 215996 3516 216002 3528
rect 215996 3488 258672 3516
rect 215996 3476 216002 3488
rect 6454 3408 6460 3460
rect 6512 3448 6518 3460
rect 192478 3448 192484 3460
rect 6512 3420 192484 3448
rect 6512 3408 6518 3420
rect 192478 3408 192484 3420
rect 192536 3408 192542 3460
rect 196618 3408 196624 3460
rect 196676 3448 196682 3460
rect 196676 3420 258074 3448
rect 196676 3408 196682 3420
rect 135254 3340 135260 3392
rect 135312 3380 135318 3392
rect 136450 3380 136456 3392
rect 135312 3352 136456 3380
rect 135312 3340 135318 3352
rect 136450 3340 136456 3352
rect 136508 3340 136514 3392
rect 235810 3340 235816 3392
rect 235868 3380 235874 3392
rect 238018 3380 238024 3392
rect 235868 3352 238024 3380
rect 235868 3340 235874 3352
rect 238018 3340 238024 3352
rect 238076 3340 238082 3392
rect 242894 3340 242900 3392
rect 242952 3380 242958 3392
rect 244090 3380 244096 3392
rect 242952 3352 244096 3380
rect 242952 3340 242958 3352
rect 244090 3340 244096 3352
rect 244148 3340 244154 3392
rect 249978 3340 249984 3392
rect 250036 3380 250042 3392
rect 253198 3380 253204 3392
rect 250036 3352 253204 3380
rect 250036 3340 250042 3352
rect 253198 3340 253204 3352
rect 253256 3340 253262 3392
rect 241698 3272 241704 3324
rect 241756 3312 241762 3324
rect 246298 3312 246304 3324
rect 241756 3284 246304 3312
rect 241756 3272 241762 3284
rect 246298 3272 246304 3284
rect 246356 3272 246362 3324
rect 258046 3312 258074 3420
rect 258644 3380 258672 3488
rect 258810 3476 258816 3528
rect 258868 3516 258874 3528
rect 261754 3516 261760 3528
rect 258868 3488 261760 3516
rect 258868 3476 258874 3488
rect 261754 3476 261760 3488
rect 261812 3476 261818 3528
rect 271138 3476 271144 3528
rect 271196 3516 271202 3528
rect 326798 3516 326804 3528
rect 271196 3488 326804 3516
rect 271196 3476 271202 3488
rect 326798 3476 326804 3488
rect 326856 3476 326862 3528
rect 329098 3476 329104 3528
rect 329156 3516 329162 3528
rect 330386 3516 330392 3528
rect 329156 3488 330392 3516
rect 329156 3476 329162 3488
rect 330386 3476 330392 3488
rect 330444 3476 330450 3528
rect 333238 3476 333244 3528
rect 333296 3516 333302 3528
rect 344554 3516 344560 3528
rect 333296 3488 344560 3516
rect 333296 3476 333302 3488
rect 344554 3476 344560 3488
rect 344612 3476 344618 3528
rect 349154 3476 349160 3528
rect 349212 3516 349218 3528
rect 350442 3516 350448 3528
rect 349212 3488 350448 3516
rect 349212 3476 349218 3488
rect 350442 3476 350448 3488
rect 350500 3476 350506 3528
rect 292574 3448 292580 3460
rect 267706 3420 292580 3448
rect 266538 3380 266544 3392
rect 258644 3352 266544 3380
rect 266538 3340 266544 3352
rect 266596 3340 266602 3392
rect 267706 3312 267734 3420
rect 292574 3408 292580 3420
rect 292632 3408 292638 3460
rect 298922 3408 298928 3460
rect 298980 3448 298986 3460
rect 301958 3448 301964 3460
rect 298980 3420 301964 3448
rect 298980 3408 298986 3420
rect 301958 3408 301964 3420
rect 302016 3408 302022 3460
rect 322106 3448 322112 3460
rect 306346 3420 322112 3448
rect 297358 3340 297364 3392
rect 297416 3380 297422 3392
rect 306346 3380 306374 3420
rect 322106 3408 322112 3420
rect 322164 3408 322170 3460
rect 323302 3408 323308 3460
rect 323360 3448 323366 3460
rect 340874 3448 340880 3460
rect 323360 3420 340880 3448
rect 323360 3408 323366 3420
rect 340874 3408 340880 3420
rect 340932 3408 340938 3460
rect 342162 3408 342168 3460
rect 342220 3448 342226 3460
rect 343634 3448 343640 3460
rect 342220 3420 343640 3448
rect 342220 3408 342226 3420
rect 343634 3408 343640 3420
rect 343692 3408 343698 3460
rect 297416 3352 306374 3380
rect 297416 3340 297422 3352
rect 309778 3340 309784 3392
rect 309836 3380 309842 3392
rect 317322 3380 317328 3392
rect 309836 3352 317328 3380
rect 309836 3340 309842 3352
rect 317322 3340 317328 3352
rect 317380 3340 317386 3392
rect 323578 3340 323584 3392
rect 323636 3380 323642 3392
rect 325602 3380 325608 3392
rect 323636 3352 325608 3380
rect 323636 3340 323642 3352
rect 325602 3340 325608 3352
rect 325660 3340 325666 3392
rect 258046 3284 267734 3312
rect 309870 3272 309876 3324
rect 309928 3312 309934 3324
rect 315022 3312 315028 3324
rect 309928 3284 315028 3312
rect 309928 3272 309934 3284
rect 315022 3272 315028 3284
rect 315080 3272 315086 3324
rect 258258 3000 258264 3052
rect 258316 3040 258322 3052
rect 260098 3040 260104 3052
rect 258316 3012 260104 3040
rect 258316 3000 258322 3012
rect 260098 3000 260104 3012
rect 260156 3000 260162 3052
rect 308490 2932 308496 2984
rect 308548 2972 308554 2984
rect 310238 2972 310244 2984
rect 308548 2944 310244 2972
rect 308548 2932 308554 2944
rect 310238 2932 310244 2944
rect 310296 2932 310302 2984
rect 346946 2932 346952 2984
rect 347004 2972 347010 2984
rect 351914 2972 351920 2984
rect 347004 2944 351920 2972
rect 347004 2932 347010 2944
rect 351914 2932 351920 2944
rect 351972 2932 351978 2984
rect 278038 2864 278044 2916
rect 278096 2904 278102 2916
rect 283098 2904 283104 2916
rect 278096 2876 283104 2904
rect 278096 2864 278102 2876
rect 283098 2864 283104 2876
rect 283156 2864 283162 2916
rect 118786 2116 118792 2168
rect 118844 2156 118850 2168
rect 295978 2156 295984 2168
rect 118844 2128 295984 2156
rect 118844 2116 118850 2128
rect 295978 2116 295984 2128
rect 296036 2116 296042 2168
rect 19426 2048 19432 2100
rect 19484 2088 19490 2100
rect 269758 2088 269764 2100
rect 19484 2060 269764 2088
rect 19484 2048 19490 2060
rect 269758 2048 269764 2060
rect 269816 2048 269822 2100
<< via1 >>
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 206284 702448 206336 702500
rect 559656 702448 559708 702500
rect 300124 700408 300176 700460
rect 310520 700408 310572 700460
rect 149704 700340 149756 700392
rect 170312 700340 170364 700392
rect 218980 700340 219032 700392
rect 309140 700340 309192 700392
rect 354588 700340 354640 700392
rect 364984 700340 365036 700392
rect 383568 700340 383620 700392
rect 478512 700340 478564 700392
rect 559656 700340 559708 700392
rect 582380 700340 582432 700392
rect 72976 700272 73028 700324
rect 94504 700272 94556 700324
rect 105452 700272 105504 700324
rect 193220 700272 193272 700324
rect 235172 700272 235224 700324
rect 299480 700272 299532 700324
rect 302056 700272 302108 700324
rect 429844 700272 429896 700324
rect 527180 700272 527232 700324
rect 565820 700272 565872 700324
rect 24308 699660 24360 699712
rect 25504 699660 25556 699712
rect 307668 698912 307720 698964
rect 397460 698912 397512 698964
rect 179052 697552 179104 697604
rect 267648 697552 267700 697604
rect 212448 696192 212500 696244
rect 348792 696192 348844 696244
rect 3424 684156 3476 684208
rect 8944 684156 8996 684208
rect 567844 683136 567896 683188
rect 580172 683136 580224 683188
rect 3516 670692 3568 670744
rect 66904 670692 66956 670744
rect 6920 669944 6972 669996
rect 62764 669944 62816 669996
rect 3424 656888 3476 656940
rect 32404 656888 32456 656940
rect 574744 643084 574796 643136
rect 580172 643084 580224 643136
rect 3424 632068 3476 632120
rect 44824 632068 44876 632120
rect 502984 630640 503036 630692
rect 580172 630640 580224 630692
rect 3148 618264 3200 618316
rect 22744 618264 22796 618316
rect 3240 605820 3292 605872
rect 90364 605820 90416 605872
rect 530584 590656 530636 590708
rect 579804 590656 579856 590708
rect 391204 576852 391256 576904
rect 580172 576852 580224 576904
rect 3424 565836 3476 565888
rect 57244 565836 57296 565888
rect 3424 553392 3476 553444
rect 36544 553392 36596 553444
rect 576124 536800 576176 536852
rect 580172 536800 580224 536852
rect 3424 527144 3476 527196
rect 39304 527144 39356 527196
rect 3424 514768 3476 514820
rect 48964 514768 49016 514820
rect 3056 500964 3108 501016
rect 120724 500964 120776 501016
rect 536104 484372 536156 484424
rect 580172 484372 580224 484424
rect 3424 474716 3476 474768
rect 31024 474716 31076 474768
rect 274548 470568 274600 470620
rect 580172 470568 580224 470620
rect 3240 462340 3292 462392
rect 98644 462340 98696 462392
rect 573364 458804 573416 458856
rect 580264 458804 580316 458856
rect 3148 448536 3200 448588
rect 53104 448536 53156 448588
rect 392584 430584 392636 430636
rect 580172 430584 580224 430636
rect 3424 422288 3476 422340
rect 13084 422288 13136 422340
rect 577504 418140 577556 418192
rect 579620 418140 579672 418192
rect 3148 409844 3200 409896
rect 50344 409844 50396 409896
rect 388444 404336 388496 404388
rect 580172 404336 580224 404388
rect 3424 397468 3476 397520
rect 58624 397468 58676 397520
rect 48964 381488 49016 381540
rect 247040 381488 247092 381540
rect 153200 380128 153252 380180
rect 270500 380128 270552 380180
rect 55036 378768 55088 378820
rect 138020 378768 138072 378820
rect 295340 378768 295392 378820
rect 574100 377408 574152 377460
rect 580172 377408 580224 377460
rect 209044 376728 209096 376780
rect 574100 376728 574152 376780
rect 195244 374620 195296 374672
rect 331220 374620 331272 374672
rect 53104 372580 53156 372632
rect 53748 372580 53800 372632
rect 291844 372580 291896 372632
rect 98644 371832 98696 371884
rect 125600 371832 125652 371884
rect 126612 371832 126664 371884
rect 232504 371288 232556 371340
rect 313924 371288 313976 371340
rect 3424 371220 3476 371272
rect 111064 371220 111116 371272
rect 126612 371220 126664 371272
rect 267004 371220 267056 371272
rect 8944 370472 8996 370524
rect 144092 370472 144144 370524
rect 143540 369860 143592 369912
rect 144092 369860 144144 369912
rect 198740 369860 198792 369912
rect 211804 369860 211856 369912
rect 212448 369860 212500 369912
rect 583024 369860 583076 369912
rect 31024 369112 31076 369164
rect 146944 369112 146996 369164
rect 146944 368636 146996 368688
rect 202880 368636 202932 368688
rect 140044 368568 140096 368620
rect 282920 368568 282972 368620
rect 170956 368500 171008 368552
rect 578240 368500 578292 368552
rect 578884 368500 578936 368552
rect 39304 368432 39356 368484
rect 39948 368432 40000 368484
rect 282920 367752 282972 367804
rect 293960 367752 294012 367804
rect 226340 367276 226392 367328
rect 340880 367276 340932 367328
rect 114560 367208 114612 367260
rect 295984 367208 296036 367260
rect 39948 367140 40000 367192
rect 264244 367140 264296 367192
rect 175096 367072 175148 367124
rect 561956 367072 562008 367124
rect 171784 366392 171836 366444
rect 201500 366392 201552 366444
rect 32404 366324 32456 366376
rect 234620 366324 234672 366376
rect 189080 365780 189132 365832
rect 307024 365780 307076 365832
rect 219440 365712 219492 365764
rect 571432 365712 571484 365764
rect 208400 365644 208452 365696
rect 209044 365644 209096 365696
rect 238760 364556 238812 364608
rect 302240 364556 302292 364608
rect 162308 364488 162360 364540
rect 208400 364488 208452 364540
rect 251180 364488 251232 364540
rect 331220 364488 331272 364540
rect 129004 364420 129056 364472
rect 282920 364420 282972 364472
rect 120724 364352 120776 364404
rect 296904 364352 296956 364404
rect 570512 364352 570564 364404
rect 580172 364352 580224 364404
rect 228824 363128 228876 363180
rect 318064 363128 318116 363180
rect 166264 363060 166316 363112
rect 287428 363060 287480 363112
rect 130384 362992 130436 363044
rect 298284 362992 298336 363044
rect 178684 362924 178736 362976
rect 580356 362924 580408 362976
rect 138664 361904 138716 361956
rect 193220 361904 193272 361956
rect 134524 361836 134576 361888
rect 231676 361836 231728 361888
rect 315304 361836 315356 361888
rect 181628 361768 181680 361820
rect 319444 361768 319496 361820
rect 111156 361700 111208 361752
rect 299572 361700 299624 361752
rect 179512 361632 179564 361684
rect 463424 361632 463476 361684
rect 64788 361564 64840 361616
rect 195244 361564 195296 361616
rect 243636 361564 243688 361616
rect 563704 361564 563756 361616
rect 126244 360612 126296 360664
rect 279332 360612 279384 360664
rect 280068 360612 280120 360664
rect 250536 360544 250588 360596
rect 297364 360544 297416 360596
rect 176108 360476 176160 360528
rect 237472 360476 237524 360528
rect 329196 360476 329248 360528
rect 176016 360408 176068 360460
rect 219440 360408 219492 360460
rect 220268 360408 220320 360460
rect 233792 360408 233844 360460
rect 332600 360408 332652 360460
rect 113180 360340 113232 360392
rect 296812 360340 296864 360392
rect 275008 360272 275060 360324
rect 538864 360272 538916 360324
rect 79324 360204 79376 360256
rect 245844 360204 245896 360256
rect 280068 360204 280120 360256
rect 578332 360204 578384 360256
rect 172428 359116 172480 359168
rect 218336 359116 218388 359168
rect 173164 359048 173216 359100
rect 296720 359048 296772 359100
rect 142804 358980 142856 359032
rect 201592 358980 201644 359032
rect 234620 358980 234672 359032
rect 235540 358980 235592 359032
rect 374644 358980 374696 359032
rect 109040 358912 109092 358964
rect 253940 358912 253992 358964
rect 264244 358912 264296 358964
rect 264888 358912 264940 358964
rect 305644 358912 305696 358964
rect 101404 358844 101456 358896
rect 293132 358844 293184 358896
rect 179236 358776 179288 358828
rect 421564 358776 421616 358828
rect 213920 358708 213972 358760
rect 214472 358708 214524 358760
rect 282920 358708 282972 358760
rect 283564 358708 283616 358760
rect 217048 358096 217100 358148
rect 232504 358096 232556 358148
rect 214564 358028 214616 358080
rect 275008 358028 275060 358080
rect 276940 358028 276992 358080
rect 387708 358028 387760 358080
rect 570512 358028 570564 358080
rect 158628 357756 158680 357808
rect 182916 357756 182968 357808
rect 275652 357756 275704 357808
rect 300860 357756 300912 357808
rect 164148 357688 164200 357740
rect 186780 357688 186832 357740
rect 195244 357688 195296 357740
rect 200028 357688 200080 357740
rect 267004 357688 267056 357740
rect 293224 357688 293276 357740
rect 179880 357620 179932 357672
rect 214472 357620 214524 357672
rect 223488 357620 223540 357672
rect 298100 357620 298152 357672
rect 154488 357552 154540 357604
rect 184940 357552 184992 357604
rect 191748 357552 191800 357604
rect 285680 357552 285732 357604
rect 287428 357552 287480 357604
rect 292212 357552 292264 357604
rect 292304 357552 292356 357604
rect 363604 357552 363656 357604
rect 135904 357484 135956 357536
rect 256792 357484 256844 357536
rect 283564 357484 283616 357536
rect 435088 357484 435140 357536
rect 80060 357416 80112 357468
rect 300952 357416 301004 357468
rect 200028 357348 200080 357400
rect 201500 357348 201552 357400
rect 305092 357348 305144 357400
rect 305736 357348 305788 357400
rect 273536 356736 273588 356788
rect 274548 356736 274600 356788
rect 40040 356668 40092 356720
rect 126980 356668 127032 356720
rect 214564 356668 214616 356720
rect 285680 356668 285732 356720
rect 307760 356668 307812 356720
rect 253940 356396 253992 356448
rect 300124 356396 300176 356448
rect 171048 356328 171100 356380
rect 197728 356328 197780 356380
rect 225420 356328 225472 356380
rect 303620 356328 303672 356380
rect 175924 356260 175976 356312
rect 273536 356260 273588 356312
rect 68836 356192 68888 356244
rect 270500 356192 270552 356244
rect 347044 356192 347096 356244
rect 67548 356124 67600 356176
rect 305092 356124 305144 356176
rect 68928 356056 68980 356108
rect 262772 356056 262824 356108
rect 582840 356056 582892 356108
rect 96620 355104 96672 355156
rect 294052 355104 294104 355156
rect 75920 355036 75972 355088
rect 293040 355036 293092 355088
rect 126428 354968 126480 355020
rect 235080 354968 235132 355020
rect 107660 354900 107712 354952
rect 298192 354900 298244 354952
rect 290464 354832 290516 354884
rect 309784 354832 309836 354884
rect 285956 354764 286008 354816
rect 311900 354764 311952 354816
rect 72424 354696 72476 354748
rect 241704 354696 241756 354748
rect 260748 354696 260800 354748
rect 305000 354696 305052 354748
rect 84292 354016 84344 354068
rect 179788 354016 179840 354068
rect 44824 353948 44876 354000
rect 45468 353948 45520 354000
rect 176660 353948 176712 354000
rect 62028 352520 62080 352572
rect 176108 352520 176160 352572
rect 296168 352520 296220 352572
rect 415768 352520 415820 352572
rect 117964 351228 118016 351280
rect 179880 351228 179932 351280
rect 60648 351160 60700 351212
rect 176016 351160 176068 351212
rect 295340 349800 295392 349852
rect 359464 349800 359516 349852
rect 389088 349800 389140 349852
rect 580356 349800 580408 349852
rect 124956 347760 125008 347812
rect 179512 347760 179564 347812
rect 295984 346400 296036 346452
rect 351184 346400 351236 346452
rect 3516 345176 3568 345228
rect 8944 345176 8996 345228
rect 157248 345040 157300 345092
rect 176660 345040 176712 345092
rect 296076 342864 296128 342916
rect 349804 342864 349856 342916
rect 175188 342252 175240 342304
rect 176844 342252 176896 342304
rect 520924 341504 520976 341556
rect 536104 341504 536156 341556
rect 160744 340892 160796 340944
rect 179328 340892 179380 340944
rect 295340 339464 295392 339516
rect 308404 339464 308456 339516
rect 293868 338104 293920 338156
rect 360844 338104 360896 338156
rect 293224 337356 293276 337408
rect 498844 337356 498896 337408
rect 295340 336676 295392 336728
rect 298284 336676 298336 336728
rect 299388 336676 299440 336728
rect 299388 335996 299440 336048
rect 582932 335996 582984 336048
rect 106280 333956 106332 334008
rect 176844 333956 176896 334008
rect 293960 333956 294012 334008
rect 531964 333956 532016 334008
rect 175096 333684 175148 333736
rect 176660 333684 176712 333736
rect 104164 333208 104216 333260
rect 175096 333208 175148 333260
rect 295340 331848 295392 331900
rect 296904 331848 296956 331900
rect 367744 331848 367796 331900
rect 294328 329808 294380 329860
rect 369124 329808 369176 329860
rect 175096 327088 175148 327140
rect 176660 327088 176712 327140
rect 293040 327088 293092 327140
rect 575572 327088 575624 327140
rect 151728 325660 151780 325712
rect 176660 325660 176712 325712
rect 3424 324912 3476 324964
rect 98644 324912 98696 324964
rect 573548 324300 573600 324352
rect 580172 324300 580224 324352
rect 295340 320152 295392 320204
rect 323584 320152 323636 320204
rect 3424 318792 3476 318844
rect 116584 318792 116636 318844
rect 295340 318792 295392 318844
rect 325056 318792 325108 318844
rect 295340 317364 295392 317416
rect 299572 317364 299624 317416
rect 300768 317364 300820 317416
rect 300768 316684 300820 316736
rect 337476 316684 337528 316736
rect 129280 314644 129332 314696
rect 176660 314644 176712 314696
rect 295340 313896 295392 313948
rect 296812 313896 296864 313948
rect 570052 313896 570104 313948
rect 160560 312536 160612 312588
rect 176660 312536 176712 312588
rect 99380 311856 99432 311908
rect 160560 311856 160612 311908
rect 295340 311856 295392 311908
rect 471244 311856 471296 311908
rect 8944 311108 8996 311160
rect 118700 311108 118752 311160
rect 122104 311108 122156 311160
rect 160744 311108 160796 311160
rect 118700 310428 118752 310480
rect 173164 310428 173216 310480
rect 295340 310428 295392 310480
rect 300952 310428 301004 310480
rect 301320 310428 301372 310480
rect 301320 309748 301372 309800
rect 468484 309748 468536 309800
rect 295340 307776 295392 307828
rect 313280 307776 313332 307828
rect 570236 307776 570288 307828
rect 25504 307028 25556 307080
rect 84384 307028 84436 307080
rect 91100 307028 91152 307080
rect 99380 307028 99432 307080
rect 154396 307028 154448 307080
rect 176476 307028 176528 307080
rect 114744 306348 114796 306400
rect 154396 306348 154448 306400
rect 81440 305124 81492 305176
rect 138756 305124 138808 305176
rect 88432 305056 88484 305108
rect 162124 305056 162176 305108
rect 3240 304988 3292 305040
rect 122196 304988 122248 305040
rect 173808 304988 173860 305040
rect 176660 304988 176712 305040
rect 295340 304988 295392 305040
rect 310612 304988 310664 305040
rect 13084 304920 13136 304972
rect 72240 304920 72292 304972
rect 94504 304920 94556 304972
rect 114744 304920 114796 304972
rect 90364 304716 90416 304768
rect 94596 304716 94648 304768
rect 388996 304240 389048 304292
rect 542360 304240 542412 304292
rect 74540 303628 74592 303680
rect 142896 303628 142948 303680
rect 88340 303560 88392 303612
rect 103796 303560 103848 303612
rect 104164 303560 104216 303612
rect 295340 303560 295392 303612
rect 298192 303560 298244 303612
rect 412640 303560 412692 303612
rect 413284 303560 413336 303612
rect 89720 302404 89772 302456
rect 134708 302404 134760 302456
rect 99380 302336 99432 302388
rect 148324 302336 148376 302388
rect 92848 302268 92900 302320
rect 152556 302268 152608 302320
rect 98736 302200 98788 302252
rect 178684 302200 178736 302252
rect 104164 301180 104216 301232
rect 144184 301180 144236 301232
rect 102140 301112 102192 301164
rect 149796 301112 149848 301164
rect 76104 301044 76156 301096
rect 130568 301044 130620 301096
rect 85580 300976 85632 301028
rect 153844 300976 153896 301028
rect 85672 300908 85724 300960
rect 155224 300908 155276 300960
rect 160008 300908 160060 300960
rect 176660 300908 176712 300960
rect 75368 300840 75420 300892
rect 165068 300840 165120 300892
rect 293224 300840 293276 300892
rect 300216 300840 300268 300892
rect 98000 300772 98052 300824
rect 98644 300772 98696 300824
rect 53748 300092 53800 300144
rect 70952 300092 71004 300144
rect 296076 300092 296128 300144
rect 305092 300092 305144 300144
rect 88340 299752 88392 299804
rect 123484 299752 123536 299804
rect 98552 299684 98604 299736
rect 136088 299684 136140 299736
rect 98000 299616 98052 299668
rect 148416 299616 148468 299668
rect 84384 299548 84436 299600
rect 144368 299548 144420 299600
rect 22836 299480 22888 299532
rect 117964 299480 118016 299532
rect 111064 298732 111116 298784
rect 124220 298732 124272 298784
rect 102876 298392 102928 298444
rect 124864 298392 124916 298444
rect 90640 298324 90692 298376
rect 137284 298324 137336 298376
rect 116584 298256 116636 298308
rect 169116 298256 169168 298308
rect 75184 298188 75236 298240
rect 131764 298188 131816 298240
rect 73252 298120 73304 298172
rect 159364 298120 159416 298172
rect 169760 298052 169812 298104
rect 170956 298052 171008 298104
rect 176660 298052 176712 298104
rect 502340 298052 502392 298104
rect 502984 298052 503036 298104
rect 158444 297372 158496 297424
rect 176660 297372 176712 297424
rect 129648 297032 129700 297084
rect 158444 297032 158496 297084
rect 87420 296964 87472 297016
rect 133236 296964 133288 297016
rect 83556 296896 83608 296948
rect 133144 296896 133196 296948
rect 104348 296828 104400 296880
rect 156696 296828 156748 296880
rect 66168 296760 66220 296812
rect 140228 296760 140280 296812
rect 68560 296692 68612 296744
rect 157340 296692 157392 296744
rect 327724 296692 327776 296744
rect 502340 296692 502392 296744
rect 84200 295672 84252 295724
rect 84476 295672 84528 295724
rect 111892 295672 111944 295724
rect 151176 295672 151228 295724
rect 78404 295604 78456 295656
rect 82268 295536 82320 295588
rect 88984 295536 89036 295588
rect 117228 295604 117280 295656
rect 164976 295604 165028 295656
rect 137376 295536 137428 295588
rect 84476 295468 84528 295520
rect 145564 295468 145616 295520
rect 32404 295400 32456 295452
rect 101404 295400 101456 295452
rect 105452 295400 105504 295452
rect 171140 295400 171192 295452
rect 88984 295332 89036 295384
rect 156604 295332 156656 295384
rect 295340 295332 295392 295384
rect 302884 295332 302936 295384
rect 79692 294652 79744 294704
rect 104164 294652 104216 294704
rect 70032 294584 70084 294636
rect 117228 294584 117280 294636
rect 300216 294584 300268 294636
rect 492404 294584 492456 294636
rect 80980 294380 81032 294432
rect 135996 294380 136048 294432
rect 106096 294312 106148 294364
rect 123576 294312 123628 294364
rect 114468 294244 114520 294296
rect 140136 294244 140188 294296
rect 82912 294176 82964 294228
rect 116860 294176 116912 294228
rect 93860 294108 93912 294160
rect 138848 294108 138900 294160
rect 67456 294040 67508 294092
rect 79324 294040 79376 294092
rect 49608 293972 49660 294024
rect 96436 293972 96488 294024
rect 103796 293972 103848 294024
rect 104532 293972 104584 294024
rect 114560 293972 114612 294024
rect 115388 293972 115440 294024
rect 117228 293972 117280 294024
rect 173164 293972 173216 294024
rect 295340 293972 295392 294024
rect 302148 293972 302200 294024
rect 75920 293904 75972 293956
rect 76748 293904 76800 293956
rect 84292 293904 84344 293956
rect 85212 293904 85264 293956
rect 85580 293904 85632 293956
rect 86500 293904 86552 293956
rect 88340 293904 88392 293956
rect 89076 293904 89128 293956
rect 92572 292884 92624 292936
rect 121000 292884 121052 292936
rect 110604 292816 110656 292868
rect 126336 292816 126388 292868
rect 88064 292748 88116 292800
rect 129096 292748 129148 292800
rect 53656 292680 53708 292732
rect 71964 292680 72016 292732
rect 91928 292680 91980 292732
rect 134616 292680 134668 292732
rect 53104 292612 53156 292664
rect 92572 292612 92624 292664
rect 109316 292612 109368 292664
rect 162216 292612 162268 292664
rect 3424 292544 3476 292596
rect 46204 292544 46256 292596
rect 68744 292544 68796 292596
rect 141516 292544 141568 292596
rect 319536 292544 319588 292596
rect 520740 292544 520792 292596
rect 71688 292476 71740 292528
rect 111156 292476 111208 292528
rect 121460 292476 121512 292528
rect 126428 292476 126480 292528
rect 117320 291932 117372 291984
rect 119712 291932 119764 291984
rect 101312 291864 101364 291916
rect 112812 291864 112864 291916
rect 116860 291864 116912 291916
rect 119344 291864 119396 291916
rect 119988 291864 120040 291916
rect 147036 291796 147088 291848
rect 160744 291796 160796 291848
rect 176660 291796 176712 291848
rect 119988 291320 120040 291372
rect 129188 291320 129240 291372
rect 127716 291252 127768 291304
rect 345664 291252 345716 291304
rect 583852 291320 583904 291372
rect 131856 291184 131908 291236
rect 323676 291184 323728 291236
rect 566464 291184 566516 291236
rect 31024 290436 31076 290488
rect 68744 290436 68796 290488
rect 362224 289960 362276 290012
rect 533620 289960 533672 290012
rect 121460 289892 121512 289944
rect 149704 289892 149756 289944
rect 318156 289892 318208 289944
rect 583668 289892 583720 289944
rect 56416 289824 56468 289876
rect 67640 289824 67692 289876
rect 121552 289824 121604 289876
rect 164884 289824 164936 289876
rect 169024 289824 169076 289876
rect 176660 289824 176712 289876
rect 302148 289824 302200 289876
rect 449900 289824 449952 289876
rect 121460 289756 121512 289808
rect 162308 289756 162360 289808
rect 4068 289076 4120 289128
rect 67456 289076 67508 289128
rect 369308 288532 369360 288584
rect 418988 288532 419040 288584
rect 52368 288464 52420 288516
rect 67732 288464 67784 288516
rect 385868 288464 385920 288516
rect 566556 288464 566608 288516
rect 50988 288396 51040 288448
rect 67640 288396 67692 288448
rect 356796 288396 356848 288448
rect 583576 288396 583628 288448
rect 121460 288328 121512 288380
rect 126244 288328 126296 288380
rect 296720 287648 296772 287700
rect 406108 287648 406160 287700
rect 413284 287648 413336 287700
rect 456984 287648 457036 287700
rect 468484 287648 468536 287700
rect 486424 287648 486476 287700
rect 121460 287580 121512 287632
rect 122196 287580 122248 287632
rect 337384 287104 337436 287156
rect 571616 287104 571668 287156
rect 59268 287036 59320 287088
rect 67640 287036 67692 287088
rect 121552 287036 121604 287088
rect 167736 287036 167788 287088
rect 342904 287036 342956 287088
rect 583116 287036 583168 287088
rect 153108 286288 153160 286340
rect 171784 286288 171836 286340
rect 363788 285812 363840 285864
rect 514300 285812 514352 285864
rect 54944 285744 54996 285796
rect 67732 285744 67784 285796
rect 121644 285744 121696 285796
rect 153108 285744 153160 285796
rect 370596 285744 370648 285796
rect 536840 285744 536892 285796
rect 41328 285676 41380 285728
rect 67640 285676 67692 285728
rect 123668 285676 123720 285728
rect 162768 285676 162820 285728
rect 176660 285676 176712 285728
rect 295340 285676 295392 285728
rect 298928 285676 298980 285728
rect 381544 285676 381596 285728
rect 582748 285676 582800 285728
rect 583300 285676 583352 285728
rect 121460 285608 121512 285660
rect 175924 285608 175976 285660
rect 471244 284928 471296 284980
rect 527180 284928 527232 284980
rect 530584 284928 530636 284980
rect 531964 284928 532016 284980
rect 546500 284928 546552 284980
rect 387616 284588 387668 284640
rect 392584 284588 392636 284640
rect 366364 284520 366416 284572
rect 428648 284520 428700 284572
rect 365076 284452 365128 284504
rect 473084 284452 473136 284504
rect 371884 284384 371936 284436
rect 575480 284384 575532 284436
rect 57888 284316 57940 284368
rect 67640 284316 67692 284368
rect 301504 284316 301556 284368
rect 302056 284316 302108 284368
rect 583484 284316 583536 284368
rect 66168 284248 66220 284300
rect 67824 284248 67876 284300
rect 574284 283772 574336 283824
rect 574744 283772 574796 283824
rect 120816 283568 120868 283620
rect 155868 283568 155920 283620
rect 389916 283228 389968 283280
rect 441528 283228 441580 283280
rect 359648 283160 359700 283212
rect 507860 283160 507912 283212
rect 371976 283092 372028 283144
rect 574284 283092 574336 283144
rect 373356 283024 373408 283076
rect 581184 283024 581236 283076
rect 341524 282956 341576 283008
rect 555516 282956 555568 283008
rect 45376 282888 45428 282940
rect 67732 282888 67784 282940
rect 121460 282888 121512 282940
rect 142988 282888 143040 282940
rect 155868 282888 155920 282940
rect 176660 282888 176712 282940
rect 295340 282888 295392 282940
rect 569960 282888 570012 282940
rect 573548 282888 573600 282940
rect 64788 282820 64840 282872
rect 67640 282820 67692 282872
rect 121000 282140 121052 282192
rect 158720 282140 158772 282192
rect 374828 281868 374880 281920
rect 438308 281868 438360 281920
rect 374736 281800 374788 281852
rect 482744 281800 482796 281852
rect 369216 281732 369268 281784
rect 523960 281732 524012 281784
rect 377496 281664 377548 281716
rect 567844 281664 567896 281716
rect 568396 281664 568448 281716
rect 384212 281596 384264 281648
rect 576952 281596 577004 281648
rect 577504 281596 577556 281648
rect 121460 281528 121512 281580
rect 157984 281528 158036 281580
rect 158720 281528 158772 281580
rect 159916 281528 159968 281580
rect 176660 281528 176712 281580
rect 295340 281528 295392 281580
rect 295524 281528 295576 281580
rect 356704 281528 356756 281580
rect 362316 281528 362368 281580
rect 582472 281528 582524 281580
rect 157156 281460 157208 281512
rect 157340 281460 157392 281512
rect 121552 280780 121604 280832
rect 167828 280780 167880 280832
rect 169116 280780 169168 280832
rect 175280 280780 175332 280832
rect 377680 280508 377732 280560
rect 397092 280508 397144 280560
rect 367928 280440 367980 280492
rect 409236 280440 409288 280492
rect 376024 280372 376076 280424
rect 469864 280372 469916 280424
rect 297548 280304 297600 280356
rect 425428 280304 425480 280356
rect 573456 280304 573508 280356
rect 389640 280236 389692 280288
rect 574192 280236 574244 280288
rect 53748 280168 53800 280220
rect 67640 280168 67692 280220
rect 121460 280168 121512 280220
rect 138940 280168 138992 280220
rect 157156 280168 157208 280220
rect 326344 280168 326396 280220
rect 581092 280168 581144 280220
rect 176660 280100 176712 280152
rect 378876 279080 378928 279132
rect 393872 279080 393924 279132
rect 381636 279012 381688 279064
rect 403532 279012 403584 279064
rect 300216 278944 300268 278996
rect 447968 278944 448020 278996
rect 583760 278944 583812 278996
rect 373264 278876 373316 278928
rect 400312 278876 400364 278928
rect 421564 278876 421616 278928
rect 421840 278876 421892 278928
rect 581644 278876 581696 278928
rect 121460 278808 121512 278860
rect 151084 278808 151136 278860
rect 158536 278808 158588 278860
rect 171140 278808 171192 278860
rect 35808 278740 35860 278792
rect 67640 278740 67692 278792
rect 121552 278740 121604 278792
rect 171784 278740 171836 278792
rect 295340 278808 295392 278860
rect 298836 278808 298888 278860
rect 391940 278808 391992 278860
rect 580448 278808 580500 278860
rect 379428 278740 379480 278792
rect 583392 278740 583444 278792
rect 176660 278672 176712 278724
rect 501420 278672 501472 278724
rect 502340 278672 502392 278724
rect 538864 278672 538916 278724
rect 543280 278672 543332 278724
rect 563704 278672 563756 278724
rect 565176 278672 565228 278724
rect 577596 278672 577648 278724
rect 580264 278672 580316 278724
rect 352564 278060 352616 278112
rect 384212 278060 384264 278112
rect 314016 277992 314068 278044
rect 385868 277992 385920 278044
rect 65984 277788 66036 277840
rect 68100 277788 68152 277840
rect 389824 277720 389876 277772
rect 549076 277720 549128 277772
rect 364984 277652 365036 277704
rect 431868 277652 431920 277704
rect 452660 277652 452712 277704
rect 489184 277652 489236 277704
rect 385684 277584 385736 277636
rect 453764 277584 453816 277636
rect 486424 277584 486476 277636
rect 576216 277584 576268 277636
rect 380164 277516 380216 277568
rect 495624 277516 495676 277568
rect 121552 277448 121604 277500
rect 133328 277448 133380 277500
rect 385776 277448 385828 277500
rect 517520 277448 517572 277500
rect 63408 277380 63460 277432
rect 67640 277380 67692 277432
rect 121460 277380 121512 277432
rect 163504 277380 163556 277432
rect 566464 277040 566516 277092
rect 568672 277040 568724 277092
rect 301320 276632 301372 276684
rect 381544 276632 381596 276684
rect 382188 276632 382240 276684
rect 391940 276632 391992 276684
rect 566556 276632 566608 276684
rect 571524 276632 571576 276684
rect 410340 276360 410392 276412
rect 582656 276360 582708 276412
rect 385868 276292 385920 276344
rect 466644 276292 466696 276344
rect 382924 276224 382976 276276
rect 530400 276224 530452 276276
rect 367836 276156 367888 276208
rect 412548 276156 412600 276208
rect 52276 276088 52328 276140
rect 67732 276088 67784 276140
rect 121552 276088 121604 276140
rect 147220 276088 147272 276140
rect 383016 276088 383068 276140
rect 570144 276088 570196 276140
rect 48228 276020 48280 276072
rect 67640 276020 67692 276072
rect 121460 276020 121512 276072
rect 170588 276020 170640 276072
rect 172336 276020 172388 276072
rect 175280 276020 175332 276072
rect 295340 276020 295392 276072
rect 300952 276020 301004 276072
rect 301320 276020 301372 276072
rect 353944 276020 353996 276072
rect 354588 276020 354640 276072
rect 571340 276020 571392 276072
rect 177488 275952 177540 276004
rect 363604 275952 363656 276004
rect 364248 275952 364300 276004
rect 410340 275952 410392 276004
rect 295984 275340 296036 275392
rect 409696 275544 409748 275596
rect 370504 275272 370556 275324
rect 389640 275272 389692 275324
rect 452660 275544 452712 275596
rect 580172 275272 580224 275324
rect 389732 275204 389784 275256
rect 389916 275204 389968 275256
rect 64696 274728 64748 274780
rect 67640 274728 67692 274780
rect 121460 274728 121512 274780
rect 126244 274728 126296 274780
rect 121552 274660 121604 274712
rect 145748 274660 145800 274712
rect 295340 274660 295392 274712
rect 298744 274660 298796 274712
rect 121460 274592 121512 274644
rect 166264 274592 166316 274644
rect 385040 274592 385092 274644
rect 22744 273912 22796 273964
rect 60096 273912 60148 273964
rect 61936 273300 61988 273352
rect 67640 273300 67692 273352
rect 60096 273232 60148 273284
rect 60372 273232 60424 273284
rect 67732 273232 67784 273284
rect 121460 273232 121512 273284
rect 141424 273232 141476 273284
rect 345756 273232 345808 273284
rect 386880 273232 386932 273284
rect 121000 272484 121052 272536
rect 124220 272484 124272 272536
rect 160100 272484 160152 272536
rect 121460 272008 121512 272060
rect 125048 272008 125100 272060
rect 64788 271872 64840 271924
rect 67640 271872 67692 271924
rect 160100 271872 160152 271924
rect 161204 271872 161256 271924
rect 176660 271872 176712 271924
rect 295340 271872 295392 271924
rect 306472 271872 306524 271924
rect 381544 271872 381596 271924
rect 64604 271804 64656 271856
rect 67732 271804 67784 271856
rect 325056 271124 325108 271176
rect 350540 271124 350592 271176
rect 46848 270512 46900 270564
rect 67640 270512 67692 270564
rect 121460 270512 121512 270564
rect 130660 270512 130712 270564
rect 140688 269764 140740 269816
rect 169024 269764 169076 269816
rect 366456 269764 366508 269816
rect 387156 269764 387208 269816
rect 121552 269152 121604 269204
rect 125140 269152 125192 269204
rect 49516 269084 49568 269136
rect 67640 269084 67692 269136
rect 121460 269084 121512 269136
rect 143080 269084 143132 269136
rect 295340 269084 295392 269136
rect 325056 269084 325108 269136
rect 66168 268200 66220 268252
rect 68192 268200 68244 268252
rect 13084 267724 13136 267776
rect 57612 267724 57664 267776
rect 67640 267724 67692 267776
rect 161388 267724 161440 267776
rect 176660 267724 176712 267776
rect 57244 267656 57296 267708
rect 68928 267656 68980 267708
rect 62764 267044 62816 267096
rect 63316 267044 63368 267096
rect 67640 267044 67692 267096
rect 298928 267044 298980 267096
rect 328460 267044 328512 267096
rect 306288 266976 306340 267028
rect 389732 266976 389784 267028
rect 3056 266364 3108 266416
rect 25504 266364 25556 266416
rect 121460 266364 121512 266416
rect 166448 266364 166500 266416
rect 165620 266296 165672 266348
rect 176660 266296 176712 266348
rect 45468 265616 45520 265668
rect 60740 265616 60792 265668
rect 60740 265004 60792 265056
rect 61844 265004 61896 265056
rect 67640 265004 67692 265056
rect 48136 264936 48188 264988
rect 67732 264936 67784 264988
rect 121460 264936 121512 264988
rect 166264 264936 166316 264988
rect 59176 264188 59228 264240
rect 67640 264188 67692 264240
rect 295340 264188 295392 264240
rect 331864 264188 331916 264240
rect 50896 263644 50948 263696
rect 67640 263644 67692 263696
rect 121460 263644 121512 263696
rect 136180 263644 136232 263696
rect 21364 263576 21416 263628
rect 59176 263576 59228 263628
rect 121552 263576 121604 263628
rect 163596 263576 163648 263628
rect 121460 263508 121512 263560
rect 146944 263508 146996 263560
rect 140228 262964 140280 263016
rect 162308 262964 162360 263016
rect 146944 262896 146996 262948
rect 169116 262896 169168 262948
rect 36544 262828 36596 262880
rect 57796 262828 57848 262880
rect 122196 262828 122248 262880
rect 169024 262828 169076 262880
rect 57796 262284 57848 262336
rect 67732 262284 67784 262336
rect 56508 262216 56560 262268
rect 67640 262216 67692 262268
rect 121460 262216 121512 262268
rect 141608 262216 141660 262268
rect 331956 262216 332008 262268
rect 386880 262216 386932 262268
rect 121460 261468 121512 261520
rect 143540 261468 143592 261520
rect 144460 261468 144512 261520
rect 162308 261468 162360 261520
rect 162676 261468 162728 261520
rect 176660 261468 176712 261520
rect 295340 261128 295392 261180
rect 297456 261128 297508 261180
rect 66076 260924 66128 260976
rect 68192 260924 68244 260976
rect 56324 260856 56376 260908
rect 67732 260856 67784 260908
rect 121552 260856 121604 260908
rect 155316 260856 155368 260908
rect 39948 260788 40000 260840
rect 67640 260788 67692 260840
rect 360844 260788 360896 260840
rect 386880 260788 386932 260840
rect 572628 260788 572680 260840
rect 581184 260788 581236 260840
rect 575572 260720 575624 260772
rect 576308 260720 576360 260772
rect 122380 260108 122432 260160
rect 165160 260108 165212 260160
rect 121460 259496 121512 259548
rect 146944 259496 146996 259548
rect 63224 259428 63276 259480
rect 67640 259428 67692 259480
rect 121552 259428 121604 259480
rect 153936 259428 153988 259480
rect 166908 259428 166960 259480
rect 176660 259428 176712 259480
rect 576308 258680 576360 258732
rect 580172 258680 580224 258732
rect 60464 258136 60516 258188
rect 67640 258136 67692 258188
rect 121460 258136 121512 258188
rect 148508 258136 148560 258188
rect 54852 258068 54904 258120
rect 67732 258068 67784 258120
rect 121552 258068 121604 258120
rect 167644 258068 167696 258120
rect 60648 258000 60700 258052
rect 67640 258000 67692 258052
rect 17224 257320 17276 257372
rect 60648 257320 60700 257372
rect 156512 257320 156564 257372
rect 179052 257320 179104 257372
rect 121552 256776 121604 256828
rect 144276 256776 144328 256828
rect 55128 256708 55180 256760
rect 67640 256708 67692 256760
rect 121460 256708 121512 256760
rect 175924 256708 175976 256760
rect 360844 256708 360896 256760
rect 363788 256708 363840 256760
rect 121552 255348 121604 255400
rect 149888 255348 149940 255400
rect 60556 255280 60608 255332
rect 67640 255280 67692 255332
rect 121460 255280 121512 255332
rect 159456 255280 159508 255332
rect 355416 255280 355468 255332
rect 386880 255280 386932 255332
rect 2780 254056 2832 254108
rect 4804 254056 4856 254108
rect 157340 253988 157392 254040
rect 158444 253988 158496 254040
rect 176660 253988 176712 254040
rect 63132 253920 63184 253972
rect 67732 253920 67784 253972
rect 121460 253920 121512 253972
rect 171876 253920 171928 253972
rect 295616 253920 295668 253972
rect 298928 253920 298980 253972
rect 60740 253852 60792 253904
rect 62028 253852 62080 253904
rect 67640 253852 67692 253904
rect 302148 253852 302200 253904
rect 306380 253852 306432 253904
rect 26884 253172 26936 253224
rect 60740 253172 60792 253224
rect 64512 253172 64564 253224
rect 68284 253172 68336 253224
rect 298836 253172 298888 253224
rect 299572 253172 299624 253224
rect 121552 252628 121604 252680
rect 152648 252628 152700 252680
rect 121460 252560 121512 252612
rect 170404 252560 170456 252612
rect 327816 252560 327868 252612
rect 386880 252560 386932 252612
rect 297180 252220 297232 252272
rect 301504 252220 301556 252272
rect 60648 251812 60700 251864
rect 68376 251812 68428 251864
rect 121460 251268 121512 251320
rect 137468 251268 137520 251320
rect 121552 251200 121604 251252
rect 174636 251200 174688 251252
rect 572628 251132 572680 251184
rect 582472 251132 582524 251184
rect 120724 250996 120776 251048
rect 124956 250996 125008 251048
rect 64604 249840 64656 249892
rect 67640 249840 67692 249892
rect 59084 249772 59136 249824
rect 67732 249772 67784 249824
rect 121460 249772 121512 249824
rect 131948 249772 132000 249824
rect 55036 249704 55088 249756
rect 67640 249704 67692 249756
rect 57796 248412 57848 248464
rect 67640 248412 67692 248464
rect 121460 248412 121512 248464
rect 174544 248412 174596 248464
rect 572628 248208 572680 248260
rect 576952 248208 577004 248260
rect 122288 247664 122340 247716
rect 167000 247664 167052 247716
rect 301320 247664 301372 247716
rect 307668 247664 307720 247716
rect 378784 247664 378836 247716
rect 62028 247120 62080 247172
rect 67640 247120 67692 247172
rect 59176 247052 59228 247104
rect 67732 247052 67784 247104
rect 121460 247052 121512 247104
rect 126428 247052 126480 247104
rect 295524 247052 295576 247104
rect 301044 247052 301096 247104
rect 301320 247052 301372 247104
rect 379428 246984 379480 247036
rect 386880 246984 386932 247036
rect 353300 246372 353352 246424
rect 379428 246372 379480 246424
rect 295524 246304 295576 246356
rect 298192 246304 298244 246356
rect 358084 246304 358136 246356
rect 121460 245760 121512 245812
rect 140228 245760 140280 245812
rect 121552 245692 121604 245744
rect 147128 245692 147180 245744
rect 124128 245624 124180 245676
rect 176660 245624 176712 245676
rect 50344 245556 50396 245608
rect 68100 245556 68152 245608
rect 582748 245556 582800 245608
rect 583668 245556 583720 245608
rect 342996 244876 343048 244928
rect 387524 244876 387576 244928
rect 121460 244332 121512 244384
rect 160100 244332 160152 244384
rect 65892 244264 65944 244316
rect 68008 244264 68060 244316
rect 121552 244264 121604 244316
rect 173256 244264 173308 244316
rect 577504 244264 577556 244316
rect 582748 244264 582800 244316
rect 121460 244196 121512 244248
rect 140044 244196 140096 244248
rect 295800 244196 295852 244248
rect 353300 244196 353352 244248
rect 363788 243516 363840 243568
rect 364248 243516 364300 243568
rect 386604 243516 386656 243568
rect 121552 242904 121604 242956
rect 166356 242904 166408 242956
rect 121644 242836 121696 242888
rect 130476 242836 130528 242888
rect 120908 242224 120960 242276
rect 149980 242224 150032 242276
rect 121460 242156 121512 242208
rect 160744 242156 160796 242208
rect 296720 242156 296772 242208
rect 333980 242156 334032 242208
rect 337476 242156 337528 242208
rect 387156 242156 387208 242208
rect 61752 241612 61804 241664
rect 67640 241612 67692 241664
rect 168380 241476 168432 241528
rect 169668 241476 169720 241528
rect 177580 241476 177632 241528
rect 161204 241408 161256 241460
rect 377680 241408 377732 241460
rect 572628 241408 572680 241460
rect 582564 241408 582616 241460
rect 141516 240728 141568 240780
rect 298928 240728 298980 240780
rect 335360 240728 335412 240780
rect 173808 240592 173860 240644
rect 180432 240592 180484 240644
rect 184020 240592 184072 240644
rect 291936 240592 291988 240644
rect 293316 240592 293368 240644
rect 3424 240116 3476 240168
rect 14464 240116 14516 240168
rect 121460 240116 121512 240168
rect 148600 240116 148652 240168
rect 363604 240116 363656 240168
rect 386880 240116 386932 240168
rect 159916 240048 159968 240100
rect 362316 240048 362368 240100
rect 180432 239980 180484 240032
rect 359648 239980 359700 240032
rect 167000 239912 167052 239964
rect 298744 239912 298796 239964
rect 179512 239844 179564 239896
rect 180018 239844 180070 239896
rect 289820 239844 289872 239896
rect 294236 239844 294288 239896
rect 63224 239368 63276 239420
rect 76564 239368 76616 239420
rect 111064 239368 111116 239420
rect 295616 239368 295668 239420
rect 121552 238892 121604 238944
rect 148968 238892 149020 238944
rect 110420 238824 110472 238876
rect 110604 238824 110656 238876
rect 142804 238824 142856 238876
rect 148416 238824 148468 238876
rect 195980 238824 196032 238876
rect 61844 238756 61896 238808
rect 180892 238756 180944 238808
rect 255228 238756 255280 238808
rect 387064 238756 387116 238808
rect 25504 238688 25556 238740
rect 86776 238688 86828 238740
rect 114468 238688 114520 238740
rect 125600 238688 125652 238740
rect 172336 238688 172388 238740
rect 374828 238688 374880 238740
rect 81624 238620 81676 238672
rect 279516 238620 279568 238672
rect 287888 238620 287940 238672
rect 377588 238620 377640 238672
rect 58624 238552 58676 238604
rect 82268 238552 82320 238604
rect 82912 238552 82964 238604
rect 111064 238552 111116 238604
rect 117688 238552 117740 238604
rect 250812 238552 250864 238604
rect 273996 238552 274048 238604
rect 377496 238552 377548 238604
rect 86776 238484 86828 238536
rect 210424 238484 210476 238536
rect 278044 238484 278096 238536
rect 365076 238484 365128 238536
rect 118332 238416 118384 238468
rect 240508 238416 240560 238468
rect 250812 238416 250864 238468
rect 300216 238416 300268 238468
rect 89352 238348 89404 238400
rect 138664 238348 138716 238400
rect 204812 238348 204864 238400
rect 255228 238348 255280 238400
rect 263048 238348 263100 238400
rect 297548 238348 297600 238400
rect 77116 238076 77168 238128
rect 106924 238076 106976 238128
rect 253112 238076 253164 238128
rect 263600 238076 263652 238128
rect 63316 238008 63368 238060
rect 117228 238008 117280 238060
rect 236276 238008 236328 238060
rect 273904 238008 273956 238060
rect 79048 237396 79100 237448
rect 86224 237396 86276 237448
rect 14464 237328 14516 237380
rect 103520 237328 103572 237380
rect 104716 237328 104768 237380
rect 113180 237328 113232 237380
rect 354680 237328 354732 237380
rect 355416 237328 355468 237380
rect 109684 237260 109736 237312
rect 140688 237260 140740 237312
rect 365168 237260 365220 237312
rect 99012 237192 99064 237244
rect 121000 237192 121052 237244
rect 157156 237192 157208 237244
rect 345664 237192 345716 237244
rect 175924 237124 175976 237176
rect 295432 237124 295484 237176
rect 269856 237056 269908 237108
rect 319536 237056 319588 237108
rect 169116 236716 169168 236768
rect 192484 236716 192536 236768
rect 64512 236648 64564 236700
rect 98644 236648 98696 236700
rect 167828 236648 167880 236700
rect 273260 236648 273312 236700
rect 67548 235900 67600 235952
rect 381636 235900 381688 235952
rect 4804 235832 4856 235884
rect 112536 235832 112588 235884
rect 129004 235832 129056 235884
rect 154396 235832 154448 235884
rect 373356 235832 373408 235884
rect 119712 235764 119764 235816
rect 323676 235764 323728 235816
rect 72608 235696 72660 235748
rect 123668 235696 123720 235748
rect 162768 235696 162820 235748
rect 366456 235696 366508 235748
rect 91284 235628 91336 235680
rect 129280 235628 129332 235680
rect 174636 235628 174688 235680
rect 273996 235628 274048 235680
rect 113824 235560 113876 235612
rect 152464 235560 152516 235612
rect 265624 235560 265676 235612
rect 310520 235560 310572 235612
rect 56324 235220 56376 235272
rect 116584 235220 116636 235272
rect 380900 234812 380952 234864
rect 381636 234812 381688 234864
rect 63132 234540 63184 234592
rect 263048 234540 263100 234592
rect 572628 234540 572680 234592
rect 581092 234540 581144 234592
rect 69296 234472 69348 234524
rect 219256 234472 219308 234524
rect 369216 234472 369268 234524
rect 95792 234404 95844 234456
rect 126980 234404 127032 234456
rect 140136 233996 140188 234048
rect 273996 233996 274048 234048
rect 69112 233928 69164 233980
rect 69756 233928 69808 233980
rect 74540 233928 74592 233980
rect 75184 233928 75236 233980
rect 80060 233928 80112 233980
rect 80980 233928 81032 233980
rect 84200 233928 84252 233980
rect 84844 233928 84896 233980
rect 95148 233928 95200 233980
rect 120724 233928 120776 233980
rect 242256 233928 242308 233980
rect 386512 233928 386564 233980
rect 64604 233860 64656 233912
rect 86960 233860 87012 233912
rect 88064 233860 88116 233912
rect 95240 233860 95292 233912
rect 96436 233860 96488 233912
rect 100760 233860 100812 233912
rect 101588 233860 101640 233912
rect 107660 233860 107712 233912
rect 108672 233860 108724 233912
rect 114560 233860 114612 233912
rect 115756 233860 115808 233912
rect 148968 233860 149020 233912
rect 311164 233860 311216 233912
rect 361028 233860 361080 233912
rect 386788 233860 386840 233912
rect 95884 233792 95936 233844
rect 61660 233180 61712 233232
rect 341524 233180 341576 233232
rect 86132 233112 86184 233164
rect 157248 233112 157300 233164
rect 184020 233112 184072 233164
rect 295616 233112 295668 233164
rect 76472 233044 76524 233096
rect 134524 233044 134576 233096
rect 144368 233044 144420 233096
rect 254676 233044 254728 233096
rect 273260 233044 273312 233096
rect 325700 233112 325752 233164
rect 326344 233112 326396 233164
rect 70676 232568 70728 232620
rect 88984 232568 89036 232620
rect 170496 232568 170548 232620
rect 186964 232568 187016 232620
rect 1308 232500 1360 232552
rect 120080 232500 120132 232552
rect 155316 232500 155368 232552
rect 275284 232500 275336 232552
rect 129280 231752 129332 231804
rect 367928 231752 367980 231804
rect 82268 231684 82320 231736
rect 278044 231684 278096 231736
rect 279516 231684 279568 231736
rect 280068 231684 280120 231736
rect 309140 231684 309192 231736
rect 104716 231616 104768 231668
rect 293224 231616 293276 231668
rect 91928 231548 91980 231600
rect 135904 231548 135956 231600
rect 149888 231548 149940 231600
rect 189080 231548 189132 231600
rect 189724 231548 189776 231600
rect 215208 231548 215260 231600
rect 363696 231548 363748 231600
rect 173256 231140 173308 231192
rect 246304 231140 246356 231192
rect 88708 231072 88760 231124
rect 315396 231072 315448 231124
rect 107384 230392 107436 230444
rect 151728 230392 151780 230444
rect 169668 230392 169720 230444
rect 371884 230392 371936 230444
rect 158444 230324 158496 230376
rect 327724 230324 327776 230376
rect 233884 230256 233936 230308
rect 353944 230256 353996 230308
rect 163596 230188 163648 230240
rect 269856 230188 269908 230240
rect 166448 229848 166500 229900
rect 203616 229848 203668 229900
rect 151728 229780 151780 229832
rect 242164 229780 242216 229832
rect 65984 229712 66036 229764
rect 380348 229712 380400 229764
rect 386420 229712 386472 229764
rect 83556 229032 83608 229084
rect 130384 229032 130436 229084
rect 162676 229032 162728 229084
rect 387800 229032 387852 229084
rect 60372 228964 60424 229016
rect 242256 228964 242308 229016
rect 167736 228896 167788 228948
rect 333244 228896 333296 228948
rect 137376 228828 137428 228880
rect 223580 228828 223632 228880
rect 352564 228828 352616 228880
rect 387156 228692 387208 228744
rect 387708 228692 387760 228744
rect 387800 228420 387852 228472
rect 388444 228420 388496 228472
rect 7564 228352 7616 228404
rect 83556 228352 83608 228404
rect 332692 228284 332744 228336
rect 333244 228284 333296 228336
rect 52368 227672 52420 227724
rect 345020 227672 345072 227724
rect 345756 227672 345808 227724
rect 160744 227604 160796 227656
rect 318156 227604 318208 227656
rect 572628 227332 572680 227384
rect 576860 227332 576912 227384
rect 177672 227264 177724 227316
rect 196624 227264 196676 227316
rect 61752 227196 61804 227248
rect 198004 227196 198056 227248
rect 195980 227128 196032 227180
rect 353944 227128 353996 227180
rect 48136 227060 48188 227112
rect 269764 227060 269816 227112
rect 67364 226992 67416 227044
rect 386972 226992 387024 227044
rect 48228 226244 48280 226296
rect 361028 226244 361080 226296
rect 133328 226176 133380 226228
rect 378876 226176 378928 226228
rect 158536 226108 158588 226160
rect 342904 226108 342956 226160
rect 54852 225632 54904 225684
rect 160744 225632 160796 225684
rect 170588 225632 170640 225684
rect 243544 225632 243596 225684
rect 271880 225632 271932 225684
rect 294144 225632 294196 225684
rect 100300 225564 100352 225616
rect 222844 225564 222896 225616
rect 256700 225564 256752 225616
rect 268384 225564 268436 225616
rect 291844 225564 291896 225616
rect 316040 225564 316092 225616
rect 360292 225428 360344 225480
rect 361028 225428 361080 225480
rect 378140 225156 378192 225208
rect 378876 225156 378928 225208
rect 149980 224884 150032 224936
rect 360200 224884 360252 224936
rect 148508 224816 148560 224868
rect 276020 224816 276072 224868
rect 347136 224816 347188 224868
rect 347780 224816 347832 224868
rect 360200 224476 360252 224528
rect 360844 224476 360896 224528
rect 276020 224408 276072 224460
rect 276664 224408 276716 224460
rect 59084 223524 59136 223576
rect 327172 223524 327224 223576
rect 327816 223524 327868 223576
rect 153844 223456 153896 223508
rect 385132 223524 385184 223576
rect 385868 223524 385920 223576
rect 145748 223388 145800 223440
rect 298192 223388 298244 223440
rect 125140 222912 125192 222964
rect 220084 222912 220136 222964
rect 56416 222844 56468 222896
rect 117964 222844 118016 222896
rect 165160 222844 165212 222896
rect 278136 222844 278188 222896
rect 45376 222096 45428 222148
rect 342352 222096 342404 222148
rect 342996 222096 343048 222148
rect 162308 222028 162360 222080
rect 263600 222028 263652 222080
rect 264244 222028 264296 222080
rect 310428 222028 310480 222080
rect 314016 222028 314068 222080
rect 141424 221620 141476 221672
rect 211896 221620 211948 221672
rect 131856 221552 131908 221604
rect 247684 221552 247736 221604
rect 87420 221484 87472 221536
rect 207664 221484 207716 221536
rect 3424 221416 3476 221468
rect 120172 221416 120224 221468
rect 151176 221416 151228 221468
rect 310428 221416 310480 221468
rect 144460 220736 144512 220788
rect 386880 220736 386932 220788
rect 156696 220668 156748 220720
rect 385040 220668 385092 220720
rect 385776 220668 385828 220720
rect 102876 220192 102928 220244
rect 252744 220192 252796 220244
rect 69204 220124 69256 220176
rect 251180 220124 251232 220176
rect 50896 220056 50948 220108
rect 356060 220056 356112 220108
rect 153936 219376 153988 219428
rect 363788 219376 363840 219428
rect 576216 219376 576268 219428
rect 580080 219376 580132 219428
rect 155868 219308 155920 219360
rect 360936 219308 360988 219360
rect 57704 218832 57756 218884
rect 162768 218832 162820 218884
rect 53656 218764 53708 218816
rect 153844 218764 153896 218816
rect 160744 218764 160796 218816
rect 274640 218764 274692 218816
rect 137468 218696 137520 218748
rect 338212 218696 338264 218748
rect 153108 217948 153160 218000
rect 270500 217948 270552 218000
rect 114560 217472 114612 217524
rect 289084 217472 289136 217524
rect 77392 217404 77444 217456
rect 252836 217404 252888 217456
rect 280896 217404 280948 217456
rect 311900 217404 311952 217456
rect 52276 217336 52328 217388
rect 233884 217336 233936 217388
rect 248420 217336 248472 217388
rect 291200 217336 291252 217388
rect 169024 217268 169076 217320
rect 357992 217268 358044 217320
rect 270500 216656 270552 216708
rect 271236 216656 271288 216708
rect 242164 216588 242216 216640
rect 387524 216588 387576 216640
rect 357992 216520 358044 216572
rect 358176 216520 358228 216572
rect 373264 216520 373316 216572
rect 141608 216112 141660 216164
rect 261484 216112 261536 216164
rect 104992 216044 105044 216096
rect 283656 216044 283708 216096
rect 70400 215976 70452 216028
rect 249800 215976 249852 216028
rect 92572 215908 92624 215960
rect 314016 215908 314068 215960
rect 3332 215228 3384 215280
rect 21364 215228 21416 215280
rect 162768 215228 162820 215280
rect 287704 215228 287756 215280
rect 155224 214752 155276 214804
rect 256700 214752 256752 214804
rect 100852 214684 100904 214736
rect 263600 214684 263652 214736
rect 325056 214684 325108 214736
rect 349160 214684 349212 214736
rect 96712 214616 96764 214668
rect 336740 214616 336792 214668
rect 76564 214548 76616 214600
rect 330484 214548 330536 214600
rect 64696 213868 64748 213920
rect 331312 213868 331364 213920
rect 331956 213868 332008 213920
rect 130568 213324 130620 213376
rect 191104 213324 191156 213376
rect 202144 213324 202196 213376
rect 283564 213324 283616 213376
rect 127716 213256 127768 213308
rect 270500 213256 270552 213308
rect 60464 213188 60516 213240
rect 238024 213188 238076 213240
rect 273996 213188 274048 213240
rect 346400 213188 346452 213240
rect 347688 213188 347740 213240
rect 347688 212508 347740 212560
rect 386880 212508 386932 212560
rect 572628 212508 572680 212560
rect 582748 212508 582800 212560
rect 148600 211964 148652 212016
rect 242164 211964 242216 212016
rect 111800 211896 111852 211948
rect 273260 211896 273312 211948
rect 92480 211828 92532 211880
rect 259552 211828 259604 211880
rect 88984 211760 89036 211812
rect 312544 211760 312596 211812
rect 323584 211760 323636 211812
rect 340972 211760 341024 211812
rect 344284 211760 344336 211812
rect 387156 211760 387208 211812
rect 572628 211080 572680 211132
rect 583576 211080 583628 211132
rect 142896 210672 142948 210724
rect 229744 210672 229796 210724
rect 95884 210604 95936 210656
rect 166172 210604 166224 210656
rect 203524 210604 203576 210656
rect 340144 210604 340196 210656
rect 137284 210536 137336 210588
rect 277400 210536 277452 210588
rect 103612 210468 103664 210520
rect 352564 210468 352616 210520
rect 78680 210400 78732 210452
rect 329840 210400 329892 210452
rect 80152 209380 80204 209432
rect 162308 209380 162360 209432
rect 144184 209312 144236 209364
rect 280160 209312 280212 209364
rect 86224 209244 86276 209296
rect 240784 209244 240836 209296
rect 136088 209176 136140 209228
rect 327080 209176 327132 209228
rect 327908 209176 327960 209228
rect 49516 209108 49568 209160
rect 269304 209108 269356 209160
rect 107752 209040 107804 209092
rect 335544 209040 335596 209092
rect 327908 208360 327960 208412
rect 386880 208360 386932 208412
rect 149704 207816 149756 207868
rect 259460 207816 259512 207868
rect 86960 207748 87012 207800
rect 252652 207748 252704 207800
rect 84384 207680 84436 207732
rect 267740 207680 267792 207732
rect 60556 207612 60608 207664
rect 336832 207612 336884 207664
rect 572444 206932 572496 206984
rect 575480 206932 575532 206984
rect 143080 206524 143132 206576
rect 265072 206524 265124 206576
rect 89812 206456 89864 206508
rect 249892 206456 249944 206508
rect 65892 206388 65944 206440
rect 255412 206388 255464 206440
rect 281540 206388 281592 206440
rect 342260 206388 342312 206440
rect 118700 206320 118752 206372
rect 315488 206320 315540 206372
rect 57888 206252 57940 206304
rect 300216 206252 300268 206304
rect 351276 205640 351328 205692
rect 386880 205640 386932 205692
rect 576216 205640 576268 205692
rect 580908 205640 580960 205692
rect 162124 205164 162176 205216
rect 225604 205164 225656 205216
rect 107660 205096 107712 205148
rect 167736 205096 167788 205148
rect 224960 205096 225012 205148
rect 308496 205096 308548 205148
rect 166172 205028 166224 205080
rect 281540 205028 281592 205080
rect 53748 204960 53800 205012
rect 238116 204960 238168 205012
rect 134708 204892 134760 204944
rect 340144 204892 340196 204944
rect 571524 203872 571576 203924
rect 574284 203872 574336 203924
rect 145564 203736 145616 203788
rect 235264 203736 235316 203788
rect 73252 203668 73304 203720
rect 148416 203668 148468 203720
rect 149796 203668 149848 203720
rect 278780 203668 278832 203720
rect 315304 203668 315356 203720
rect 360844 203668 360896 203720
rect 129188 203600 129240 203652
rect 347872 203600 347924 203652
rect 69020 203532 69072 203584
rect 324320 203532 324372 203584
rect 147036 202376 147088 202428
rect 239404 202376 239456 202428
rect 129096 202308 129148 202360
rect 232504 202308 232556 202360
rect 245660 202308 245712 202360
rect 309876 202308 309928 202360
rect 126336 202240 126388 202292
rect 264980 202240 265032 202292
rect 110512 202172 110564 202224
rect 255596 202172 255648 202224
rect 340144 202172 340196 202224
rect 386880 202172 386932 202224
rect 159364 202104 159416 202156
rect 347964 202104 348016 202156
rect 96620 200948 96672 201000
rect 160100 200948 160152 201000
rect 136180 200880 136232 200932
rect 262312 200880 262364 200932
rect 140228 200812 140280 200864
rect 269212 200812 269264 200864
rect 103704 200744 103756 200796
rect 322940 200744 322992 200796
rect 100760 199588 100812 199640
rect 255504 199588 255556 199640
rect 318064 199588 318116 199640
rect 335452 199588 335504 199640
rect 162216 199520 162268 199572
rect 318156 199520 318208 199572
rect 116584 199452 116636 199504
rect 333244 199452 333296 199504
rect 120724 199384 120776 199436
rect 340236 199384 340288 199436
rect 572628 198636 572680 198688
rect 579712 198636 579764 198688
rect 151084 198228 151136 198280
rect 233976 198228 234028 198280
rect 261484 198228 261536 198280
rect 334164 198228 334216 198280
rect 138940 198160 138992 198212
rect 260932 198160 260984 198212
rect 269764 198160 269816 198212
rect 347780 198160 347832 198212
rect 133236 198092 133288 198144
rect 277492 198092 277544 198144
rect 57796 198024 57848 198076
rect 276112 198024 276164 198076
rect 99380 197956 99432 198008
rect 345296 197956 345348 198008
rect 300124 197276 300176 197328
rect 382188 197276 382240 197328
rect 386880 197276 386932 197328
rect 152648 196868 152700 196920
rect 262404 196868 262456 196920
rect 124864 196800 124916 196852
rect 273352 196800 273404 196852
rect 80060 196732 80112 196784
rect 319536 196732 319588 196784
rect 93952 196664 94004 196716
rect 343732 196664 343784 196716
rect 69112 196596 69164 196648
rect 320824 196596 320876 196648
rect 130660 195440 130712 195492
rect 196716 195440 196768 195492
rect 160100 195372 160152 195424
rect 261024 195372 261076 195424
rect 192484 195304 192536 195356
rect 370596 195304 370648 195356
rect 153844 195236 153896 195288
rect 338856 195236 338908 195288
rect 147128 194080 147180 194132
rect 270592 194080 270644 194132
rect 134616 194012 134668 194064
rect 258172 194012 258224 194064
rect 63408 193944 63460 193996
rect 160744 193944 160796 193996
rect 227720 193944 227772 193996
rect 351920 193944 351972 193996
rect 115940 193876 115992 193928
rect 249064 193876 249116 193928
rect 74632 193808 74684 193860
rect 321652 193808 321704 193860
rect 330484 193808 330536 193860
rect 386420 193808 386472 193860
rect 583852 193128 583904 193180
rect 583852 192924 583904 192976
rect 246304 192856 246356 192908
rect 349344 192856 349396 192908
rect 148324 192788 148376 192840
rect 271972 192788 272024 192840
rect 120816 192720 120868 192772
rect 246396 192720 246448 192772
rect 89720 192652 89772 192704
rect 249984 192652 250036 192704
rect 189724 192584 189776 192636
rect 354036 192584 354088 192636
rect 138756 192516 138808 192568
rect 345204 192516 345256 192568
rect 71780 192448 71832 192500
rect 343824 192448 343876 192500
rect 306288 191836 306340 191888
rect 334072 191836 334124 191888
rect 278136 191768 278188 191820
rect 571708 191700 571760 191752
rect 574192 191700 574244 191752
rect 231860 191360 231912 191412
rect 278044 191360 278096 191412
rect 163504 191292 163556 191344
rect 324412 191292 324464 191344
rect 56508 191224 56560 191276
rect 242256 191224 242308 191276
rect 273904 191224 273956 191276
rect 358084 191224 358136 191276
rect 142988 191156 143040 191208
rect 358820 191156 358872 191208
rect 84292 191088 84344 191140
rect 321560 191088 321612 191140
rect 324964 191088 325016 191140
rect 329104 191088 329156 191140
rect 102048 190476 102100 190528
rect 192484 190476 192536 190528
rect 324412 190408 324464 190460
rect 380256 190408 380308 190460
rect 333244 190340 333296 190392
rect 387064 190340 387116 190392
rect 126428 190000 126480 190052
rect 246488 190000 246540 190052
rect 152556 189932 152608 189984
rect 273444 189932 273496 189984
rect 117964 189864 118016 189916
rect 209044 189864 209096 189916
rect 210424 189864 210476 189916
rect 332048 189864 332100 189916
rect 40684 189796 40736 189848
rect 109684 189796 109736 189848
rect 171784 189796 171836 189848
rect 324504 189796 324556 189848
rect 62028 189728 62080 189780
rect 259644 189728 259696 189780
rect 103428 189048 103480 189100
rect 171968 189048 172020 189100
rect 3424 188980 3476 189032
rect 53104 188980 53156 189032
rect 324504 188980 324556 189032
rect 325056 188980 325108 189032
rect 383016 188980 383068 189032
rect 243544 188572 243596 188624
rect 330484 188572 330536 188624
rect 156604 188504 156656 188556
rect 246304 188504 246356 188556
rect 138848 188436 138900 188488
rect 247776 188436 247828 188488
rect 144276 188368 144328 188420
rect 262220 188368 262272 188420
rect 135996 188300 136048 188352
rect 274732 188300 274784 188352
rect 100668 187688 100720 187740
rect 171784 187688 171836 187740
rect 329196 187620 329248 187672
rect 386788 187620 386840 187672
rect 572628 187620 572680 187672
rect 583484 187620 583536 187672
rect 330484 187552 330536 187604
rect 370504 187552 370556 187604
rect 161388 187144 161440 187196
rect 195244 187144 195296 187196
rect 104900 187076 104952 187128
rect 188344 187076 188396 187128
rect 162308 187008 162360 187060
rect 327264 187008 327316 187060
rect 95240 186940 95292 186992
rect 320180 186940 320232 186992
rect 126888 186328 126940 186380
rect 169116 186328 169168 186380
rect 131948 185852 132000 185904
rect 243544 185852 243596 185904
rect 170404 185784 170456 185836
rect 324964 185784 325016 185836
rect 60648 185716 60700 185768
rect 254032 185716 254084 185768
rect 102140 185648 102192 185700
rect 323124 185648 323176 185700
rect 66076 185580 66128 185632
rect 324504 185580 324556 185632
rect 329196 185580 329248 185632
rect 386880 185580 386932 185632
rect 115848 184968 115900 185020
rect 170496 184968 170548 185020
rect 122748 184900 122800 184952
rect 211988 184900 212040 184952
rect 571432 184832 571484 184884
rect 574100 184832 574152 184884
rect 160008 184424 160060 184476
rect 189724 184424 189776 184476
rect 126244 184356 126296 184408
rect 266544 184356 266596 184408
rect 148416 184288 148468 184340
rect 337476 184288 337528 184340
rect 84200 184220 84252 184272
rect 321836 184220 321888 184272
rect 77300 184152 77352 184204
rect 318064 184152 318116 184204
rect 119988 183540 120040 183592
rect 170680 183540 170732 183592
rect 237380 182996 237432 183048
rect 271144 182996 271196 183048
rect 93860 182928 93912 182980
rect 253940 182928 253992 182980
rect 283656 182928 283708 182980
rect 342536 182928 342588 182980
rect 167644 182860 167696 182912
rect 339500 182860 339552 182912
rect 106924 182792 106976 182844
rect 350632 182792 350684 182844
rect 130752 182248 130804 182300
rect 206376 182248 206428 182300
rect 110696 182180 110748 182232
rect 214564 182180 214616 182232
rect 341524 182180 341576 182232
rect 386420 182180 386472 182232
rect 222844 181636 222896 181688
rect 266452 181636 266504 181688
rect 311164 181636 311216 181688
rect 341064 181636 341116 181688
rect 211068 181568 211120 181620
rect 220820 181568 220872 181620
rect 225604 181568 225656 181620
rect 335636 181568 335688 181620
rect 171876 181500 171928 181552
rect 251272 181500 251324 181552
rect 271236 181500 271288 181552
rect 381636 181500 381688 181552
rect 154488 181432 154540 181484
rect 198004 181432 198056 181484
rect 203616 181432 203668 181484
rect 356888 181432 356940 181484
rect 121092 180956 121144 181008
rect 166540 180956 166592 181008
rect 112996 180888 113048 180940
rect 167736 180888 167788 180940
rect 128084 180820 128136 180872
rect 214656 180820 214708 180872
rect 242164 180412 242216 180464
rect 256792 180412 256844 180464
rect 240784 180344 240836 180396
rect 258356 180344 258408 180396
rect 166908 180276 166960 180328
rect 182824 180276 182876 180328
rect 238116 180276 238168 180328
rect 263692 180276 263744 180328
rect 315396 180276 315448 180328
rect 346492 180276 346544 180328
rect 158628 180208 158680 180260
rect 184204 180208 184256 180260
rect 209044 180208 209096 180260
rect 272064 180208 272116 180260
rect 300216 180208 300268 180260
rect 345112 180208 345164 180260
rect 66168 180140 66220 180192
rect 251364 180140 251416 180192
rect 280068 180140 280120 180192
rect 380440 180140 380492 180192
rect 68928 180072 68980 180124
rect 321744 180072 321796 180124
rect 132040 179528 132092 179580
rect 165344 179528 165396 179580
rect 110236 179460 110288 179512
rect 167828 179460 167880 179512
rect 114376 179392 114428 179444
rect 210424 179392 210476 179444
rect 246488 178984 246540 179036
rect 252560 178984 252612 179036
rect 247776 178916 247828 178968
rect 249340 178916 249392 178968
rect 233976 178848 234028 178900
rect 249432 178848 249484 178900
rect 220084 178780 220136 178832
rect 265164 178780 265216 178832
rect 317328 178780 317380 178832
rect 337384 178780 337436 178832
rect 211896 178712 211948 178764
rect 258080 178712 258132 178764
rect 289084 178712 289136 178764
rect 325792 178712 325844 178764
rect 146944 178644 146996 178696
rect 254124 178644 254176 178696
rect 305644 178644 305696 178696
rect 363696 178644 363748 178696
rect 318064 178508 318116 178560
rect 323032 178508 323084 178560
rect 148232 178236 148284 178288
rect 166448 178236 166500 178288
rect 123024 178168 123076 178220
rect 169300 178168 169352 178220
rect 118424 178100 118476 178152
rect 166632 178100 166684 178152
rect 129464 178032 129516 178084
rect 214196 178032 214248 178084
rect 326436 177964 326488 178016
rect 386880 177964 386932 178016
rect 572076 177964 572128 178016
rect 576308 177964 576360 178016
rect 258172 177760 258224 177812
rect 242256 177556 242308 177608
rect 258264 177556 258316 177608
rect 171048 177488 171100 177540
rect 215944 177488 215996 177540
rect 239404 177488 239456 177540
rect 256976 177488 257028 177540
rect 196716 177420 196768 177472
rect 249248 177420 249300 177472
rect 314016 177556 314068 177608
rect 332784 177556 332836 177608
rect 311256 177488 311308 177540
rect 338764 177488 338816 177540
rect 269120 177420 269172 177472
rect 275284 177420 275336 177472
rect 328552 177420 328604 177472
rect 164884 177352 164936 177404
rect 251456 177352 251508 177404
rect 264244 177352 264296 177404
rect 365076 177352 365128 177404
rect 166356 177284 166408 177336
rect 325884 177284 325936 177336
rect 104624 177012 104676 177064
rect 170588 177012 170640 177064
rect 133144 176944 133196 176996
rect 164516 176944 164568 176996
rect 128176 176876 128228 176928
rect 165436 176876 165488 176928
rect 108120 176808 108172 176860
rect 169024 176808 169076 176860
rect 107016 176740 107068 176792
rect 171876 176740 171928 176792
rect 158996 176672 159048 176724
rect 166264 176672 166316 176724
rect 135720 176604 135772 176656
rect 213920 176604 213972 176656
rect 235264 176604 235316 176656
rect 248052 176604 248104 176656
rect 324320 176604 324372 176656
rect 380348 176604 380400 176656
rect 246304 176536 246356 176588
rect 255320 176536 255372 176588
rect 134432 176196 134484 176248
rect 165528 176196 165580 176248
rect 124496 176128 124548 176180
rect 167920 176128 167972 176180
rect 319536 176128 319588 176180
rect 334256 176128 334308 176180
rect 116952 176060 117004 176112
rect 169208 176060 169260 176112
rect 312544 176060 312596 176112
rect 327356 176060 327408 176112
rect 98368 175992 98420 176044
rect 170404 175992 170456 176044
rect 307024 175992 307076 176044
rect 343640 175992 343692 176044
rect 4804 175924 4856 175976
rect 110420 175924 110472 175976
rect 160744 175924 160796 175976
rect 259736 175924 259788 175976
rect 283564 175924 283616 175976
rect 329932 175924 329984 175976
rect 243544 175788 243596 175840
rect 249156 175788 249208 175840
rect 164516 175176 164568 175228
rect 214012 175176 214064 175228
rect 324320 175176 324372 175228
rect 360292 175176 360344 175228
rect 165528 175108 165580 175160
rect 213920 175108 213972 175160
rect 3700 163480 3752 163532
rect 4068 163480 4120 163532
rect 66904 163480 66956 163532
rect 3424 150356 3476 150408
rect 31024 150356 31076 150408
rect 3240 137912 3292 137964
rect 17224 137912 17276 137964
rect 60648 128324 60700 128376
rect 66076 128324 66128 128376
rect 57888 125604 57940 125656
rect 66168 125604 66220 125656
rect 63316 122816 63368 122868
rect 66076 122816 66128 122868
rect 63408 121456 63460 121508
rect 66168 121456 66220 121508
rect 2780 110712 2832 110764
rect 4804 110712 4856 110764
rect 3424 97588 3476 97640
rect 7564 97588 7616 97640
rect 165436 174496 165488 174548
rect 214104 174496 214156 174548
rect 283748 174020 283800 174072
rect 307300 174020 307352 174072
rect 274088 173952 274140 174004
rect 306748 173952 306800 174004
rect 264244 173884 264296 173936
rect 307668 173884 307720 173936
rect 165344 173816 165396 173868
rect 213920 173816 213972 173868
rect 354036 173816 354088 173868
rect 387156 173816 387208 173868
rect 387616 173816 387668 173868
rect 206376 173748 206428 173800
rect 214012 173748 214064 173800
rect 283656 172660 283708 172712
rect 307576 172660 307628 172712
rect 269764 172592 269816 172644
rect 307300 172592 307352 172644
rect 261668 172524 261720 172576
rect 307668 172524 307720 172576
rect 324320 172456 324372 172508
rect 385132 172456 385184 172508
rect 251824 171844 251876 171896
rect 258080 171844 258132 171896
rect 167000 171776 167052 171828
rect 214656 171776 214708 171828
rect 289452 171232 289504 171284
rect 306932 171232 306984 171284
rect 268476 171164 268528 171216
rect 307668 171164 307720 171216
rect 262864 171096 262916 171148
rect 306564 171096 306616 171148
rect 324872 171096 324924 171148
rect 354036 171096 354088 171148
rect 169116 171028 169168 171080
rect 213920 171028 213972 171080
rect 251732 171028 251784 171080
rect 256700 171028 256752 171080
rect 324320 171028 324372 171080
rect 382280 171028 382332 171080
rect 356888 170280 356940 170332
rect 359648 170280 359700 170332
rect 282276 169872 282328 169924
rect 307668 169872 307720 169924
rect 251824 169804 251876 169856
rect 259644 169804 259696 169856
rect 265624 169804 265676 169856
rect 307300 169804 307352 169856
rect 257344 169736 257396 169788
rect 306748 169736 306800 169788
rect 324320 169736 324372 169788
rect 356796 169736 356848 169788
rect 572628 169736 572680 169788
rect 576860 169736 576912 169788
rect 167920 169668 167972 169720
rect 213920 169668 213972 169720
rect 324504 169668 324556 169720
rect 329196 169668 329248 169720
rect 332048 169668 332100 169720
rect 386880 169668 386932 169720
rect 169300 169600 169352 169652
rect 214012 169600 214064 169652
rect 252468 169600 252520 169652
rect 261024 169600 261076 169652
rect 324320 168988 324372 169040
rect 327264 168988 327316 169040
rect 331956 168988 332008 169040
rect 279424 168444 279476 168496
rect 306748 168444 306800 168496
rect 258908 168376 258960 168428
rect 307300 168376 307352 168428
rect 166540 168308 166592 168360
rect 213920 168308 213972 168360
rect 252376 168308 252428 168360
rect 262404 168308 262456 168360
rect 324320 168308 324372 168360
rect 380900 168308 380952 168360
rect 211988 168240 212040 168292
rect 214012 168240 214064 168292
rect 324412 168240 324464 168292
rect 324688 168240 324740 168292
rect 376024 168240 376076 168292
rect 252468 168172 252520 168224
rect 256976 168172 257028 168224
rect 271236 167628 271288 167680
rect 307576 167628 307628 167680
rect 252468 167220 252520 167272
rect 258172 167220 258224 167272
rect 279608 167084 279660 167136
rect 307668 167084 307720 167136
rect 262956 167016 263008 167068
rect 307484 167016 307536 167068
rect 166632 166948 166684 167000
rect 214104 166948 214156 167000
rect 252468 166948 252520 167000
rect 258264 166948 258316 167000
rect 324320 166948 324372 167000
rect 344284 166948 344336 167000
rect 169208 166880 169260 166932
rect 214012 166880 214064 166932
rect 170680 166812 170732 166864
rect 213920 166812 213972 166864
rect 252376 166812 252428 166864
rect 256792 166812 256844 166864
rect 252284 166268 252336 166320
rect 259552 166268 259604 166320
rect 337476 166268 337528 166320
rect 386880 166268 386932 166320
rect 278228 165724 278280 165776
rect 306564 165724 306616 165776
rect 268568 165656 268620 165708
rect 307668 165656 307720 165708
rect 257528 165588 257580 165640
rect 307484 165588 307536 165640
rect 572352 165588 572404 165640
rect 574100 165588 574152 165640
rect 170496 165520 170548 165572
rect 213920 165520 213972 165572
rect 252468 165520 252520 165572
rect 264980 165520 265032 165572
rect 252468 164976 252520 165028
rect 259736 164976 259788 165028
rect 264428 164840 264480 164892
rect 307300 164840 307352 164892
rect 292028 164296 292080 164348
rect 307576 164296 307628 164348
rect 324320 164296 324372 164348
rect 337384 164296 337436 164348
rect 275284 164228 275336 164280
rect 307668 164228 307720 164280
rect 323400 164228 323452 164280
rect 380256 164228 380308 164280
rect 167736 164160 167788 164212
rect 213920 164160 213972 164212
rect 252192 164160 252244 164212
rect 262312 164160 262364 164212
rect 324320 164160 324372 164212
rect 333244 164160 333296 164212
rect 210424 164092 210476 164144
rect 214012 164092 214064 164144
rect 324412 164092 324464 164144
rect 330576 164092 330628 164144
rect 260380 163480 260432 163532
rect 307392 163480 307444 163532
rect 289268 162936 289320 162988
rect 307484 162936 307536 162988
rect 261484 162868 261536 162920
rect 307668 162868 307720 162920
rect 167828 162800 167880 162852
rect 213920 162800 213972 162852
rect 252100 162800 252152 162852
rect 265164 162800 265216 162852
rect 380440 162800 380492 162852
rect 386880 162800 386932 162852
rect 252468 162732 252520 162784
rect 263692 162732 263744 162784
rect 260840 162120 260892 162172
rect 284944 162120 284996 162172
rect 325884 162120 325936 162172
rect 369216 162120 369268 162172
rect 251548 162052 251600 162104
rect 252836 162052 252888 162104
rect 287704 161576 287756 161628
rect 306748 161576 306800 161628
rect 281080 161508 281132 161560
rect 307668 161508 307720 161560
rect 260104 161440 260156 161492
rect 307484 161440 307536 161492
rect 169024 161372 169076 161424
rect 213920 161372 213972 161424
rect 171876 161304 171928 161356
rect 214012 161304 214064 161356
rect 177764 160692 177816 160744
rect 216036 160692 216088 160744
rect 324320 160692 324372 160744
rect 331496 160692 331548 160744
rect 251548 160216 251600 160268
rect 254216 160216 254268 160268
rect 297548 160216 297600 160268
rect 307668 160216 307720 160268
rect 263140 160148 263192 160200
rect 306748 160148 306800 160200
rect 257436 160080 257488 160132
rect 307576 160080 307628 160132
rect 170588 160012 170640 160064
rect 213920 160012 213972 160064
rect 324320 159332 324372 159384
rect 327356 159332 327408 159384
rect 367928 159332 367980 159384
rect 289084 158856 289136 158908
rect 307668 158856 307720 158908
rect 261576 158788 261628 158840
rect 307576 158788 307628 158840
rect 253296 158720 253348 158772
rect 307484 158720 307536 158772
rect 359648 158720 359700 158772
rect 380348 158720 380400 158772
rect 572628 158720 572680 158772
rect 575480 158720 575532 158772
rect 171968 158652 172020 158704
rect 213920 158652 213972 158704
rect 252468 158652 252520 158704
rect 273444 158652 273496 158704
rect 324412 158652 324464 158704
rect 360200 158652 360252 158704
rect 324320 158584 324372 158636
rect 359648 158584 359700 158636
rect 279700 157972 279752 158024
rect 307300 157972 307352 158024
rect 265716 157428 265768 157480
rect 307484 157428 307536 157480
rect 258816 157360 258868 157412
rect 307668 157360 307720 157412
rect 171784 157292 171836 157344
rect 214012 157292 214064 157344
rect 324320 157292 324372 157344
rect 385040 157292 385092 157344
rect 192484 157224 192536 157276
rect 213920 157224 213972 157276
rect 324412 157224 324464 157276
rect 345296 157224 345348 157276
rect 346308 157224 346360 157276
rect 251180 157088 251232 157140
rect 254032 157088 254084 157140
rect 251364 157020 251416 157072
rect 254124 157020 254176 157072
rect 290648 156612 290700 156664
rect 307576 156612 307628 156664
rect 346308 156612 346360 156664
rect 377496 156612 377548 156664
rect 267004 156000 267056 156052
rect 307668 156000 307720 156052
rect 257620 155932 257672 155984
rect 306748 155932 306800 155984
rect 170404 155864 170456 155916
rect 213920 155864 213972 155916
rect 251824 155864 251876 155916
rect 277400 155864 277452 155916
rect 324320 155864 324372 155916
rect 342444 155864 342496 155916
rect 252468 155796 252520 155848
rect 267740 155796 267792 155848
rect 252376 155728 252428 155780
rect 263600 155728 263652 155780
rect 252284 155252 252336 155304
rect 266544 155252 266596 155304
rect 287888 155252 287940 155304
rect 306932 155252 306984 155304
rect 264980 155184 265032 155236
rect 293132 155184 293184 155236
rect 342444 155184 342496 155236
rect 384396 155184 384448 155236
rect 574744 155184 574796 155236
rect 580356 155184 580408 155236
rect 300216 154640 300268 154692
rect 307668 154640 307720 154692
rect 260288 154572 260340 154624
rect 307484 154572 307536 154624
rect 252468 154504 252520 154556
rect 269304 154504 269356 154556
rect 324320 154504 324372 154556
rect 346492 154504 346544 154556
rect 347688 154504 347740 154556
rect 324412 154436 324464 154488
rect 334256 154436 334308 154488
rect 334624 154436 334676 154488
rect 252100 154300 252152 154352
rect 257344 154300 257396 154352
rect 347688 153892 347740 153944
rect 360936 153892 360988 153944
rect 276020 153824 276072 153876
rect 291936 153824 291988 153876
rect 334624 153824 334676 153876
rect 385776 153824 385828 153876
rect 575388 153824 575440 153876
rect 581000 153824 581052 153876
rect 296260 153348 296312 153400
rect 307668 153348 307720 153400
rect 192484 153280 192536 153332
rect 213920 153280 213972 153332
rect 264336 153280 264388 153332
rect 307576 153280 307628 153332
rect 177304 153212 177356 153264
rect 214012 153212 214064 153264
rect 258724 153212 258776 153264
rect 306564 153212 306616 153264
rect 324964 153212 325016 153264
rect 376024 153212 376076 153264
rect 572628 153212 572680 153264
rect 575388 153212 575440 153264
rect 252376 153144 252428 153196
rect 272064 153144 272116 153196
rect 349804 153144 349856 153196
rect 386880 153144 386932 153196
rect 252468 153076 252520 153128
rect 270500 153076 270552 153128
rect 254584 153008 254636 153060
rect 255412 153008 255464 153060
rect 256240 152464 256292 152516
rect 305000 152464 305052 152516
rect 273996 151920 274048 151972
rect 307668 151920 307720 151972
rect 202236 151852 202288 151904
rect 213920 151852 213972 151904
rect 257344 151852 257396 151904
rect 306564 151852 306616 151904
rect 171784 151784 171836 151836
rect 214012 151784 214064 151836
rect 254124 151784 254176 151836
rect 307576 151784 307628 151836
rect 252468 151716 252520 151768
rect 273260 151716 273312 151768
rect 324320 151716 324372 151768
rect 337476 151716 337528 151768
rect 251916 151648 251968 151700
rect 266452 151648 266504 151700
rect 167644 151036 167696 151088
rect 205640 151036 205692 151088
rect 250628 151036 250680 151088
rect 259460 151036 259512 151088
rect 572628 151036 572680 151088
rect 579620 151036 579672 151088
rect 304356 150560 304408 150612
rect 307668 150560 307720 150612
rect 211896 150492 211948 150544
rect 214012 150492 214064 150544
rect 289360 150492 289412 150544
rect 307484 150492 307536 150544
rect 203616 150424 203668 150476
rect 213920 150424 213972 150476
rect 256056 150424 256108 150476
rect 307576 150424 307628 150476
rect 324412 150424 324464 150476
rect 333888 150424 333940 150476
rect 335544 150424 335596 150476
rect 579620 150424 579672 150476
rect 580264 150424 580316 150476
rect 166448 150356 166500 150408
rect 214012 150356 214064 150408
rect 324320 150356 324372 150408
rect 331312 150356 331364 150408
rect 334164 150356 334216 150408
rect 386604 150356 386656 150408
rect 205640 150288 205692 150340
rect 213920 150288 213972 150340
rect 324412 150288 324464 150340
rect 338212 150288 338264 150340
rect 251180 150152 251232 150204
rect 253940 150152 253992 150204
rect 295984 149676 296036 149728
rect 307208 149676 307260 149728
rect 338212 149676 338264 149728
rect 388444 149676 388496 149728
rect 260196 149064 260248 149116
rect 307484 149064 307536 149116
rect 329196 149064 329248 149116
rect 334164 149064 334216 149116
rect 166264 148996 166316 149048
rect 213920 148996 213972 149048
rect 252468 148996 252520 149048
rect 278780 148996 278832 149048
rect 177856 148316 177908 148368
rect 216128 148316 216180 148368
rect 272616 147772 272668 147824
rect 307576 147772 307628 147824
rect 269856 147704 269908 147756
rect 307668 147704 307720 147756
rect 254676 147636 254728 147688
rect 307484 147636 307536 147688
rect 322848 147636 322900 147688
rect 382924 147636 382976 147688
rect 252376 147568 252428 147620
rect 281540 147568 281592 147620
rect 324320 147568 324372 147620
rect 335636 147568 335688 147620
rect 380164 147568 380216 147620
rect 252468 147500 252520 147552
rect 277492 147500 277544 147552
rect 251732 147432 251784 147484
rect 255504 147432 255556 147484
rect 571708 147296 571760 147348
rect 574744 147296 574796 147348
rect 251548 146956 251600 147008
rect 265072 146956 265124 147008
rect 256148 146888 256200 146940
rect 306932 146888 306984 146940
rect 301596 146412 301648 146464
rect 307668 146412 307720 146464
rect 185584 146344 185636 146396
rect 213920 146344 213972 146396
rect 283840 146344 283892 146396
rect 307576 146344 307628 146396
rect 166264 146276 166316 146328
rect 214012 146276 214064 146328
rect 263048 146276 263100 146328
rect 307484 146276 307536 146328
rect 252100 146208 252152 146260
rect 274640 146208 274692 146260
rect 342444 146208 342496 146260
rect 387064 146208 387116 146260
rect 252284 146140 252336 146192
rect 258356 146140 258408 146192
rect 330576 145596 330628 145648
rect 342444 145596 342496 145648
rect 193864 145528 193916 145580
rect 214104 145528 214156 145580
rect 324320 145528 324372 145580
rect 336832 145528 336884 145580
rect 337476 145528 337528 145580
rect 254860 145052 254912 145104
rect 306932 145052 306984 145104
rect 204904 144984 204956 145036
rect 214012 144984 214064 145036
rect 255964 144984 256016 145036
rect 306564 144984 306616 145036
rect 167644 144916 167696 144968
rect 213920 144916 213972 144968
rect 373264 144916 373316 144968
rect 386604 144916 386656 144968
rect 251916 144848 251968 144900
rect 270592 144848 270644 144900
rect 324412 144848 324464 144900
rect 330484 144848 330536 144900
rect 252468 144780 252520 144832
rect 262220 144780 262272 144832
rect 324320 144780 324372 144832
rect 327172 144780 327224 144832
rect 274640 144236 274692 144288
rect 295340 144236 295392 144288
rect 254768 144168 254820 144220
rect 307392 144168 307444 144220
rect 328368 144168 328420 144220
rect 339500 144168 339552 144220
rect 212080 143624 212132 143676
rect 214656 143624 214708 143676
rect 298744 143624 298796 143676
rect 306932 143624 306984 143676
rect 189816 143556 189868 143608
rect 213920 143556 213972 143608
rect 293408 143556 293460 143608
rect 307668 143556 307720 143608
rect 572628 143556 572680 143608
rect 575572 143556 575624 143608
rect 252376 143488 252428 143540
rect 274732 143488 274784 143540
rect 324412 143488 324464 143540
rect 332692 143488 332744 143540
rect 338856 143488 338908 143540
rect 385684 143488 385736 143540
rect 252468 143420 252520 143472
rect 269212 143420 269264 143472
rect 324320 143352 324372 143404
rect 326344 143352 326396 143404
rect 251824 142808 251876 142860
rect 265716 142808 265768 142860
rect 210516 142672 210568 142724
rect 213920 142672 213972 142724
rect 301504 142264 301556 142316
rect 306748 142264 306800 142316
rect 278320 142196 278372 142248
rect 307484 142196 307536 142248
rect 267096 142128 267148 142180
rect 307668 142128 307720 142180
rect 360108 142128 360160 142180
rect 380164 142128 380216 142180
rect 252468 142060 252520 142112
rect 260932 142060 260984 142112
rect 324412 142060 324464 142112
rect 345204 142060 345256 142112
rect 384304 142060 384356 142112
rect 324320 141992 324372 142044
rect 359556 141992 359608 142044
rect 360108 141992 360160 142044
rect 275468 141448 275520 141500
rect 298100 141448 298152 141500
rect 253480 141380 253532 141432
rect 307116 141380 307168 141432
rect 186964 140836 187016 140888
rect 214012 140836 214064 140888
rect 173348 140768 173400 140820
rect 213920 140768 213972 140820
rect 299112 140768 299164 140820
rect 307668 140768 307720 140820
rect 252100 140700 252152 140752
rect 280160 140700 280212 140752
rect 324320 140700 324372 140752
rect 358176 140700 358228 140752
rect 251732 140632 251784 140684
rect 273352 140632 273404 140684
rect 167828 140020 167880 140072
rect 211896 140020 211948 140072
rect 252192 140020 252244 140072
rect 279424 140020 279476 140072
rect 373448 140020 373500 140072
rect 387616 140020 387668 140072
rect 251732 139748 251784 139800
rect 255596 139748 255648 139800
rect 211988 139476 212040 139528
rect 214656 139476 214708 139528
rect 282368 139476 282420 139528
rect 307576 139476 307628 139528
rect 202144 139408 202196 139460
rect 213920 139408 213972 139460
rect 253388 139408 253440 139460
rect 307668 139408 307720 139460
rect 572628 139408 572680 139460
rect 582656 139408 582708 139460
rect 251364 138728 251416 138780
rect 254584 138728 254636 138780
rect 271420 138660 271472 138712
rect 307300 138660 307352 138712
rect 188436 138048 188488 138100
rect 213920 138048 213972 138100
rect 171876 137980 171928 138032
rect 214012 137980 214064 138032
rect 250536 137980 250588 138032
rect 306932 137980 306984 138032
rect 322848 137980 322900 138032
rect 384304 137980 384356 138032
rect 574744 137980 574796 138032
rect 580172 137980 580224 138032
rect 252468 137912 252520 137964
rect 276112 137912 276164 137964
rect 324320 137912 324372 137964
rect 328552 137912 328604 137964
rect 373264 137912 373316 137964
rect 572628 137912 572680 137964
rect 583024 137912 583076 137964
rect 252100 137844 252152 137896
rect 271972 137844 272024 137896
rect 324412 137844 324464 137896
rect 329840 137844 329892 137896
rect 330300 137844 330352 137896
rect 252008 137300 252060 137352
rect 267004 137300 267056 137352
rect 177488 137232 177540 137284
rect 214748 137232 214800 137284
rect 264520 137232 264572 137284
rect 306564 137232 306616 137284
rect 330300 137232 330352 137284
rect 388628 137232 388680 137284
rect 279424 136688 279476 136740
rect 306932 136688 306984 136740
rect 250444 136620 250496 136672
rect 307668 136620 307720 136672
rect 252376 136552 252428 136604
rect 283748 136552 283800 136604
rect 324320 136552 324372 136604
rect 343824 136552 343876 136604
rect 344468 136552 344520 136604
rect 252100 136484 252152 136536
rect 274088 136484 274140 136536
rect 324412 136484 324464 136536
rect 338856 136484 338908 136536
rect 251732 136416 251784 136468
rect 264244 136416 264296 136468
rect 369124 135940 369176 135992
rect 386420 135940 386472 135992
rect 386696 135940 386748 135992
rect 344468 135872 344520 135924
rect 385684 135872 385736 135924
rect 273904 135464 273956 135516
rect 306932 135464 306984 135516
rect 285036 135396 285088 135448
rect 307484 135396 307536 135448
rect 170404 135328 170456 135380
rect 213920 135328 213972 135380
rect 283564 135328 283616 135380
rect 307576 135328 307628 135380
rect 169116 135260 169168 135312
rect 214012 135260 214064 135312
rect 304264 135260 304316 135312
rect 307668 135260 307720 135312
rect 252468 135192 252520 135244
rect 283656 135192 283708 135244
rect 324320 135192 324372 135244
rect 347964 135192 348016 135244
rect 388536 135192 388588 135244
rect 252284 135124 252336 135176
rect 269764 135124 269816 135176
rect 324412 135124 324464 135176
rect 353300 135124 353352 135176
rect 364984 135124 365036 135176
rect 325516 134512 325568 134564
rect 366364 134512 366416 134564
rect 282184 133968 282236 134020
rect 306748 133968 306800 134020
rect 207756 133900 207808 133952
rect 213920 133900 213972 133952
rect 271328 133900 271380 133952
rect 307668 133900 307720 133952
rect 252376 133832 252428 133884
rect 289452 133832 289504 133884
rect 324320 133832 324372 133884
rect 341064 133832 341116 133884
rect 341248 133832 341300 133884
rect 251732 133764 251784 133816
rect 262864 133764 262916 133816
rect 252468 133696 252520 133748
rect 261668 133696 261720 133748
rect 341248 133220 341300 133272
rect 359556 133220 359608 133272
rect 261760 133152 261812 133204
rect 307392 133152 307444 133204
rect 337476 133152 337528 133204
rect 387616 133152 387668 133204
rect 289176 132540 289228 132592
rect 307484 132540 307536 132592
rect 173256 132472 173308 132524
rect 213920 132472 213972 132524
rect 280988 132472 281040 132524
rect 306932 132472 306984 132524
rect 252468 132404 252520 132456
rect 268476 132404 268528 132456
rect 324320 132404 324372 132456
rect 358820 132404 358872 132456
rect 373448 132404 373500 132456
rect 324412 132336 324464 132388
rect 347136 132336 347188 132388
rect 278780 131724 278832 131776
rect 293040 131724 293092 131776
rect 373264 131724 373316 131776
rect 386420 131724 386472 131776
rect 252468 131588 252520 131640
rect 260380 131588 260432 131640
rect 290556 131248 290608 131300
rect 307484 131248 307536 131300
rect 286416 131180 286468 131232
rect 307576 131180 307628 131232
rect 192576 131112 192628 131164
rect 213920 131112 213972 131164
rect 262864 131112 262916 131164
rect 307668 131112 307720 131164
rect 328368 131112 328420 131164
rect 378876 131112 378928 131164
rect 252468 131044 252520 131096
rect 282276 131044 282328 131096
rect 324412 131044 324464 131096
rect 332784 131044 332836 131096
rect 252376 130976 252428 131028
rect 265624 130976 265676 131028
rect 324320 130976 324372 131028
rect 328368 130976 328420 131028
rect 332784 130364 332836 130416
rect 381728 130364 381780 130416
rect 572628 130160 572680 130212
rect 577596 130160 577648 130212
rect 303160 129956 303212 130008
rect 306748 129956 306800 130008
rect 298928 129888 298980 129940
rect 307668 129888 307720 129940
rect 286324 129820 286376 129872
rect 307116 129820 307168 129872
rect 265716 129752 265768 129804
rect 307576 129752 307628 129804
rect 252468 129684 252520 129736
rect 271236 129684 271288 129736
rect 373356 129684 373408 129736
rect 386604 129684 386656 129736
rect 252376 129616 252428 129668
rect 264428 129616 264480 129668
rect 324320 129004 324372 129056
rect 340788 129004 340840 129056
rect 356704 129004 356756 129056
rect 387064 129004 387116 129056
rect 251732 128460 251784 128512
rect 258908 128460 258960 128512
rect 196716 128392 196768 128444
rect 214012 128392 214064 128444
rect 278136 128392 278188 128444
rect 307484 128392 307536 128444
rect 169024 128324 169076 128376
rect 213920 128324 213972 128376
rect 265624 128324 265676 128376
rect 307668 128324 307720 128376
rect 252468 128256 252520 128308
rect 279608 128256 279660 128308
rect 324320 128256 324372 128308
rect 354772 128256 354824 128308
rect 355968 128256 356020 128308
rect 252376 128188 252428 128240
rect 268568 128188 268620 128240
rect 172336 127576 172388 127628
rect 198096 127576 198148 127628
rect 355968 127576 356020 127628
rect 374736 127576 374788 127628
rect 252100 127168 252152 127220
rect 253296 127168 253348 127220
rect 280804 127100 280856 127152
rect 307668 127100 307720 127152
rect 279516 127032 279568 127084
rect 307484 127032 307536 127084
rect 206468 126964 206520 127016
rect 213920 126964 213972 127016
rect 269764 126964 269816 127016
rect 307576 126964 307628 127016
rect 252376 126896 252428 126948
rect 292028 126896 292080 126948
rect 324320 126896 324372 126948
rect 378140 126896 378192 126948
rect 252468 126828 252520 126880
rect 278228 126828 278280 126880
rect 252468 126556 252520 126608
rect 257528 126556 257580 126608
rect 257712 126216 257764 126268
rect 280896 126216 280948 126268
rect 569224 126216 569276 126268
rect 578332 126216 578384 126268
rect 579620 126216 579672 126268
rect 196808 125672 196860 125724
rect 214012 125672 214064 125724
rect 291936 125672 291988 125724
rect 307576 125672 307628 125724
rect 173440 125604 173492 125656
rect 213920 125604 213972 125656
rect 268476 125604 268528 125656
rect 307668 125604 307720 125656
rect 324320 125536 324372 125588
rect 349252 125536 349304 125588
rect 349620 125536 349672 125588
rect 252468 125468 252520 125520
rect 275284 125468 275336 125520
rect 324412 125468 324464 125520
rect 347872 125468 347924 125520
rect 367836 125468 367888 125520
rect 252376 125400 252428 125452
rect 279700 125400 279752 125452
rect 251180 125332 251232 125384
rect 253480 125332 253532 125384
rect 280160 124924 280212 124976
rect 291844 124924 291896 124976
rect 275376 124856 275428 124908
rect 307024 124856 307076 124908
rect 349620 124856 349672 124908
rect 389824 124856 389876 124908
rect 260380 124380 260432 124432
rect 306748 124380 306800 124432
rect 296076 124312 296128 124364
rect 307484 124312 307536 124364
rect 170496 124244 170548 124296
rect 213920 124244 213972 124296
rect 278228 124244 278280 124296
rect 307668 124244 307720 124296
rect 166356 124176 166408 124228
rect 214012 124176 214064 124228
rect 252284 124108 252336 124160
rect 295984 124108 296036 124160
rect 324504 124108 324556 124160
rect 350632 124108 350684 124160
rect 572628 124108 572680 124160
rect 583300 124108 583352 124160
rect 252468 124040 252520 124092
rect 289268 124040 289320 124092
rect 324320 124040 324372 124092
rect 334072 124040 334124 124092
rect 252376 123972 252428 124024
rect 261484 123972 261536 124024
rect 324412 123972 324464 124024
rect 329196 123972 329248 124024
rect 350632 123428 350684 123480
rect 385868 123428 385920 123480
rect 294604 122952 294656 123004
rect 307116 122952 307168 123004
rect 170588 122884 170640 122936
rect 213920 122884 213972 122936
rect 293224 122884 293276 122936
rect 307668 122884 307720 122936
rect 167736 122816 167788 122868
rect 214012 122816 214064 122868
rect 287796 122816 287848 122868
rect 307484 122816 307536 122868
rect 252468 122748 252520 122800
rect 287704 122748 287756 122800
rect 321652 122748 321704 122800
rect 341524 122748 341576 122800
rect 377404 122748 377456 122800
rect 386788 122748 386840 122800
rect 252376 122680 252428 122732
rect 281080 122680 281132 122732
rect 324320 122476 324372 122528
rect 327080 122476 327132 122528
rect 167920 122068 167972 122120
rect 203616 122068 203668 122120
rect 337476 122068 337528 122120
rect 387156 122068 387208 122120
rect 252468 121864 252520 121916
rect 260104 121864 260156 121916
rect 290464 121592 290516 121644
rect 307668 121592 307720 121644
rect 206560 121524 206612 121576
rect 214012 121524 214064 121576
rect 283748 121524 283800 121576
rect 307576 121524 307628 121576
rect 184296 121456 184348 121508
rect 213920 121456 213972 121508
rect 267004 121456 267056 121508
rect 307484 121456 307536 121508
rect 252376 121388 252428 121440
rect 297548 121388 297600 121440
rect 324320 121388 324372 121440
rect 343732 121388 343784 121440
rect 252468 121320 252520 121372
rect 263140 121320 263192 121372
rect 324412 121320 324464 121372
rect 327540 121320 327592 121372
rect 251548 121252 251600 121304
rect 257436 121252 257488 121304
rect 343732 120708 343784 120760
rect 383108 120708 383160 120760
rect 297640 120232 297692 120284
rect 307576 120232 307628 120284
rect 187056 120164 187108 120216
rect 213920 120164 213972 120216
rect 291844 120164 291896 120216
rect 307668 120164 307720 120216
rect 182916 120096 182968 120148
rect 214012 120096 214064 120148
rect 262956 120096 263008 120148
rect 306748 120096 306800 120148
rect 252376 120028 252428 120080
rect 289084 120028 289136 120080
rect 324320 120028 324372 120080
rect 349344 120028 349396 120080
rect 370596 120028 370648 120080
rect 386880 120028 386932 120080
rect 252468 119960 252520 120012
rect 261576 119960 261628 120012
rect 340236 119960 340288 120012
rect 363604 119960 363656 120012
rect 251732 119348 251784 119400
rect 298744 119348 298796 119400
rect 349344 119348 349396 119400
rect 378968 119348 379020 119400
rect 210608 118804 210660 118856
rect 214104 118804 214156 118856
rect 302976 118804 303028 118856
rect 307668 118804 307720 118856
rect 212172 118736 212224 118788
rect 214012 118736 214064 118788
rect 296168 118736 296220 118788
rect 307116 118736 307168 118788
rect 166448 118668 166500 118720
rect 213920 118668 213972 118720
rect 287704 118668 287756 118720
rect 306564 118668 306616 118720
rect 252376 118600 252428 118652
rect 290648 118600 290700 118652
rect 324412 118600 324464 118652
rect 340236 118600 340288 118652
rect 252468 118532 252520 118584
rect 258816 118532 258868 118584
rect 324320 118532 324372 118584
rect 330576 118532 330628 118584
rect 252100 117920 252152 117972
rect 301596 117920 301648 117972
rect 324504 117920 324556 117972
rect 354680 117920 354732 117972
rect 300124 117444 300176 117496
rect 306564 117444 306616 117496
rect 203616 117376 203668 117428
rect 213920 117376 213972 117428
rect 301780 117376 301832 117428
rect 307668 117376 307720 117428
rect 195336 117308 195388 117360
rect 214012 117308 214064 117360
rect 289268 117308 289320 117360
rect 306932 117308 306984 117360
rect 252468 117240 252520 117292
rect 287980 117240 288032 117292
rect 324320 117240 324372 117292
rect 356060 117240 356112 117292
rect 357348 117240 357400 117292
rect 572628 117240 572680 117292
rect 583208 117240 583260 117292
rect 251824 116560 251876 116612
rect 264336 116560 264388 116612
rect 252008 116356 252060 116408
rect 257620 116356 257672 116408
rect 298744 116084 298796 116136
rect 307576 116084 307628 116136
rect 282276 116016 282328 116068
rect 307668 116016 307720 116068
rect 193956 115948 194008 116000
rect 213920 115948 213972 116000
rect 261576 115948 261628 116000
rect 307484 115948 307536 116000
rect 252008 115880 252060 115932
rect 300216 115880 300268 115932
rect 324412 115880 324464 115932
rect 345112 115880 345164 115932
rect 346308 115880 346360 115932
rect 252284 115812 252336 115864
rect 287888 115812 287940 115864
rect 324780 115200 324832 115252
rect 340144 115200 340196 115252
rect 324320 115064 324372 115116
rect 327724 115064 327776 115116
rect 210424 114588 210476 114640
rect 214012 114588 214064 114640
rect 293316 114588 293368 114640
rect 307484 114588 307536 114640
rect 177396 114520 177448 114572
rect 213920 114520 213972 114572
rect 249156 114520 249208 114572
rect 307116 114520 307168 114572
rect 352564 114520 352616 114572
rect 354680 114520 354732 114572
rect 386880 114520 386932 114572
rect 251548 114452 251600 114504
rect 271420 114452 271472 114504
rect 324412 114452 324464 114504
rect 374000 114452 374052 114504
rect 252468 114384 252520 114436
rect 260288 114384 260340 114436
rect 324320 114384 324372 114436
rect 336740 114384 336792 114436
rect 338028 114384 338080 114436
rect 252192 114316 252244 114368
rect 254860 114316 254912 114368
rect 260104 113772 260156 113824
rect 284300 113772 284352 113824
rect 338028 113772 338080 113824
rect 388536 113772 388588 113824
rect 289084 113296 289136 113348
rect 307668 113296 307720 113348
rect 184388 113228 184440 113280
rect 213920 113228 213972 113280
rect 254584 113228 254636 113280
rect 171968 113160 172020 113212
rect 214012 113160 214064 113212
rect 272524 113228 272576 113280
rect 307576 113228 307628 113280
rect 306564 113160 306616 113212
rect 251548 113092 251600 113144
rect 296260 113092 296312 113144
rect 324320 113092 324372 113144
rect 338120 113092 338172 113144
rect 252468 113024 252520 113076
rect 275376 113024 275428 113076
rect 338120 112480 338172 112532
rect 376116 112480 376168 112532
rect 325056 112412 325108 112464
rect 387156 112412 387208 112464
rect 252376 112208 252428 112260
rect 258724 112208 258776 112260
rect 199384 111868 199436 111920
rect 213920 111868 213972 111920
rect 299020 111868 299072 111920
rect 307576 111868 307628 111920
rect 192668 111800 192720 111852
rect 214012 111800 214064 111852
rect 295984 111800 296036 111852
rect 307668 111800 307720 111852
rect 570604 111800 570656 111852
rect 579896 111800 579948 111852
rect 252468 111732 252520 111784
rect 273996 111732 274048 111784
rect 324320 111732 324372 111784
rect 347780 111732 347832 111784
rect 252376 111664 252428 111716
rect 257344 111664 257396 111716
rect 347780 111052 347832 111104
rect 388720 111052 388772 111104
rect 324412 110712 324464 110764
rect 327080 110712 327132 110764
rect 300216 110576 300268 110628
rect 307668 110576 307720 110628
rect 189908 110508 189960 110560
rect 213920 110508 213972 110560
rect 274088 110508 274140 110560
rect 307484 110508 307536 110560
rect 169208 110440 169260 110492
rect 214012 110440 214064 110492
rect 258724 110440 258776 110492
rect 307576 110440 307628 110492
rect 252376 110372 252428 110424
rect 304356 110372 304408 110424
rect 324320 110372 324372 110424
rect 329932 110372 329984 110424
rect 252468 110304 252520 110356
rect 289360 110304 289412 110356
rect 252100 109964 252152 110016
rect 256056 109964 256108 110016
rect 301596 109148 301648 109200
rect 307668 109148 307720 109200
rect 209044 109080 209096 109132
rect 214012 109080 214064 109132
rect 304540 109080 304592 109132
rect 306932 109080 306984 109132
rect 167920 109012 167972 109064
rect 213920 109012 213972 109064
rect 273996 109012 274048 109064
rect 307576 109012 307628 109064
rect 168104 108944 168156 108996
rect 177488 108944 177540 108996
rect 252468 108944 252520 108996
rect 283932 108944 283984 108996
rect 353944 108944 353996 108996
rect 386604 108944 386656 108996
rect 252376 108876 252428 108928
rect 260196 108876 260248 108928
rect 252100 108672 252152 108724
rect 256148 108672 256200 108724
rect 214748 108400 214800 108452
rect 214656 108196 214708 108248
rect 324320 108332 324372 108384
rect 325792 108332 325844 108384
rect 329196 108332 329248 108384
rect 324412 108264 324464 108316
rect 351276 108264 351328 108316
rect 258816 107856 258868 107908
rect 307668 107856 307720 107908
rect 300308 107788 300360 107840
rect 307576 107788 307628 107840
rect 207848 107720 207900 107772
rect 213920 107720 213972 107772
rect 264244 107720 264296 107772
rect 307392 107720 307444 107772
rect 188528 107652 188580 107704
rect 214012 107652 214064 107704
rect 304448 107652 304500 107704
rect 307484 107652 307536 107704
rect 252468 107584 252520 107636
rect 272616 107584 272668 107636
rect 252376 107516 252428 107568
rect 269856 107516 269908 107568
rect 251548 107040 251600 107092
rect 254676 107040 254728 107092
rect 252468 106904 252520 106956
rect 263048 106904 263100 106956
rect 575388 106904 575440 106956
rect 580356 106904 580408 106956
rect 256056 106428 256108 106480
rect 307668 106428 307720 106480
rect 185676 106360 185728 106412
rect 213920 106360 213972 106412
rect 271420 106360 271472 106412
rect 307576 106360 307628 106412
rect 170680 106292 170732 106344
rect 214012 106292 214064 106344
rect 321560 106292 321612 106344
rect 387248 106292 387300 106344
rect 571248 106292 571300 106344
rect 574836 106292 574888 106344
rect 252100 106224 252152 106276
rect 283840 106224 283892 106276
rect 324320 106224 324372 106276
rect 354680 106224 354732 106276
rect 251640 106156 251692 106208
rect 254768 106156 254820 106208
rect 252008 105544 252060 105596
rect 301504 105544 301556 105596
rect 337384 105544 337436 105596
rect 389732 105544 389784 105596
rect 205088 105000 205140 105052
rect 213920 105000 213972 105052
rect 203708 104932 203760 104984
rect 214012 104932 214064 104984
rect 301688 104932 301740 104984
rect 307576 104932 307628 104984
rect 191196 104864 191248 104916
rect 214104 104864 214156 104916
rect 283656 104864 283708 104916
rect 307668 104864 307720 104916
rect 252100 104796 252152 104848
rect 305736 104796 305788 104848
rect 252284 104388 252336 104440
rect 255964 104388 256016 104440
rect 285128 103640 285180 103692
rect 307484 103640 307536 103692
rect 198280 103572 198332 103624
rect 213920 103572 213972 103624
rect 296260 103572 296312 103624
rect 307668 103572 307720 103624
rect 194048 103504 194100 103556
rect 214012 103504 214064 103556
rect 322940 103504 322992 103556
rect 385960 103504 386012 103556
rect 252468 103436 252520 103488
rect 264520 103436 264572 103488
rect 324412 103436 324464 103488
rect 346400 103436 346452 103488
rect 252376 102756 252428 102808
rect 293408 102756 293460 102808
rect 304356 102280 304408 102332
rect 306748 102280 306800 102332
rect 200764 102212 200816 102264
rect 214012 102212 214064 102264
rect 292028 102212 292080 102264
rect 307484 102212 307536 102264
rect 198188 102144 198240 102196
rect 213920 102144 213972 102196
rect 269856 102144 269908 102196
rect 307668 102144 307720 102196
rect 572628 102144 572680 102196
rect 574192 102144 574244 102196
rect 252100 102076 252152 102128
rect 278320 102076 278372 102128
rect 251824 102008 251876 102060
rect 267096 102008 267148 102060
rect 292672 101396 292724 101448
rect 302240 101396 302292 101448
rect 324596 101396 324648 101448
rect 337476 101396 337528 101448
rect 303068 100920 303120 100972
rect 306748 100920 306800 100972
rect 287888 100852 287940 100904
rect 307484 100852 307536 100904
rect 275376 100784 275428 100836
rect 307668 100784 307720 100836
rect 204996 100716 205048 100768
rect 213920 100716 213972 100768
rect 271236 100716 271288 100768
rect 307576 100716 307628 100768
rect 251916 100648 251968 100700
rect 297732 100648 297784 100700
rect 252100 100580 252152 100632
rect 261760 100580 261812 100632
rect 169300 100036 169352 100088
rect 214656 100036 214708 100088
rect 166540 99968 166592 100020
rect 214380 99968 214432 100020
rect 252284 99968 252336 100020
rect 306012 99968 306064 100020
rect 297548 99356 297600 99408
rect 307484 99356 307536 99408
rect 172428 99288 172480 99340
rect 217968 99288 218020 99340
rect 324320 99288 324372 99340
rect 368480 99288 368532 99340
rect 381636 99288 381688 99340
rect 386880 99288 386932 99340
rect 252376 99220 252428 99272
rect 299112 99220 299164 99272
rect 324412 99220 324464 99272
rect 345020 99220 345072 99272
rect 251180 98948 251232 99000
rect 253204 98948 253256 99000
rect 191104 98676 191156 98728
rect 217324 98676 217376 98728
rect 188344 98608 188396 98660
rect 217416 98608 217468 98660
rect 251916 98608 251968 98660
rect 282368 98608 282420 98660
rect 301504 98132 301556 98184
rect 306564 98132 306616 98184
rect 298836 98064 298888 98116
rect 307576 98064 307628 98116
rect 167828 97996 167880 98048
rect 213920 97996 213972 98048
rect 255964 97996 256016 98048
rect 307668 97996 307720 98048
rect 389640 96772 389692 96824
rect 389824 96772 389876 96824
rect 275284 96704 275336 96756
rect 307668 96704 307720 96756
rect 207940 96636 207992 96688
rect 213920 96636 213972 96688
rect 253296 96636 253348 96688
rect 307484 96636 307536 96688
rect 198096 96568 198148 96620
rect 321744 96568 321796 96620
rect 324320 96568 324372 96620
rect 342352 96568 342404 96620
rect 378876 96568 378928 96620
rect 575572 96568 575624 96620
rect 383016 96500 383068 96552
rect 568580 96500 568632 96552
rect 165528 95888 165580 95940
rect 214012 95888 214064 95940
rect 261484 95888 261536 95940
rect 292580 95888 292632 95940
rect 367928 95412 367980 95464
rect 392584 95412 392636 95464
rect 385776 95344 385828 95396
rect 428004 95344 428056 95396
rect 380256 95276 380308 95328
rect 500776 95276 500828 95328
rect 172060 95208 172112 95260
rect 213920 95208 213972 95260
rect 249064 95208 249116 95260
rect 307668 95208 307720 95260
rect 355324 95208 355376 95260
rect 507216 95208 507268 95260
rect 523316 95208 523368 95260
rect 578240 95208 578292 95260
rect 174544 95140 174596 95192
rect 324688 95140 324740 95192
rect 388720 95140 388772 95192
rect 399024 95140 399076 95192
rect 548432 95140 548484 95192
rect 576124 95140 576176 95192
rect 207664 95072 207716 95124
rect 325700 95072 325752 95124
rect 385684 95072 385736 95124
rect 395804 95072 395856 95124
rect 418344 95072 418396 95124
rect 574744 95072 574796 95124
rect 331956 95004 332008 95056
rect 424784 95004 424836 95056
rect 541992 95004 542044 95056
rect 569224 95004 569276 95056
rect 382924 94936 382976 94988
rect 437020 94936 437072 94988
rect 322940 94868 322992 94920
rect 513656 94868 513708 94920
rect 388628 94800 388680 94852
rect 421564 94800 421616 94852
rect 126888 94460 126940 94512
rect 214104 94460 214156 94512
rect 246304 94460 246356 94512
rect 257712 94460 257764 94512
rect 151912 94052 151964 94104
rect 171784 94052 171836 94104
rect 123208 93984 123260 94036
rect 173348 93984 173400 94036
rect 112352 93916 112404 93968
rect 166448 93916 166500 93968
rect 113180 93848 113232 93900
rect 169116 93848 169168 93900
rect 67640 93780 67692 93832
rect 205088 93780 205140 93832
rect 217416 93780 217468 93832
rect 322940 93848 322992 93900
rect 325700 93848 325752 93900
rect 564532 93780 564584 93832
rect 582932 93780 582984 93832
rect 443460 93712 443512 93764
rect 456340 93712 456392 93764
rect 582380 93712 582432 93764
rect 384304 93644 384356 93696
rect 475660 93644 475712 93696
rect 487804 93644 487856 93696
rect 573364 93644 573416 93696
rect 356796 93576 356848 93628
rect 402244 93576 402296 93628
rect 529756 93576 529808 93628
rect 569316 93576 569368 93628
rect 387156 93508 387208 93560
rect 415124 93508 415176 93560
rect 567752 93508 567804 93560
rect 582840 93508 582892 93560
rect 385868 93440 385920 93492
rect 411904 93440 411956 93492
rect 376024 93372 376076 93424
rect 572720 93372 572772 93424
rect 121736 93304 121788 93356
rect 167736 93304 167788 93356
rect 151544 93236 151596 93288
rect 202236 93236 202288 93288
rect 93952 93168 94004 93220
rect 207848 93168 207900 93220
rect 107752 93100 107804 93152
rect 193956 93100 194008 93152
rect 206376 93100 206428 93152
rect 324320 93100 324372 93152
rect 88984 92420 89036 92472
rect 165528 92420 165580 92472
rect 380348 92420 380400 92472
rect 576860 92420 576912 92472
rect 118056 92352 118108 92404
rect 188436 92352 188488 92404
rect 388444 92352 388496 92404
rect 571432 92352 571484 92404
rect 87236 92284 87288 92336
rect 126888 92284 126940 92336
rect 129464 92284 129516 92336
rect 189816 92284 189868 92336
rect 387708 92284 387760 92336
rect 570604 92284 570656 92336
rect 107476 92216 107528 92268
rect 128360 92216 128412 92268
rect 135720 92216 135772 92268
rect 193864 92216 193916 92268
rect 360844 92216 360896 92268
rect 509884 92216 509936 92268
rect 510528 92216 510580 92268
rect 114192 92148 114244 92200
rect 169300 92148 169352 92200
rect 351184 92148 351236 92200
rect 418344 92148 418396 92200
rect 449900 92148 449952 92200
rect 576216 92148 576268 92200
rect 125784 92080 125836 92132
rect 166540 92080 166592 92132
rect 381544 92080 381596 92132
rect 446680 92080 446732 92132
rect 238024 91876 238076 91928
rect 250996 91876 251048 91928
rect 167000 91808 167052 91860
rect 204904 91808 204956 91860
rect 228364 91808 228416 91860
rect 260380 91808 260432 91860
rect 198740 91740 198792 91792
rect 276112 91740 276164 91792
rect 430488 91740 430540 91792
rect 431224 91740 431276 91792
rect 109684 91128 109736 91180
rect 116676 91128 116728 91180
rect 85764 91060 85816 91112
rect 116584 91060 116636 91112
rect 64788 90992 64840 91044
rect 198280 90992 198332 91044
rect 324320 90992 324372 91044
rect 569960 90992 570012 91044
rect 111616 90924 111668 90976
rect 195336 90924 195388 90976
rect 469220 90924 469272 90976
rect 577504 90924 577556 90976
rect 100484 90856 100536 90908
rect 169208 90856 169260 90908
rect 378784 90856 378836 90908
rect 478880 90856 478932 90908
rect 124496 90788 124548 90840
rect 186964 90788 187016 90840
rect 387248 90788 387300 90840
rect 434444 90788 434496 90840
rect 125416 90720 125468 90772
rect 173440 90720 173492 90772
rect 388536 90720 388588 90772
rect 472440 90720 472492 90772
rect 151728 90652 151780 90704
rect 177304 90652 177356 90704
rect 308404 90312 308456 90364
rect 317420 90312 317472 90364
rect 63316 89632 63368 89684
rect 200764 89632 200816 89684
rect 217324 89632 217376 89684
rect 327080 89632 327132 89684
rect 328368 89632 328420 89684
rect 378968 89632 379020 89684
rect 554872 89632 554924 89684
rect 115388 89564 115440 89616
rect 210608 89564 210660 89616
rect 363696 89564 363748 89616
rect 526536 89564 526588 89616
rect 128176 89496 128228 89548
rect 212080 89496 212132 89548
rect 429200 89496 429252 89548
rect 430488 89496 430540 89548
rect 583852 89496 583904 89548
rect 104256 89428 104308 89480
rect 171968 89428 172020 89480
rect 354036 89428 354088 89480
rect 482100 89428 482152 89480
rect 151360 89360 151412 89412
rect 192484 89360 192536 89412
rect 359464 89360 359516 89412
rect 440240 89360 440292 89412
rect 132224 89292 132276 89344
rect 167000 89292 167052 89344
rect 211896 88952 211948 89004
rect 307300 88952 307352 89004
rect 206284 88272 206336 88324
rect 429200 88272 429252 88324
rect 90732 88204 90784 88256
rect 203708 88204 203760 88256
rect 369216 88204 369268 88256
rect 571616 88204 571668 88256
rect 117136 88136 117188 88188
rect 182916 88136 182968 88188
rect 328368 88136 328420 88188
rect 459560 88136 459612 88188
rect 133144 88068 133196 88120
rect 185584 88068 185636 88120
rect 383108 88068 383160 88120
rect 462780 88068 462832 88120
rect 120724 88000 120776 88052
rect 170588 88000 170640 88052
rect 64696 87932 64748 87984
rect 207940 87932 207992 87984
rect 184204 87592 184256 87644
rect 233884 87592 233936 87644
rect 302884 87592 302936 87644
rect 324504 87592 324556 87644
rect 67732 86912 67784 86964
rect 214840 86912 214892 86964
rect 327908 86912 327960 86964
rect 560300 86912 560352 86964
rect 573456 86912 573508 86964
rect 580172 86912 580224 86964
rect 63408 86844 63460 86896
rect 198188 86844 198240 86896
rect 384396 86844 384448 86896
rect 489920 86844 489972 86896
rect 110144 86776 110196 86828
rect 203616 86776 203668 86828
rect 381728 86776 381780 86828
rect 465080 86776 465132 86828
rect 118240 86708 118292 86760
rect 184296 86708 184348 86760
rect 130752 86640 130804 86692
rect 167644 86640 167696 86692
rect 253204 86300 253256 86352
rect 266360 86300 266412 86352
rect 242900 86232 242952 86284
rect 293960 86232 294012 86284
rect 3148 85484 3200 85536
rect 26884 85484 26936 85536
rect 113916 85484 113968 85536
rect 212172 85484 212224 85536
rect 329196 85484 329248 85536
rect 531320 85484 531372 85536
rect 101864 85416 101916 85468
rect 192668 85416 192720 85468
rect 338764 85416 338816 85468
rect 487804 85416 487856 85468
rect 108488 85348 108540 85400
rect 173256 85348 173308 85400
rect 385960 85348 386012 85400
rect 496820 85348 496872 85400
rect 119896 85280 119948 85332
rect 171876 85280 171928 85332
rect 360936 85280 360988 85332
rect 452660 85280 452712 85332
rect 124036 85212 124088 85264
rect 166356 85212 166408 85264
rect 134708 85144 134760 85196
rect 166264 85144 166316 85196
rect 176384 84804 176436 84856
rect 267740 84804 267792 84856
rect 510528 84804 510580 84856
rect 522304 84804 522356 84856
rect 99104 84124 99156 84176
rect 206468 84124 206520 84176
rect 359556 84124 359608 84176
rect 557540 84124 557592 84176
rect 107568 84056 107620 84108
rect 210424 84056 210476 84108
rect 374736 84056 374788 84108
rect 516140 84056 516192 84108
rect 96528 83988 96580 84040
rect 167920 83988 167972 84040
rect 115848 83920 115900 83972
rect 187056 83920 187108 83972
rect 124128 83852 124180 83904
rect 170496 83852 170548 83904
rect 212540 83444 212592 83496
rect 327080 83444 327132 83496
rect 67272 82764 67324 82816
rect 324412 82764 324464 82816
rect 358084 82764 358136 82816
rect 548524 82764 548576 82816
rect 97908 82696 97960 82748
rect 209044 82696 209096 82748
rect 367744 82696 367796 82748
rect 503720 82696 503772 82748
rect 111708 82628 111760 82680
rect 207756 82628 207808 82680
rect 377496 82628 377548 82680
rect 494060 82628 494112 82680
rect 103336 82560 103388 82612
rect 184388 82560 184440 82612
rect 46848 81336 46900 81388
rect 321560 81336 321612 81388
rect 582748 81336 582800 81388
rect 92388 81268 92440 81320
rect 185676 81268 185728 81320
rect 333888 81268 333940 81320
rect 518900 81268 518952 81320
rect 126888 81200 126940 81252
rect 210516 81200 210568 81252
rect 373448 81200 373500 81252
rect 550640 81200 550692 81252
rect 126796 81132 126848 81184
rect 196808 81132 196860 81184
rect 210424 80656 210476 80708
rect 307208 80656 307260 80708
rect 95148 79976 95200 80028
rect 188528 79976 188580 80028
rect 324964 79976 325016 80028
rect 570144 79976 570196 80028
rect 121368 79908 121420 79960
rect 211988 79908 212040 79960
rect 365076 79908 365128 79960
rect 574192 79908 574244 79960
rect 119988 79840 120040 79892
rect 206560 79840 206612 79892
rect 86868 79772 86920 79824
rect 167828 79772 167880 79824
rect 99196 79704 99248 79756
rect 169024 79704 169076 79756
rect 238760 79364 238812 79416
rect 294052 79364 294104 79416
rect 179328 79296 179380 79348
rect 245660 79296 245712 79348
rect 297456 79296 297508 79348
rect 320180 79296 320232 79348
rect 116676 78616 116728 78668
rect 213184 78616 213236 78668
rect 276664 78616 276716 78668
rect 570052 78616 570104 78668
rect 102048 78548 102100 78600
rect 196716 78548 196768 78600
rect 99288 78480 99340 78532
rect 189908 78480 189960 78532
rect 122748 78412 122800 78464
rect 202144 78412 202196 78464
rect 93768 78344 93820 78396
rect 170680 78344 170732 78396
rect 257988 78004 258040 78056
rect 275468 78004 275520 78056
rect 200120 77936 200172 77988
rect 311900 77936 311952 77988
rect 66904 77188 66956 77240
rect 484400 77188 484452 77240
rect 75828 77120 75880 77172
rect 172060 77120 172112 77172
rect 347044 77120 347096 77172
rect 545120 77120 545172 77172
rect 106188 77052 106240 77104
rect 177396 77052 177448 77104
rect 120080 76508 120132 76560
rect 250536 76508 250588 76560
rect 100576 75828 100628 75880
rect 199384 75828 199436 75880
rect 113088 75760 113140 75812
rect 170404 75760 170456 75812
rect 175096 75216 175148 75268
rect 331312 75216 331364 75268
rect 49700 75148 49752 75200
rect 265716 75148 265768 75200
rect 116584 74468 116636 74520
rect 214564 74468 214616 74520
rect 104808 74400 104860 74452
rect 192576 74400 192628 74452
rect 52460 73856 52512 73908
rect 301780 73856 301832 73908
rect 27620 73788 27672 73840
rect 279516 73788 279568 73840
rect 85488 73108 85540 73160
rect 204996 73108 205048 73160
rect 574836 73108 574888 73160
rect 579988 73108 580040 73160
rect 114560 72496 114612 72548
rect 274088 72496 274140 72548
rect 66260 72428 66312 72480
rect 296168 72428 296220 72480
rect 3424 71680 3476 71732
rect 32404 71680 32456 71732
rect 179144 71136 179196 71188
rect 296720 71136 296772 71188
rect 103520 71068 103572 71120
rect 304540 71068 304592 71120
rect 30380 71000 30432 71052
rect 249156 71000 249208 71052
rect 124220 69708 124272 69760
rect 253388 69708 253440 69760
rect 89720 69640 89772 69692
rect 304448 69640 304500 69692
rect 184940 68416 184992 68468
rect 316132 68416 316184 68468
rect 93860 68348 93912 68400
rect 264244 68348 264296 68400
rect 62120 68280 62172 68332
rect 289268 68280 289320 68332
rect 96620 66852 96672 66904
rect 273996 66852 274048 66904
rect 80060 65560 80112 65612
rect 297640 65560 297692 65612
rect 45560 65492 45612 65544
rect 298928 65492 298980 65544
rect 60740 64132 60792 64184
rect 286416 64132 286468 64184
rect 63500 62840 63552 62892
rect 290556 62840 290608 62892
rect 46940 62772 46992 62824
rect 304356 62772 304408 62824
rect 70400 61412 70452 61464
rect 289176 61412 289228 61464
rect 51080 61344 51132 61396
rect 305920 61344 305972 61396
rect 387616 60664 387668 60716
rect 580172 60664 580224 60716
rect 53840 59984 53892 60036
rect 296260 59984 296312 60036
rect 3056 59304 3108 59356
rect 373264 59304 373316 59356
rect 74540 58624 74592 58676
rect 280988 58624 281040 58676
rect 81440 57264 81492 57316
rect 271328 57264 271380 57316
rect 57980 57196 58032 57248
rect 285128 57196 285180 57248
rect 85580 55904 85632 55956
rect 282184 55904 282236 55956
rect 64880 55836 64932 55888
rect 301688 55836 301740 55888
rect 52552 54476 52604 54528
rect 303160 54476 303212 54528
rect 121460 53116 121512 53168
rect 299020 53116 299072 53168
rect 9680 53048 9732 53100
rect 291936 53048 291988 53100
rect 110420 51756 110472 51808
rect 300216 51756 300268 51808
rect 44180 51688 44232 51740
rect 261576 51688 261628 51740
rect 85672 50396 85724 50448
rect 258816 50396 258868 50448
rect 34520 50328 34572 50380
rect 293316 50328 293368 50380
rect 82820 49036 82872 49088
rect 300308 49036 300360 49088
rect 37280 48968 37332 49020
rect 307116 48968 307168 49020
rect 49608 48220 49660 48272
rect 249248 48220 249300 48272
rect 48964 47880 49016 47932
rect 49608 47880 49660 47932
rect 179604 47540 179656 47592
rect 306380 47540 306432 47592
rect 88340 46180 88392 46232
rect 304264 46180 304316 46232
rect 3424 45500 3476 45552
rect 40684 45500 40736 45552
rect 78680 44888 78732 44940
rect 305828 44888 305880 44940
rect 41420 44820 41472 44872
rect 282276 44820 282328 44872
rect 187700 43596 187752 43648
rect 258816 43596 258868 43648
rect 201500 43528 201552 43580
rect 333244 43528 333296 43580
rect 4160 43460 4212 43512
rect 249064 43460 249116 43512
rect 44272 43392 44324 43444
rect 292028 43392 292080 43444
rect 104900 42100 104952 42152
rect 287796 42100 287848 42152
rect 75920 42032 75972 42084
rect 271420 42032 271472 42084
rect 122840 40672 122892 40724
rect 268476 40672 268528 40724
rect 107660 39380 107712 39432
rect 258724 39380 258776 39432
rect 77300 39312 77352 39364
rect 291844 39312 291896 39364
rect 179512 38020 179564 38072
rect 293960 38020 294012 38072
rect 93952 37952 94004 38004
rect 267004 37952 267056 38004
rect 42800 37884 42852 37936
rect 286324 37884 286376 37936
rect 16580 36524 16632 36576
rect 297548 36524 297600 36576
rect 177948 35300 178000 35352
rect 298928 35300 298980 35352
rect 27712 35232 27764 35284
rect 272524 35232 272576 35284
rect 20720 35164 20772 35216
rect 305736 35164 305788 35216
rect 179420 33872 179472 33924
rect 332692 33872 332744 33924
rect 71780 33804 71832 33856
rect 256056 33804 256108 33856
rect 98000 33736 98052 33788
rect 294604 33736 294656 33788
rect 3516 33056 3568 33108
rect 13084 33056 13136 33108
rect 522304 33056 522356 33108
rect 580172 33056 580224 33108
rect 208400 32512 208452 32564
rect 323584 32512 323636 32564
rect 106280 32444 106332 32496
rect 250444 32444 250496 32496
rect 48320 32376 48372 32428
rect 298744 32376 298796 32428
rect 73160 31084 73212 31136
rect 302976 31084 303028 31136
rect 33140 31016 33192 31068
rect 287888 31016 287940 31068
rect 176568 29724 176620 29776
rect 262220 29724 262272 29776
rect 118700 29656 118752 29708
rect 228364 29656 228416 29708
rect 12440 29588 12492 29640
rect 289084 29588 289136 29640
rect 102140 28296 102192 28348
rect 293224 28296 293276 28348
rect 26240 28228 26292 28280
rect 275376 28228 275428 28280
rect 100760 26868 100812 26920
rect 301596 26868 301648 26920
rect 91100 25576 91152 25628
rect 283748 25576 283800 25628
rect 24860 25508 24912 25560
rect 298836 25508 298888 25560
rect 193220 24216 193272 24268
rect 242164 24216 242216 24268
rect 56600 24148 56652 24200
rect 262864 24148 262916 24200
rect 2872 24080 2924 24132
rect 275284 24080 275336 24132
rect 86960 22788 87012 22840
rect 290464 22788 290516 22840
rect 19340 22720 19392 22772
rect 255964 22720 256016 22772
rect 179236 21496 179288 21548
rect 284300 21496 284352 21548
rect 40040 21428 40092 21480
rect 269856 21428 269908 21480
rect 15200 21360 15252 21412
rect 307024 21360 307076 21412
rect 3424 20612 3476 20664
rect 22836 20612 22888 20664
rect 195244 20068 195296 20120
rect 273260 20068 273312 20120
rect 115940 20000 115992 20052
rect 296076 20000 296128 20052
rect 38660 19932 38712 19984
rect 278136 19932 278188 19984
rect 109040 18640 109092 18692
rect 278228 18640 278280 18692
rect 11152 18572 11204 18624
rect 253296 18572 253348 18624
rect 110512 17280 110564 17332
rect 279424 17280 279476 17332
rect 23480 17212 23532 17264
rect 280804 17212 280856 17264
rect 175188 15920 175240 15972
rect 311440 15920 311492 15972
rect 84200 15852 84252 15904
rect 262956 15852 263008 15904
rect 135260 14492 135312 14544
rect 203524 14492 203576 14544
rect 233884 14492 233936 14544
rect 281540 14492 281592 14544
rect 36728 14424 36780 14476
rect 303068 14424 303120 14476
rect 183560 13200 183612 13252
rect 349252 13200 349304 13252
rect 22560 13132 22612 13184
rect 254584 13132 254636 13184
rect 59360 13064 59412 13116
rect 300124 13064 300176 13116
rect 128912 11840 128964 11892
rect 216680 11840 216732 11892
rect 112352 11772 112404 11824
rect 305644 11772 305696 11824
rect 30104 11704 30156 11756
rect 271236 11704 271288 11756
rect 112 10956 164 11008
rect 1308 10956 1360 11008
rect 251180 10956 251232 11008
rect 176476 10344 176528 10396
rect 299480 10344 299532 10396
rect 92480 10276 92532 10328
rect 283564 10276 283616 10328
rect 189724 9052 189776 9104
rect 245200 9052 245252 9104
rect 96252 8984 96304 9036
rect 285036 8984 285088 9036
rect 1676 8916 1728 8968
rect 48964 8916 49016 8968
rect 62028 8916 62080 8968
rect 283656 8916 283708 8968
rect 99840 7624 99892 7676
rect 273904 7624 273956 7676
rect 7656 7556 7708 7608
rect 301504 7556 301556 7608
rect 3424 6808 3476 6860
rect 35164 6808 35216 6860
rect 180800 6332 180852 6384
rect 268844 6332 268896 6384
rect 211804 6264 211856 6316
rect 305552 6264 305604 6316
rect 309048 6264 309100 6316
rect 335452 6264 335504 6316
rect 182824 6196 182876 6248
rect 348056 6196 348108 6248
rect 70308 6128 70360 6180
rect 287704 6128 287756 6180
rect 303160 6128 303212 6180
rect 332600 6128 332652 6180
rect 198004 4836 198056 4888
rect 260656 4836 260708 4888
rect 35992 4768 36044 4820
rect 265624 4768 265676 4820
rect 216128 3680 216180 3732
rect 240508 3680 240560 3732
rect 242164 3680 242216 3732
rect 247592 3680 247644 3732
rect 253480 3680 253532 3732
rect 261484 3680 261536 3732
rect 114008 3612 114060 3664
rect 110420 3544 110472 3596
rect 111616 3544 111668 3596
rect 118700 3544 118752 3596
rect 119896 3544 119948 3596
rect 211068 3612 211120 3664
rect 248788 3612 248840 3664
rect 210424 3544 210476 3596
rect 216036 3544 216088 3596
rect 254676 3612 254728 3664
rect 268384 3612 268436 3664
rect 251088 3544 251140 3596
rect 252376 3544 252428 3596
rect 257988 3544 258040 3596
rect 264152 3544 264204 3596
rect 276020 3544 276072 3596
rect 276756 3544 276808 3596
rect 284944 3612 284996 3664
rect 298468 3612 298520 3664
rect 288992 3544 289044 3596
rect 299572 3544 299624 3596
rect 300768 3544 300820 3596
rect 319720 3544 319772 3596
rect 331220 3544 331272 3596
rect 331864 3544 331916 3596
rect 333888 3544 333940 3596
rect 11060 3476 11112 3528
rect 11980 3476 12032 3528
rect 27620 3476 27672 3528
rect 28540 3476 28592 3528
rect 44180 3476 44232 3528
rect 45100 3476 45152 3528
rect 103336 3476 103388 3528
rect 211896 3476 211948 3528
rect 215944 3476 215996 3528
rect 6460 3408 6512 3460
rect 192484 3408 192536 3460
rect 196624 3408 196676 3460
rect 135260 3340 135312 3392
rect 136456 3340 136508 3392
rect 235816 3340 235868 3392
rect 238024 3340 238076 3392
rect 242900 3340 242952 3392
rect 244096 3340 244148 3392
rect 249984 3340 250036 3392
rect 253204 3340 253256 3392
rect 241704 3272 241756 3324
rect 246304 3272 246356 3324
rect 258816 3476 258868 3528
rect 261760 3476 261812 3528
rect 271144 3476 271196 3528
rect 326804 3476 326856 3528
rect 329104 3476 329156 3528
rect 330392 3476 330444 3528
rect 333244 3476 333296 3528
rect 344560 3476 344612 3528
rect 349160 3476 349212 3528
rect 350448 3476 350500 3528
rect 266544 3340 266596 3392
rect 292580 3408 292632 3460
rect 298928 3408 298980 3460
rect 301964 3408 302016 3460
rect 297364 3340 297416 3392
rect 322112 3408 322164 3460
rect 323308 3408 323360 3460
rect 340880 3408 340932 3460
rect 342168 3408 342220 3460
rect 343640 3408 343692 3460
rect 309784 3340 309836 3392
rect 317328 3340 317380 3392
rect 323584 3340 323636 3392
rect 325608 3340 325660 3392
rect 309876 3272 309928 3324
rect 315028 3272 315080 3324
rect 258264 3000 258316 3052
rect 260104 3000 260156 3052
rect 308496 2932 308548 2984
rect 310244 2932 310296 2984
rect 346952 2932 347004 2984
rect 351920 2932 351972 2984
rect 278044 2864 278096 2916
rect 283104 2864 283156 2916
rect 118792 2116 118844 2168
rect 295984 2116 296036 2168
rect 19432 2048 19484 2100
rect 269764 2048 269816 2100
<< obsm1 >>
rect 68800 95100 164756 174600
<< metal2 >>
rect 6932 703582 7972 703610
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 684214 3464 684247
rect 3424 684208 3476 684214
rect 3424 684150 3476 684156
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 6932 670002 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 24320 699718 24348 703520
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 25504 699712 25556 699718
rect 25504 699654 25556 699660
rect 8944 684208 8996 684214
rect 8944 684150 8996 684156
rect 6920 669996 6972 670002
rect 6920 669938 6972 669944
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 553450 3464 553823
rect 3424 553444 3476 553450
rect 3424 553386 3476 553392
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 527202 3464 527847
rect 3424 527196 3476 527202
rect 3424 527138 3476 527144
rect 3422 514856 3478 514865
rect 3422 514791 3424 514800
rect 3476 514791 3478 514800
rect 3424 514762 3476 514768
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3436 474774 3464 475623
rect 3424 474768 3476 474774
rect 3424 474710 3476 474716
rect 3238 462632 3294 462641
rect 3238 462567 3294 462576
rect 3252 462398 3280 462567
rect 3240 462392 3292 462398
rect 3240 462334 3292 462340
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 3422 423600 3478 423609
rect 3422 423535 3478 423544
rect 3436 422346 3464 423535
rect 3424 422340 3476 422346
rect 3424 422282 3476 422288
rect 3146 410544 3202 410553
rect 3146 410479 3202 410488
rect 3160 409902 3188 410479
rect 3148 409896 3200 409902
rect 3148 409838 3200 409844
rect 3424 397520 3476 397526
rect 3422 397488 3424 397497
rect 3476 397488 3478 397497
rect 3422 397423 3478 397432
rect 3422 371376 3478 371385
rect 3422 371311 3478 371320
rect 3436 371278 3464 371311
rect 3424 371272 3476 371278
rect 3424 371214 3476 371220
rect 8956 370530 8984 684150
rect 22744 618316 22796 618322
rect 22744 618258 22796 618264
rect 13084 422340 13136 422346
rect 13084 422282 13136 422288
rect 8944 370524 8996 370530
rect 8944 370466 8996 370472
rect 3422 358456 3478 358465
rect 3422 358391 3478 358400
rect 3436 324970 3464 358391
rect 3514 345400 3570 345409
rect 3514 345335 3570 345344
rect 3528 345234 3556 345335
rect 3516 345228 3568 345234
rect 3516 345170 3568 345176
rect 8944 345228 8996 345234
rect 8944 345170 8996 345176
rect 3424 324964 3476 324970
rect 3424 324906 3476 324912
rect 3422 319288 3478 319297
rect 3422 319223 3478 319232
rect 3436 318850 3464 319223
rect 3424 318844 3476 318850
rect 3424 318786 3476 318792
rect 8956 311166 8984 345170
rect 8944 311160 8996 311166
rect 8944 311102 8996 311108
rect 3238 306232 3294 306241
rect 3238 306167 3294 306176
rect 3252 305046 3280 306167
rect 3240 305040 3292 305046
rect 3240 304982 3292 304988
rect 13096 304978 13124 422282
rect 13084 304972 13136 304978
rect 13084 304914 13136 304920
rect 3422 293176 3478 293185
rect 3422 293111 3478 293120
rect 3436 292602 3464 293111
rect 3424 292596 3476 292602
rect 3424 292538 3476 292544
rect 4068 289128 4120 289134
rect 4068 289070 4120 289076
rect 3054 267200 3110 267209
rect 3054 267135 3110 267144
rect 3068 266422 3096 267135
rect 3056 266416 3108 266422
rect 3056 266358 3108 266364
rect 2778 254144 2834 254153
rect 2778 254079 2780 254088
rect 2832 254079 2834 254088
rect 2780 254050 2832 254056
rect 3422 241088 3478 241097
rect 3422 241023 3478 241032
rect 3436 240174 3464 241023
rect 3424 240168 3476 240174
rect 3424 240110 3476 240116
rect 1308 232552 1360 232558
rect 1308 232494 1360 232500
rect 1320 11014 1348 232494
rect 3424 221468 3476 221474
rect 3424 221410 3476 221416
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3436 201929 3464 221410
rect 3422 201920 3478 201929
rect 3422 201855 3478 201864
rect 3424 189032 3476 189038
rect 3424 188974 3476 188980
rect 3436 188873 3464 188974
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 4080 163538 4108 289070
rect 22756 273970 22784 618258
rect 25516 307086 25544 699654
rect 32404 656940 32456 656946
rect 32404 656882 32456 656888
rect 31024 474768 31076 474774
rect 31024 474710 31076 474716
rect 31036 369170 31064 474710
rect 31024 369164 31076 369170
rect 31024 369106 31076 369112
rect 32416 366382 32444 656882
rect 36544 553444 36596 553450
rect 36544 553386 36596 553392
rect 32404 366376 32456 366382
rect 32404 366318 32456 366324
rect 25504 307080 25556 307086
rect 25504 307022 25556 307028
rect 22836 299532 22888 299538
rect 22836 299474 22888 299480
rect 22744 273964 22796 273970
rect 22744 273906 22796 273912
rect 13084 267776 13136 267782
rect 13084 267718 13136 267724
rect 4804 254108 4856 254114
rect 4804 254050 4856 254056
rect 4816 235890 4844 254050
rect 4804 235884 4856 235890
rect 4804 235826 4856 235832
rect 7564 228404 7616 228410
rect 7564 228346 7616 228352
rect 4804 175976 4856 175982
rect 4804 175918 4856 175924
rect 3700 163532 3752 163538
rect 3700 163474 3752 163480
rect 4068 163532 4120 163538
rect 4068 163474 4120 163480
rect 3712 162897 3740 163474
rect 3698 162888 3754 162897
rect 3698 162823 3754 162832
rect 3424 150408 3476 150414
rect 3424 150350 3476 150356
rect 3436 149841 3464 150350
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3240 137964 3292 137970
rect 3240 137906 3292 137912
rect 3252 136785 3280 137906
rect 3238 136776 3294 136785
rect 3238 136711 3294 136720
rect 4816 110770 4844 175918
rect 2780 110764 2832 110770
rect 2780 110706 2832 110712
rect 4804 110764 4856 110770
rect 4804 110706 4856 110712
rect 2792 110673 2820 110706
rect 2778 110664 2834 110673
rect 2778 110599 2834 110608
rect 7576 97646 7604 228346
rect 3424 97640 3476 97646
rect 3422 97608 3424 97617
rect 7564 97640 7616 97646
rect 3476 97608 3478 97617
rect 7564 97582 7616 97588
rect 3422 97543 3478 97552
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 2778 64152 2834 64161
rect 2778 64087 2834 64096
rect 112 11008 164 11014
rect 112 10950 164 10956
rect 1308 11008 1360 11014
rect 1308 10950 1360 10956
rect 124 354 152 10950
rect 1676 8968 1728 8974
rect 1676 8910 1728 8916
rect 1688 480 1716 8910
rect 2792 6914 2820 64087
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 9680 53100 9732 53106
rect 9680 53042 9732 53048
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 4160 43512 4212 43518
rect 4160 43454 4212 43460
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 2872 24132 2924 24138
rect 2872 24074 2924 24080
rect 2884 16574 2912 24074
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 4172 16574 4200 43454
rect 8298 40624 8354 40633
rect 8298 40559 8354 40568
rect 8312 16574 8340 40559
rect 2884 16546 3648 16574
rect 4172 16546 5304 16574
rect 8312 16546 8800 16574
rect 2792 6886 2912 6914
rect 2884 480 2912 6886
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 542 354 654 480
rect 124 326 654 354
rect 542 -960 654 326
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3620 354 3648 16546
rect 5276 480 5304 16546
rect 7656 7608 7708 7614
rect 7656 7550 7708 7556
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 6472 480 6500 3402
rect 7668 480 7696 7550
rect 8772 480 8800 16546
rect 4038 354 4150 480
rect 3620 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 53042
rect 11058 46200 11114 46209
rect 11058 46135 11114 46144
rect 11072 3534 11100 46135
rect 13096 33114 13124 267718
rect 21364 263628 21416 263634
rect 21364 263570 21416 263576
rect 17224 257372 17276 257378
rect 17224 257314 17276 257320
rect 14464 240168 14516 240174
rect 14464 240110 14516 240116
rect 14476 237386 14504 240110
rect 14464 237380 14516 237386
rect 14464 237322 14516 237328
rect 17236 137970 17264 257314
rect 21376 215286 21404 263570
rect 21364 215280 21416 215286
rect 21364 215222 21416 215228
rect 17224 137964 17276 137970
rect 17224 137906 17276 137912
rect 17958 75168 18014 75177
rect 17958 75103 18014 75112
rect 13818 66872 13874 66881
rect 13818 66807 13874 66816
rect 13084 33108 13136 33114
rect 13084 33050 13136 33056
rect 12440 29640 12492 29646
rect 12440 29582 12492 29588
rect 11152 18624 11204 18630
rect 11152 18566 11204 18572
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 11164 480 11192 18566
rect 12452 16574 12480 29582
rect 13832 16574 13860 66807
rect 16580 36576 16632 36582
rect 16580 36518 16632 36524
rect 15200 21412 15252 21418
rect 15200 21354 15252 21360
rect 15212 16574 15240 21354
rect 16592 16574 16620 36518
rect 12452 16546 13584 16574
rect 13832 16546 14320 16574
rect 15212 16546 15976 16574
rect 16592 16546 17080 16574
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 11992 354 12020 3470
rect 13556 480 13584 16546
rect 12318 354 12430 480
rect 11992 326 12430 354
rect 12318 -960 12430 326
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 15948 480 15976 16546
rect 17052 480 17080 16546
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 75103
rect 20720 35216 20772 35222
rect 20720 35158 20772 35164
rect 19340 22772 19392 22778
rect 19340 22714 19392 22720
rect 19352 16574 19380 22714
rect 20732 16574 20760 35158
rect 22848 20670 22876 299474
rect 32404 295452 32456 295458
rect 32404 295394 32456 295400
rect 31024 290488 31076 290494
rect 31024 290430 31076 290436
rect 25504 266416 25556 266422
rect 25504 266358 25556 266364
rect 25516 238746 25544 266358
rect 26884 253224 26936 253230
rect 26884 253166 26936 253172
rect 25504 238740 25556 238746
rect 25504 238682 25556 238688
rect 26896 85542 26924 253166
rect 31036 150414 31064 290430
rect 31024 150408 31076 150414
rect 31024 150350 31076 150356
rect 26884 85536 26936 85542
rect 26884 85478 26936 85484
rect 27620 73840 27672 73846
rect 27620 73782 27672 73788
rect 26240 28280 26292 28286
rect 26240 28222 26292 28228
rect 24860 25560 24912 25566
rect 24860 25502 24912 25508
rect 22836 20664 22888 20670
rect 22836 20606 22888 20612
rect 23480 17264 23532 17270
rect 23480 17206 23532 17212
rect 23492 16574 23520 17206
rect 24872 16574 24900 25502
rect 19352 16546 20208 16574
rect 20732 16546 21864 16574
rect 23492 16546 24256 16574
rect 24872 16546 25360 16574
rect 19432 2100 19484 2106
rect 19432 2042 19484 2048
rect 19444 480 19472 2042
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20180 354 20208 16546
rect 21836 480 21864 16546
rect 22560 13184 22612 13190
rect 22560 13126 22612 13132
rect 20598 354 20710 480
rect 20180 326 20710 354
rect 20598 -960 20710 326
rect 21794 -960 21906 480
rect 22572 354 22600 13126
rect 24228 480 24256 16546
rect 25332 480 25360 16546
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 28222
rect 27632 3534 27660 73782
rect 32416 71738 32444 295394
rect 35808 278792 35860 278798
rect 35808 278734 35860 278740
rect 35820 239465 35848 278734
rect 36556 262886 36584 553386
rect 39304 527196 39356 527202
rect 39304 527138 39356 527144
rect 39316 368490 39344 527138
rect 39304 368484 39356 368490
rect 39304 368426 39356 368432
rect 39948 368484 40000 368490
rect 39948 368426 40000 368432
rect 39960 367198 39988 368426
rect 39948 367192 40000 367198
rect 39948 367134 40000 367140
rect 36544 262880 36596 262886
rect 36544 262822 36596 262828
rect 39960 260846 39988 367134
rect 40052 356726 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 700330 73016 703520
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 72976 700324 73028 700330
rect 72976 700266 73028 700272
rect 66904 670744 66956 670750
rect 66904 670686 66956 670692
rect 62764 669996 62816 670002
rect 62764 669938 62816 669944
rect 44824 632120 44876 632126
rect 44824 632062 44876 632068
rect 40040 356720 40092 356726
rect 40040 356662 40092 356668
rect 44836 354006 44864 632062
rect 57244 565888 57296 565894
rect 57244 565830 57296 565836
rect 48964 514820 49016 514826
rect 48964 514762 49016 514768
rect 48976 381546 49004 514762
rect 53104 448588 53156 448594
rect 53104 448530 53156 448536
rect 50344 409896 50396 409902
rect 50344 409838 50396 409844
rect 48964 381540 49016 381546
rect 48964 381482 49016 381488
rect 44824 354000 44876 354006
rect 44824 353942 44876 353948
rect 45468 354000 45520 354006
rect 45468 353942 45520 353948
rect 41328 285728 41380 285734
rect 41328 285670 41380 285676
rect 39948 260840 40000 260846
rect 39948 260782 40000 260788
rect 35162 239456 35218 239465
rect 35162 239391 35218 239400
rect 35806 239456 35862 239465
rect 35806 239391 35862 239400
rect 32404 71732 32456 71738
rect 32404 71674 32456 71680
rect 30380 71052 30432 71058
rect 30380 70994 30432 71000
rect 27712 35284 27764 35290
rect 27712 35226 27764 35232
rect 27620 3528 27672 3534
rect 27620 3470 27672 3476
rect 27724 480 27752 35226
rect 30392 16574 30420 70994
rect 34520 50380 34572 50386
rect 34520 50322 34572 50328
rect 33140 31068 33192 31074
rect 33140 31010 33192 31016
rect 33152 16574 33180 31010
rect 30392 16546 30880 16574
rect 33152 16546 33640 16574
rect 30104 11756 30156 11762
rect 30104 11698 30156 11704
rect 28540 3528 28592 3534
rect 28540 3470 28592 3476
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28552 354 28580 3470
rect 30116 480 30144 11698
rect 28878 354 28990 480
rect 28552 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 32402 4856 32458 4865
rect 32402 4791 32458 4800
rect 32416 480 32444 4791
rect 33612 480 33640 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31270 -960 31382 326
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34532 354 34560 50322
rect 35176 6866 35204 239391
rect 40684 189848 40736 189854
rect 40684 189790 40736 189796
rect 37280 49020 37332 49026
rect 37280 48962 37332 48968
rect 37292 16574 37320 48962
rect 40696 45558 40724 189790
rect 41340 183025 41368 285670
rect 45376 282940 45428 282946
rect 45376 282882 45428 282888
rect 45388 222154 45416 282882
rect 45480 265674 45508 353942
rect 49608 294024 49660 294030
rect 49608 293966 49660 293972
rect 46204 292596 46256 292602
rect 46204 292538 46256 292544
rect 45468 265668 45520 265674
rect 45468 265610 45520 265616
rect 46216 243001 46244 292538
rect 48228 276072 48280 276078
rect 48228 276014 48280 276020
rect 46848 270564 46900 270570
rect 46848 270506 46900 270512
rect 46202 242992 46258 243001
rect 46202 242927 46258 242936
rect 45376 222148 45428 222154
rect 45376 222090 45428 222096
rect 41326 183016 41382 183025
rect 41326 182951 41382 182960
rect 46860 81394 46888 270506
rect 48136 264988 48188 264994
rect 48136 264930 48188 264936
rect 48148 227118 48176 264930
rect 48136 227112 48188 227118
rect 48136 227054 48188 227060
rect 48240 226302 48268 276014
rect 49516 269136 49568 269142
rect 49516 269078 49568 269084
rect 48228 226296 48280 226302
rect 48228 226238 48280 226244
rect 49528 209166 49556 269078
rect 49516 209160 49568 209166
rect 49516 209102 49568 209108
rect 46848 81388 46900 81394
rect 46848 81330 46900 81336
rect 45560 65544 45612 65550
rect 45560 65486 45612 65492
rect 44180 51740 44232 51746
rect 44180 51682 44232 51688
rect 40684 45552 40736 45558
rect 40684 45494 40736 45500
rect 41420 44872 41472 44878
rect 41420 44814 41472 44820
rect 40040 21480 40092 21486
rect 40040 21422 40092 21428
rect 38660 19984 38712 19990
rect 38660 19926 38712 19932
rect 38672 16574 38700 19926
rect 40052 16574 40080 21422
rect 41432 16574 41460 44814
rect 42800 37936 42852 37942
rect 42800 37878 42852 37884
rect 37292 16546 38424 16574
rect 38672 16546 39160 16574
rect 40052 16546 40264 16574
rect 41432 16546 41920 16574
rect 36728 14476 36780 14482
rect 36728 14418 36780 14424
rect 35164 6860 35216 6866
rect 35164 6802 35216 6808
rect 35992 4820 36044 4826
rect 35992 4762 36044 4768
rect 36004 480 36032 4762
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 14418
rect 38396 480 38424 16546
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 41892 480 41920 16546
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 42812 354 42840 37878
rect 44192 3534 44220 51682
rect 44272 43444 44324 43450
rect 44272 43386 44324 43392
rect 44180 3528 44232 3534
rect 44180 3470 44232 3476
rect 44284 480 44312 43386
rect 45572 16574 45600 65486
rect 46940 62824 46992 62830
rect 46940 62766 46992 62772
rect 46952 16574 46980 62766
rect 49620 48278 49648 293966
rect 50356 245614 50384 409838
rect 53116 372638 53144 448530
rect 55036 378820 55088 378826
rect 55036 378762 55088 378768
rect 53104 372632 53156 372638
rect 53104 372574 53156 372580
rect 53748 372632 53800 372638
rect 53748 372574 53800 372580
rect 53760 300150 53788 372574
rect 53748 300144 53800 300150
rect 53748 300086 53800 300092
rect 53656 292732 53708 292738
rect 53656 292674 53708 292680
rect 53104 292664 53156 292670
rect 53104 292606 53156 292612
rect 52368 288516 52420 288522
rect 52368 288458 52420 288464
rect 50988 288448 51040 288454
rect 50988 288390 51040 288396
rect 50896 263696 50948 263702
rect 50896 263638 50948 263644
rect 50344 245608 50396 245614
rect 50344 245550 50396 245556
rect 50908 220114 50936 263638
rect 50896 220108 50948 220114
rect 50896 220050 50948 220056
rect 51000 187105 51028 288390
rect 52276 276140 52328 276146
rect 52276 276082 52328 276088
rect 52288 217394 52316 276082
rect 52380 227730 52408 288458
rect 52368 227724 52420 227730
rect 52368 227666 52420 227672
rect 52276 217388 52328 217394
rect 52276 217330 52328 217336
rect 53116 189038 53144 292606
rect 53668 218822 53696 292674
rect 54944 285796 54996 285802
rect 54944 285738 54996 285744
rect 53748 280220 53800 280226
rect 53748 280162 53800 280168
rect 53656 218816 53708 218822
rect 53656 218758 53708 218764
rect 53760 205018 53788 280162
rect 54852 258120 54904 258126
rect 54852 258062 54904 258068
rect 54864 225690 54892 258062
rect 54852 225684 54904 225690
rect 54852 225626 54904 225632
rect 53748 205012 53800 205018
rect 53748 204954 53800 204960
rect 54956 203561 54984 285738
rect 55048 249762 55076 378762
rect 56416 289876 56468 289882
rect 56416 289818 56468 289824
rect 56324 260908 56376 260914
rect 56324 260850 56376 260856
rect 55128 256760 55180 256766
rect 55128 256702 55180 256708
rect 55036 249756 55088 249762
rect 55036 249698 55088 249704
rect 54942 203552 54998 203561
rect 54942 203487 54998 203496
rect 53104 189032 53156 189038
rect 53104 188974 53156 188980
rect 50986 187096 51042 187105
rect 50986 187031 51042 187040
rect 55140 85513 55168 256702
rect 56336 235278 56364 260850
rect 56324 235272 56376 235278
rect 56324 235214 56376 235220
rect 56428 222902 56456 289818
rect 57256 267714 57284 565830
rect 58624 397520 58676 397526
rect 58624 397462 58676 397468
rect 57888 284368 57940 284374
rect 57888 284310 57940 284316
rect 57612 267776 57664 267782
rect 57612 267718 57664 267724
rect 57244 267708 57296 267714
rect 57244 267650 57296 267656
rect 56508 262268 56560 262274
rect 56508 262210 56560 262216
rect 56416 222896 56468 222902
rect 56416 222838 56468 222844
rect 56520 191282 56548 262210
rect 57624 239873 57652 267718
rect 57796 262880 57848 262886
rect 57796 262822 57848 262828
rect 57808 262342 57836 262822
rect 57796 262336 57848 262342
rect 57796 262278 57848 262284
rect 57808 258074 57836 262278
rect 57716 258046 57836 258074
rect 57610 239864 57666 239873
rect 57610 239799 57666 239808
rect 57716 218890 57744 258046
rect 57796 248464 57848 248470
rect 57796 248406 57848 248412
rect 57704 218884 57756 218890
rect 57704 218826 57756 218832
rect 57808 198082 57836 248406
rect 57900 206310 57928 284310
rect 58636 238610 58664 397462
rect 62028 352572 62080 352578
rect 62028 352514 62080 352520
rect 60648 351212 60700 351218
rect 60648 351154 60700 351160
rect 59268 287088 59320 287094
rect 59268 287030 59320 287036
rect 59176 264240 59228 264246
rect 59176 264182 59228 264188
rect 59188 263673 59216 264182
rect 59174 263664 59230 263673
rect 59174 263599 59176 263608
rect 59228 263599 59230 263608
rect 59176 263570 59228 263576
rect 59188 263539 59216 263570
rect 59084 249824 59136 249830
rect 59084 249766 59136 249772
rect 58624 238604 58676 238610
rect 58624 238546 58676 238552
rect 59096 223582 59124 249766
rect 59176 247104 59228 247110
rect 59176 247046 59228 247052
rect 59084 223576 59136 223582
rect 59084 223518 59136 223524
rect 57888 206304 57940 206310
rect 57888 206246 57940 206252
rect 57796 198076 57848 198082
rect 57796 198018 57848 198024
rect 56508 191276 56560 191282
rect 56508 191218 56560 191224
rect 59188 188329 59216 247046
rect 59280 195265 59308 287030
rect 60096 273964 60148 273970
rect 60096 273906 60148 273912
rect 60108 273290 60136 273906
rect 60096 273284 60148 273290
rect 60096 273226 60148 273232
rect 60372 273284 60424 273290
rect 60372 273226 60424 273232
rect 60384 229022 60412 273226
rect 60464 258188 60516 258194
rect 60464 258130 60516 258136
rect 60372 229016 60424 229022
rect 60372 228958 60424 228964
rect 60476 213246 60504 258130
rect 60660 258058 60688 351154
rect 61936 273352 61988 273358
rect 61936 273294 61988 273300
rect 60740 265668 60792 265674
rect 60740 265610 60792 265616
rect 60752 265062 60780 265610
rect 60740 265056 60792 265062
rect 60740 264998 60792 265004
rect 61844 265056 61896 265062
rect 61844 264998 61896 265004
rect 60648 258052 60700 258058
rect 60648 257994 60700 258000
rect 60660 257378 60688 257994
rect 60648 257372 60700 257378
rect 60648 257314 60700 257320
rect 60556 255332 60608 255338
rect 60556 255274 60608 255280
rect 60464 213240 60516 213246
rect 60464 213182 60516 213188
rect 60568 207670 60596 255274
rect 60740 253904 60792 253910
rect 60740 253846 60792 253852
rect 60752 253230 60780 253846
rect 60740 253224 60792 253230
rect 60740 253166 60792 253172
rect 60648 251864 60700 251870
rect 60648 251806 60700 251812
rect 60556 207664 60608 207670
rect 60556 207606 60608 207612
rect 59266 195256 59322 195265
rect 59266 195191 59322 195200
rect 59174 188320 59230 188329
rect 59174 188255 59230 188264
rect 60660 185774 60688 251806
rect 61856 248414 61884 264998
rect 61672 248386 61884 248414
rect 61672 233238 61700 248386
rect 61752 241664 61804 241670
rect 61752 241606 61804 241612
rect 61660 233232 61712 233238
rect 61660 233174 61712 233180
rect 61764 227254 61792 241606
rect 61842 240136 61898 240145
rect 61842 240071 61898 240080
rect 61856 238814 61884 240071
rect 61844 238808 61896 238814
rect 61844 238750 61896 238756
rect 61752 227248 61804 227254
rect 61752 227190 61804 227196
rect 61948 218657 61976 273294
rect 62040 253910 62068 352514
rect 62776 267102 62804 669938
rect 64788 361616 64840 361622
rect 64788 361558 64840 361564
rect 64602 298208 64658 298217
rect 64602 298143 64658 298152
rect 63408 277432 63460 277438
rect 63408 277374 63460 277380
rect 62764 267096 62816 267102
rect 62764 267038 62816 267044
rect 63316 267096 63368 267102
rect 63316 267038 63368 267044
rect 63224 259480 63276 259486
rect 63224 259422 63276 259428
rect 63132 253972 63184 253978
rect 63132 253914 63184 253920
rect 62028 253904 62080 253910
rect 62028 253846 62080 253852
rect 62028 247172 62080 247178
rect 62028 247114 62080 247120
rect 61934 218648 61990 218657
rect 61934 218583 61990 218592
rect 62040 189786 62068 247114
rect 63144 234598 63172 253914
rect 63236 239426 63264 259422
rect 63224 239420 63276 239426
rect 63224 239362 63276 239368
rect 63328 238066 63356 267038
rect 63316 238060 63368 238066
rect 63316 238002 63368 238008
rect 63132 234592 63184 234598
rect 63132 234534 63184 234540
rect 63420 194002 63448 277374
rect 64616 271862 64644 298143
rect 64800 282878 64828 361558
rect 66168 296812 66220 296818
rect 66168 296754 66220 296760
rect 66180 284306 66208 296754
rect 66916 293049 66944 670686
rect 79324 360256 79376 360262
rect 79324 360198 79376 360204
rect 68836 356244 68888 356250
rect 68836 356186 68888 356192
rect 67548 356176 67600 356182
rect 67548 356118 67600 356124
rect 67456 294092 67508 294098
rect 67456 294034 67508 294040
rect 66902 293040 66958 293049
rect 66902 292975 66958 292984
rect 66916 286385 66944 292975
rect 67468 289134 67496 294034
rect 67456 289128 67508 289134
rect 67456 289070 67508 289076
rect 66902 286376 66958 286385
rect 66902 286311 66958 286320
rect 66168 284300 66220 284306
rect 66168 284242 66220 284248
rect 64788 282872 64840 282878
rect 64788 282814 64840 282820
rect 67560 278905 67588 356118
rect 68560 296744 68612 296750
rect 68560 296686 68612 296692
rect 67638 290456 67694 290465
rect 67638 290391 67694 290400
rect 67652 289882 67680 290391
rect 67640 289876 67692 289882
rect 67640 289818 67692 289824
rect 67730 289776 67786 289785
rect 67730 289711 67786 289720
rect 67638 289096 67694 289105
rect 67638 289031 67694 289040
rect 67652 288454 67680 289031
rect 67744 288522 67772 289711
rect 67732 288516 67784 288522
rect 67732 288458 67784 288464
rect 67640 288448 67692 288454
rect 67640 288390 67692 288396
rect 67638 287736 67694 287745
rect 67638 287671 67694 287680
rect 67652 287094 67680 287671
rect 67640 287088 67692 287094
rect 67640 287030 67692 287036
rect 67730 287056 67786 287065
rect 67730 286991 67786 287000
rect 67744 285802 67772 286991
rect 67732 285796 67784 285802
rect 67732 285738 67784 285744
rect 67640 285728 67692 285734
rect 67638 285696 67640 285705
rect 67692 285696 67694 285705
rect 67638 285631 67694 285640
rect 68572 285025 68600 296686
rect 68744 292596 68796 292602
rect 68744 292538 68796 292544
rect 68756 291145 68784 292538
rect 68742 291136 68798 291145
rect 68742 291071 68798 291080
rect 68756 290494 68784 291071
rect 68744 290488 68796 290494
rect 68744 290430 68796 290436
rect 68848 288425 68876 356186
rect 68928 356108 68980 356114
rect 68928 356050 68980 356056
rect 68834 288416 68890 288425
rect 68834 288351 68890 288360
rect 68558 285016 68614 285025
rect 68558 284951 68614 284960
rect 67640 284368 67692 284374
rect 67638 284336 67640 284345
rect 67692 284336 67694 284345
rect 67638 284271 67694 284280
rect 67824 284300 67876 284306
rect 67824 284242 67876 284248
rect 67730 283656 67786 283665
rect 67730 283591 67786 283600
rect 67744 282946 67772 283591
rect 67836 282985 67864 284242
rect 67822 282976 67878 282985
rect 67732 282940 67784 282946
rect 67822 282911 67878 282920
rect 67732 282882 67784 282888
rect 67640 282872 67692 282878
rect 67640 282814 67692 282820
rect 67652 281625 67680 282814
rect 67638 281616 67694 281625
rect 67638 281551 67694 281560
rect 68282 280936 68338 280945
rect 68282 280871 68338 280880
rect 67638 280256 67694 280265
rect 67638 280191 67640 280200
rect 67692 280191 67694 280200
rect 67640 280162 67692 280168
rect 67638 279576 67694 279585
rect 67638 279511 67694 279520
rect 67546 278896 67602 278905
rect 67546 278831 67602 278840
rect 67652 278798 67680 279511
rect 67640 278792 67692 278798
rect 67640 278734 67692 278740
rect 68098 278216 68154 278225
rect 68098 278151 68154 278160
rect 68112 277846 68140 278151
rect 65984 277840 66036 277846
rect 65984 277782 66036 277788
rect 68100 277840 68152 277846
rect 68100 277782 68152 277788
rect 64696 274780 64748 274786
rect 64696 274722 64748 274728
rect 64604 271856 64656 271862
rect 64604 271798 64656 271804
rect 64512 253224 64564 253230
rect 64512 253166 64564 253172
rect 64524 236706 64552 253166
rect 64604 249892 64656 249898
rect 64604 249834 64656 249840
rect 64512 236700 64564 236706
rect 64512 236642 64564 236648
rect 64616 233918 64644 249834
rect 64604 233912 64656 233918
rect 64604 233854 64656 233860
rect 64708 213926 64736 274722
rect 64788 271924 64840 271930
rect 64788 271866 64840 271872
rect 64696 213920 64748 213926
rect 64696 213862 64748 213868
rect 63408 193996 63460 194002
rect 63408 193938 63460 193944
rect 62028 189780 62080 189786
rect 62028 189722 62080 189728
rect 60648 185768 60700 185774
rect 60648 185710 60700 185716
rect 64800 181529 64828 271866
rect 65892 244316 65944 244322
rect 65892 244258 65944 244264
rect 65904 206446 65932 244258
rect 65996 229770 66024 277782
rect 67638 277536 67694 277545
rect 67638 277471 67694 277480
rect 67652 277438 67680 277471
rect 67640 277432 67692 277438
rect 67640 277374 67692 277380
rect 67730 276856 67786 276865
rect 67730 276791 67786 276800
rect 67638 276176 67694 276185
rect 67744 276146 67772 276791
rect 67638 276111 67694 276120
rect 67732 276140 67784 276146
rect 67652 276078 67680 276111
rect 67732 276082 67784 276088
rect 67640 276072 67692 276078
rect 67640 276014 67692 276020
rect 67638 275496 67694 275505
rect 67638 275431 67694 275440
rect 67454 274816 67510 274825
rect 67652 274786 67680 275431
rect 67454 274751 67510 274760
rect 67640 274780 67692 274786
rect 67362 269376 67418 269385
rect 67362 269311 67418 269320
rect 66168 268252 66220 268258
rect 66168 268194 66220 268200
rect 66076 260976 66128 260982
rect 66076 260918 66128 260924
rect 65984 229764 66036 229770
rect 65984 229706 66036 229712
rect 65892 206440 65944 206446
rect 65892 206382 65944 206388
rect 66088 185638 66116 260918
rect 66076 185632 66128 185638
rect 66076 185574 66128 185580
rect 64786 181520 64842 181529
rect 64786 181455 64842 181464
rect 66180 180198 66208 268194
rect 67270 251696 67326 251705
rect 67270 251631 67326 251640
rect 66168 180192 66220 180198
rect 66168 180134 66220 180140
rect 66904 163532 66956 163538
rect 66904 163474 66956 163480
rect 66074 129296 66130 129305
rect 66074 129231 66130 129240
rect 66088 128382 66116 129231
rect 60648 128376 60700 128382
rect 60648 128318 60700 128324
rect 66076 128376 66128 128382
rect 66076 128318 66128 128324
rect 57888 125656 57940 125662
rect 57888 125598 57940 125604
rect 57900 89729 57928 125598
rect 60660 94897 60688 128318
rect 66166 126304 66222 126313
rect 66166 126239 66222 126248
rect 66180 125662 66208 126239
rect 66168 125656 66220 125662
rect 66168 125598 66220 125604
rect 66166 125216 66222 125225
rect 66166 125151 66222 125160
rect 66180 124273 66208 125151
rect 64786 124264 64842 124273
rect 64786 124199 64842 124208
rect 66166 124264 66222 124273
rect 66166 124199 66222 124208
rect 63316 122868 63368 122874
rect 63316 122810 63368 122816
rect 60646 94888 60702 94897
rect 60646 94823 60702 94832
rect 57886 89720 57942 89729
rect 63328 89690 63356 122810
rect 63408 121508 63460 121514
rect 63408 121450 63460 121456
rect 57886 89655 57942 89664
rect 63316 89684 63368 89690
rect 63316 89626 63368 89632
rect 63420 86902 63448 121450
rect 64694 102232 64750 102241
rect 64694 102167 64750 102176
rect 64708 87990 64736 102167
rect 64800 91050 64828 124199
rect 66074 123584 66130 123593
rect 66074 123519 66130 123528
rect 66088 122874 66116 123519
rect 66076 122868 66128 122874
rect 66076 122810 66128 122816
rect 66166 122632 66222 122641
rect 66166 122567 66222 122576
rect 66180 121514 66208 122567
rect 66168 121508 66220 121514
rect 66168 121450 66220 121456
rect 64788 91044 64840 91050
rect 64788 90986 64840 90992
rect 64696 87984 64748 87990
rect 64696 87926 64748 87932
rect 63408 86896 63460 86902
rect 63408 86838 63460 86844
rect 55126 85504 55182 85513
rect 55126 85439 55182 85448
rect 66916 77246 66944 163474
rect 67284 82822 67312 251631
rect 67376 227050 67404 269311
rect 67364 227044 67416 227050
rect 67364 226986 67416 226992
rect 67468 188465 67496 274751
rect 67640 274722 67692 274728
rect 67730 274136 67786 274145
rect 67730 274071 67786 274080
rect 67638 273456 67694 273465
rect 67638 273391 67694 273400
rect 67652 273358 67680 273391
rect 67640 273352 67692 273358
rect 67640 273294 67692 273300
rect 67744 273290 67772 274071
rect 67732 273284 67784 273290
rect 67732 273226 67784 273232
rect 67638 272776 67694 272785
rect 67638 272711 67694 272720
rect 67652 271930 67680 272711
rect 67640 271924 67692 271930
rect 67640 271866 67692 271872
rect 67732 271856 67784 271862
rect 67732 271798 67784 271804
rect 67638 271416 67694 271425
rect 67638 271351 67694 271360
rect 67652 270570 67680 271351
rect 67744 270745 67772 271798
rect 67730 270736 67786 270745
rect 67730 270671 67786 270680
rect 67640 270564 67692 270570
rect 67640 270506 67692 270512
rect 67638 270056 67694 270065
rect 67638 269991 67694 270000
rect 67652 269142 67680 269991
rect 67640 269136 67692 269142
rect 67640 269078 67692 269084
rect 68190 268696 68246 268705
rect 68190 268631 68246 268640
rect 68204 268258 68232 268631
rect 68192 268252 68244 268258
rect 68192 268194 68244 268200
rect 67638 268016 67694 268025
rect 67638 267951 67694 267960
rect 67652 267782 67680 267951
rect 67640 267776 67692 267782
rect 67640 267718 67692 267724
rect 67640 267096 67692 267102
rect 67640 267038 67692 267044
rect 67652 266665 67680 267038
rect 67638 266656 67694 266665
rect 67638 266591 67694 266600
rect 67730 265976 67786 265985
rect 67730 265911 67786 265920
rect 67638 265296 67694 265305
rect 67638 265231 67694 265240
rect 67652 265062 67680 265231
rect 67640 265056 67692 265062
rect 67640 264998 67692 265004
rect 67744 264994 67772 265911
rect 67732 264988 67784 264994
rect 67732 264930 67784 264936
rect 67638 264616 67694 264625
rect 67638 264551 67694 264560
rect 67652 264246 67680 264551
rect 67640 264240 67692 264246
rect 67640 264182 67692 264188
rect 67638 263936 67694 263945
rect 67638 263871 67694 263880
rect 67652 263702 67680 263871
rect 67640 263696 67692 263702
rect 67640 263638 67692 263644
rect 67730 263256 67786 263265
rect 67730 263191 67786 263200
rect 67638 262576 67694 262585
rect 67638 262511 67694 262520
rect 67652 262274 67680 262511
rect 67744 262342 67772 263191
rect 67732 262336 67784 262342
rect 67732 262278 67784 262284
rect 67640 262268 67692 262274
rect 67640 262210 67692 262216
rect 67730 261896 67786 261905
rect 67730 261831 67786 261840
rect 67744 260914 67772 261831
rect 68190 261216 68246 261225
rect 68190 261151 68246 261160
rect 68204 260982 68232 261151
rect 68192 260976 68244 260982
rect 68192 260918 68244 260924
rect 67732 260908 67784 260914
rect 67732 260850 67784 260856
rect 67640 260840 67692 260846
rect 67640 260782 67692 260788
rect 67652 260545 67680 260782
rect 67638 260536 67694 260545
rect 67638 260471 67694 260480
rect 67638 259856 67694 259865
rect 67638 259791 67694 259800
rect 67652 259486 67680 259791
rect 67640 259480 67692 259486
rect 67640 259422 67692 259428
rect 67730 259176 67786 259185
rect 67730 259111 67786 259120
rect 67638 258496 67694 258505
rect 67638 258431 67694 258440
rect 67652 258194 67680 258431
rect 67640 258188 67692 258194
rect 67640 258130 67692 258136
rect 67744 258126 67772 259111
rect 67732 258120 67784 258126
rect 67732 258062 67784 258068
rect 67640 258052 67692 258058
rect 67640 257994 67692 258000
rect 67652 257825 67680 257994
rect 67638 257816 67694 257825
rect 67638 257751 67694 257760
rect 67638 257136 67694 257145
rect 67638 257071 67694 257080
rect 67652 256766 67680 257071
rect 67640 256760 67692 256766
rect 67640 256702 67692 256708
rect 67638 255776 67694 255785
rect 67638 255711 67694 255720
rect 67652 255338 67680 255711
rect 67640 255332 67692 255338
rect 67640 255274 67692 255280
rect 67730 254416 67786 254425
rect 67730 254351 67786 254360
rect 67744 253978 67772 254351
rect 67732 253972 67784 253978
rect 67732 253914 67784 253920
rect 67640 253904 67692 253910
rect 67640 253846 67692 253852
rect 67652 253745 67680 253846
rect 67638 253736 67694 253745
rect 67638 253671 67694 253680
rect 68296 253230 68324 280871
rect 68374 272096 68430 272105
rect 68374 272031 68430 272040
rect 68284 253224 68336 253230
rect 68284 253166 68336 253172
rect 68388 251870 68416 272031
rect 68940 267714 68968 356050
rect 75920 355088 75972 355094
rect 75920 355030 75972 355036
rect 72424 354748 72476 354754
rect 72424 354690 72476 354696
rect 72436 306374 72464 354690
rect 72252 306346 72464 306374
rect 72252 304978 72280 306346
rect 72240 304972 72292 304978
rect 72240 304914 72292 304920
rect 70952 300144 71004 300150
rect 70952 300086 71004 300092
rect 70032 294636 70084 294642
rect 70032 294578 70084 294584
rect 70044 291924 70072 294578
rect 70674 292632 70730 292641
rect 70674 292567 70730 292576
rect 70688 291924 70716 292567
rect 70964 291938 70992 300086
rect 71964 292732 72016 292738
rect 71964 292674 72016 292680
rect 71688 292528 71740 292534
rect 71688 292470 71740 292476
rect 71700 292369 71728 292470
rect 71686 292360 71742 292369
rect 71686 292295 71742 292304
rect 70964 291910 71346 291938
rect 71976 291924 72004 292674
rect 72252 291938 72280 304914
rect 74540 303680 74592 303686
rect 74540 303622 74592 303628
rect 73252 298172 73304 298178
rect 73252 298114 73304 298120
rect 72252 291910 72634 291938
rect 73264 291924 73292 298114
rect 73894 294536 73950 294545
rect 73894 294471 73950 294480
rect 73908 291924 73936 294471
rect 74552 291924 74580 303622
rect 75368 300892 75420 300898
rect 75368 300834 75420 300840
rect 75184 298240 75236 298246
rect 75184 298182 75236 298188
rect 75196 291924 75224 298182
rect 75380 291938 75408 300834
rect 75932 293962 75960 355030
rect 76104 301096 76156 301102
rect 76104 301038 76156 301044
rect 75920 293956 75972 293962
rect 75920 293898 75972 293904
rect 76116 291938 76144 301038
rect 78404 295656 78456 295662
rect 78404 295598 78456 295604
rect 76748 293956 76800 293962
rect 76748 293898 76800 293904
rect 76760 291938 76788 293898
rect 77758 292768 77814 292777
rect 77758 292703 77814 292712
rect 75380 291910 75854 291938
rect 76116 291910 76498 291938
rect 76760 291910 77142 291938
rect 77772 291924 77800 292703
rect 78416 291924 78444 295598
rect 79336 294098 79364 360198
rect 80060 357468 80112 357474
rect 80060 357410 80112 357416
rect 79692 294704 79744 294710
rect 79692 294646 79744 294652
rect 79324 294092 79376 294098
rect 79324 294034 79376 294040
rect 79336 291938 79364 294034
rect 79074 291910 79364 291938
rect 79704 291924 79732 294646
rect 80072 291938 80100 357410
rect 84292 354068 84344 354074
rect 84292 354010 84344 354016
rect 81440 305176 81492 305182
rect 81440 305118 81492 305124
rect 80980 294432 81032 294438
rect 80980 294374 81032 294380
rect 80072 291910 80362 291938
rect 80992 291924 81020 294374
rect 81452 291938 81480 305118
rect 83556 296948 83608 296954
rect 83556 296890 83608 296896
rect 82268 295588 82320 295594
rect 82268 295530 82320 295536
rect 81452 291910 81650 291938
rect 82280 291924 82308 295530
rect 82912 294228 82964 294234
rect 82912 294170 82964 294176
rect 82924 291924 82952 294170
rect 83568 291924 83596 296890
rect 84200 295724 84252 295730
rect 84200 295666 84252 295672
rect 84212 291924 84240 295666
rect 84304 293962 84332 354010
rect 84384 307080 84436 307086
rect 84384 307022 84436 307028
rect 84396 299606 84424 307022
rect 88352 303618 88380 702406
rect 105464 700330 105492 703520
rect 94504 700324 94556 700330
rect 94504 700266 94556 700272
rect 105452 700324 105504 700330
rect 105452 700266 105504 700272
rect 90364 605872 90416 605878
rect 90364 605814 90416 605820
rect 88432 305108 88484 305114
rect 88432 305050 88484 305056
rect 88340 303612 88392 303618
rect 88340 303554 88392 303560
rect 85580 301028 85632 301034
rect 85580 300970 85632 300976
rect 84384 299600 84436 299606
rect 84384 299542 84436 299548
rect 84292 293956 84344 293962
rect 84292 293898 84344 293904
rect 84396 291938 84424 299542
rect 84476 295724 84528 295730
rect 84476 295666 84528 295672
rect 84488 295526 84516 295666
rect 84476 295520 84528 295526
rect 84476 295462 84528 295468
rect 85592 293962 85620 300970
rect 85672 300960 85724 300966
rect 85672 300902 85724 300908
rect 85212 293956 85264 293962
rect 85212 293898 85264 293904
rect 85580 293956 85632 293962
rect 85580 293898 85632 293904
rect 85224 291938 85252 293898
rect 85684 291938 85712 300902
rect 88340 299804 88392 299810
rect 88340 299746 88392 299752
rect 87420 297016 87472 297022
rect 87420 296958 87472 296964
rect 86500 293956 86552 293962
rect 86500 293898 86552 293904
rect 86512 291938 86540 293898
rect 84396 291910 84870 291938
rect 85224 291910 85514 291938
rect 85684 291910 86158 291938
rect 86512 291910 86802 291938
rect 87432 291924 87460 296958
rect 88352 293962 88380 299746
rect 88340 293956 88392 293962
rect 88340 293898 88392 293904
rect 88064 292800 88116 292806
rect 88064 292742 88116 292748
rect 88076 291924 88104 292742
rect 88444 291938 88472 305050
rect 90376 304774 90404 605814
rect 91100 307080 91152 307086
rect 91100 307022 91152 307028
rect 90364 304768 90416 304774
rect 90364 304710 90416 304716
rect 89720 302456 89772 302462
rect 89720 302398 89772 302404
rect 88984 295588 89036 295594
rect 88984 295530 89036 295536
rect 88996 295390 89024 295530
rect 88984 295384 89036 295390
rect 88984 295326 89036 295332
rect 89076 293956 89128 293962
rect 89076 293898 89128 293904
rect 89088 291938 89116 293898
rect 89732 291938 89760 302398
rect 90640 298376 90692 298382
rect 90640 298318 90692 298324
rect 88444 291910 88734 291938
rect 89088 291910 89378 291938
rect 89732 291910 90022 291938
rect 90652 291924 90680 298318
rect 91112 291938 91140 307022
rect 94516 304978 94544 700266
rect 137848 699802 137876 703520
rect 154132 702434 154160 703520
rect 153212 702406 154160 702434
rect 149704 700392 149756 700398
rect 149704 700334 149756 700340
rect 137848 699774 138060 699802
rect 120724 501016 120776 501022
rect 120724 500958 120776 500964
rect 98644 462392 98696 462398
rect 98644 462334 98696 462340
rect 98656 371890 98684 462334
rect 98644 371884 98696 371890
rect 98644 371826 98696 371832
rect 111064 371272 111116 371278
rect 111064 371214 111116 371220
rect 109040 358964 109092 358970
rect 109040 358906 109092 358912
rect 101404 358896 101456 358902
rect 101404 358838 101456 358844
rect 96620 355156 96672 355162
rect 96620 355098 96672 355104
rect 96632 306374 96660 355098
rect 98644 324964 98696 324970
rect 98644 324906 98696 324912
rect 96632 306346 96752 306374
rect 94504 304972 94556 304978
rect 94504 304914 94556 304920
rect 94596 304768 94648 304774
rect 94596 304710 94648 304716
rect 92848 302320 92900 302326
rect 92848 302262 92900 302268
rect 92572 292936 92624 292942
rect 92572 292878 92624 292884
rect 91928 292732 91980 292738
rect 91928 292674 91980 292680
rect 91112 291910 91310 291938
rect 91940 291924 91968 292674
rect 92584 292670 92612 292878
rect 92572 292664 92624 292670
rect 92572 292606 92624 292612
rect 92584 291924 92612 292606
rect 92860 291938 92888 302262
rect 94608 296993 94636 304710
rect 94594 296984 94650 296993
rect 94594 296919 94650 296928
rect 93860 294160 93912 294166
rect 93860 294102 93912 294108
rect 92860 291910 93242 291938
rect 93872 291924 93900 294102
rect 94608 291938 94636 296919
rect 95146 296032 95202 296041
rect 95146 295967 95202 295976
rect 94530 291910 94636 291938
rect 95160 291924 95188 295967
rect 95790 294128 95846 294137
rect 95790 294063 95846 294072
rect 95804 291924 95832 294063
rect 96436 294024 96488 294030
rect 96436 293966 96488 293972
rect 96448 291924 96476 293966
rect 96724 291938 96752 306346
rect 98656 300830 98684 324906
rect 99380 311908 99432 311914
rect 99380 311850 99432 311856
rect 99392 307086 99420 311850
rect 99380 307080 99432 307086
rect 99380 307022 99432 307028
rect 99380 302388 99432 302394
rect 99380 302330 99432 302336
rect 98736 302252 98788 302258
rect 98736 302194 98788 302200
rect 98000 300824 98052 300830
rect 98000 300766 98052 300772
rect 98644 300824 98696 300830
rect 98644 300766 98696 300772
rect 98012 299674 98040 300766
rect 98552 299736 98604 299742
rect 98552 299678 98604 299684
rect 98000 299668 98052 299674
rect 98000 299610 98052 299616
rect 97722 298344 97778 298353
rect 97722 298279 97778 298288
rect 96724 291910 97106 291938
rect 97736 291924 97764 298279
rect 98012 291938 98040 299610
rect 98564 291938 98592 299678
rect 98748 294545 98776 302194
rect 98734 294536 98790 294545
rect 98734 294471 98790 294480
rect 99392 291938 99420 302330
rect 101416 295458 101444 358838
rect 107660 354952 107712 354958
rect 107660 354894 107712 354900
rect 106280 334008 106332 334014
rect 106280 333950 106332 333956
rect 104164 333260 104216 333266
rect 104164 333202 104216 333208
rect 104176 303618 104204 333202
rect 106292 306374 106320 333950
rect 107672 306374 107700 354894
rect 109052 306374 109080 358906
rect 106292 306346 107056 306374
rect 107672 306346 108344 306374
rect 109052 306346 109632 306374
rect 103796 303612 103848 303618
rect 103796 303554 103848 303560
rect 104164 303612 104216 303618
rect 104164 303554 104216 303560
rect 102140 301164 102192 301170
rect 102140 301106 102192 301112
rect 101404 295452 101456 295458
rect 101404 295394 101456 295400
rect 101416 291938 101444 295394
rect 102152 291938 102180 301106
rect 102876 298444 102928 298450
rect 102876 298386 102928 298392
rect 98012 291910 98394 291938
rect 98564 291910 99038 291938
rect 99392 291910 99682 291938
rect 100970 291922 101352 291938
rect 100970 291916 101364 291922
rect 100970 291910 101312 291916
rect 101416 291910 101614 291938
rect 102152 291910 102258 291938
rect 102888 291924 102916 298386
rect 103518 294264 103574 294273
rect 103518 294199 103574 294208
rect 103532 291924 103560 294199
rect 103808 294030 103836 303554
rect 104164 301232 104216 301238
rect 104164 301174 104216 301180
rect 104176 294710 104204 301174
rect 104348 296880 104400 296886
rect 104348 296822 104400 296828
rect 104164 294704 104216 294710
rect 104164 294646 104216 294652
rect 103796 294024 103848 294030
rect 103796 293966 103848 293972
rect 104360 291938 104388 296822
rect 105452 295452 105504 295458
rect 105452 295394 105504 295400
rect 104532 294024 104584 294030
rect 104532 293966 104584 293972
rect 104190 291910 104388 291938
rect 104544 291938 104572 293966
rect 104544 291910 104834 291938
rect 105464 291924 105492 295394
rect 106096 294364 106148 294370
rect 106096 294306 106148 294312
rect 106108 291924 106136 294306
rect 106738 293992 106794 294001
rect 106738 293927 106794 293936
rect 106752 291924 106780 293927
rect 107028 291938 107056 306346
rect 108026 292904 108082 292913
rect 108026 292839 108082 292848
rect 107028 291910 107410 291938
rect 108040 291924 108068 292839
rect 108316 291938 108344 306346
rect 109316 292664 109368 292670
rect 109316 292606 109368 292612
rect 108316 291910 108698 291938
rect 109328 291924 109356 292606
rect 109604 291938 109632 306346
rect 111076 298790 111104 371214
rect 114560 367260 114612 367266
rect 114560 367202 114612 367208
rect 111156 361752 111208 361758
rect 111156 361694 111208 361700
rect 111064 298784 111116 298790
rect 111064 298726 111116 298732
rect 110604 292868 110656 292874
rect 110604 292810 110656 292816
rect 109604 291910 109986 291938
rect 110616 291924 110644 292810
rect 111168 292534 111196 361694
rect 113180 360392 113232 360398
rect 113180 360334 113232 360340
rect 111892 295724 111944 295730
rect 111892 295666 111944 295672
rect 111246 295352 111302 295361
rect 111246 295287 111302 295296
rect 111156 292528 111208 292534
rect 111156 292470 111208 292476
rect 111260 291924 111288 295287
rect 111904 291924 111932 295666
rect 112562 291922 112852 291938
rect 113192 291924 113220 360334
rect 114468 294296 114520 294302
rect 114468 294238 114520 294244
rect 114190 291952 114246 291961
rect 112562 291916 112864 291922
rect 112562 291910 112812 291916
rect 101312 291858 101364 291864
rect 113850 291910 114190 291938
rect 114480 291924 114508 294238
rect 114572 294030 114600 367202
rect 120736 364410 120764 500958
rect 138032 378826 138060 699774
rect 138020 378820 138072 378826
rect 138020 378762 138072 378768
rect 125600 371884 125652 371890
rect 125600 371826 125652 371832
rect 126612 371884 126664 371890
rect 126612 371826 126664 371832
rect 120724 364404 120776 364410
rect 120724 364346 120776 364352
rect 117964 351280 118016 351286
rect 117964 351222 118016 351228
rect 116584 318844 116636 318850
rect 116584 318786 116636 318792
rect 114744 306400 114796 306406
rect 114744 306342 114796 306348
rect 114756 304978 114784 306342
rect 114744 304972 114796 304978
rect 114744 304914 114796 304920
rect 114560 294024 114612 294030
rect 114560 293966 114612 293972
rect 114756 291938 114784 304914
rect 116596 298314 116624 318786
rect 117976 299538 118004 351222
rect 118700 311160 118752 311166
rect 118700 311102 118752 311108
rect 118712 310486 118740 311102
rect 118700 310480 118752 310486
rect 118700 310422 118752 310428
rect 118712 306374 118740 310422
rect 118712 306346 119476 306374
rect 117964 299532 118016 299538
rect 117964 299474 118016 299480
rect 116584 298308 116636 298314
rect 116584 298250 116636 298256
rect 115388 294024 115440 294030
rect 115388 293966 115440 293972
rect 115400 291938 115428 293966
rect 116596 291938 116624 298250
rect 117976 296714 118004 299474
rect 117884 296686 118004 296714
rect 117228 295656 117280 295662
rect 117228 295598 117280 295604
rect 117240 294642 117268 295598
rect 117228 294636 117280 294642
rect 117228 294578 117280 294584
rect 116860 294228 116912 294234
rect 116860 294170 116912 294176
rect 114756 291910 115138 291938
rect 115400 291910 115782 291938
rect 116426 291910 116624 291938
rect 116872 291922 116900 294170
rect 117226 294128 117282 294137
rect 117226 294063 117282 294072
rect 117686 294128 117742 294137
rect 117686 294063 117742 294072
rect 117240 294030 117268 294063
rect 117228 294024 117280 294030
rect 117228 293966 117280 293972
rect 117320 291984 117372 291990
rect 117070 291932 117320 291938
rect 117070 291926 117372 291932
rect 116860 291916 116912 291922
rect 114190 291887 114246 291896
rect 112812 291858 112864 291864
rect 117070 291910 117360 291926
rect 117700 291924 117728 294063
rect 117884 291938 117912 296686
rect 119448 291938 119476 306346
rect 119712 291984 119764 291990
rect 117884 291910 118358 291938
rect 119002 291922 119384 291938
rect 119002 291916 119396 291922
rect 119002 291910 119344 291916
rect 116860 291858 116912 291864
rect 119448 291910 119646 291938
rect 119712 291926 119764 291932
rect 119344 291858 119396 291864
rect 68928 267708 68980 267714
rect 68928 267650 68980 267656
rect 68940 267345 68968 267650
rect 68926 267336 68982 267345
rect 68926 267271 68982 267280
rect 69202 256456 69258 256465
rect 69202 256391 69258 256400
rect 69018 253056 69074 253065
rect 69018 252991 69074 253000
rect 68926 252376 68982 252385
rect 68926 252311 68982 252320
rect 68376 251864 68428 251870
rect 68376 251806 68428 251812
rect 67730 251016 67786 251025
rect 67730 250951 67786 250960
rect 67638 250336 67694 250345
rect 67638 250271 67694 250280
rect 67652 249898 67680 250271
rect 67640 249892 67692 249898
rect 67640 249834 67692 249840
rect 67744 249830 67772 250951
rect 67732 249824 67784 249830
rect 67732 249766 67784 249772
rect 67640 249756 67692 249762
rect 67640 249698 67692 249704
rect 67652 249665 67680 249698
rect 67638 249656 67694 249665
rect 67638 249591 67694 249600
rect 67638 248976 67694 248985
rect 67638 248911 67694 248920
rect 67652 248470 67680 248911
rect 67640 248464 67692 248470
rect 67640 248406 67692 248412
rect 67730 248296 67786 248305
rect 67730 248231 67786 248240
rect 67638 247616 67694 247625
rect 67638 247551 67694 247560
rect 67652 247178 67680 247551
rect 67640 247172 67692 247178
rect 67640 247114 67692 247120
rect 67744 247110 67772 248231
rect 67732 247104 67784 247110
rect 67732 247046 67784 247052
rect 68100 245608 68152 245614
rect 68098 245576 68100 245585
rect 68152 245576 68154 245585
rect 68098 245511 68154 245520
rect 68006 244896 68062 244905
rect 68006 244831 68062 244840
rect 68020 244322 68048 244831
rect 68008 244316 68060 244322
rect 68008 244258 68060 244264
rect 67546 244216 67602 244225
rect 67546 244151 67602 244160
rect 67560 235958 67588 244151
rect 67638 242176 67694 242185
rect 67638 242111 67694 242120
rect 67652 241670 67680 242111
rect 67640 241664 67692 241670
rect 67640 241606 67692 241612
rect 67548 235952 67600 235958
rect 67548 235894 67600 235900
rect 67454 188456 67510 188465
rect 67454 188391 67510 188400
rect 68940 180130 68968 252311
rect 69032 203590 69060 252991
rect 69112 233980 69164 233986
rect 69112 233922 69164 233928
rect 69020 203584 69072 203590
rect 69020 203526 69072 203532
rect 69124 196654 69152 233922
rect 69216 220182 69244 256391
rect 69294 245576 69350 245585
rect 69294 245511 69350 245520
rect 69308 234530 69336 245511
rect 69768 240094 70058 240122
rect 69296 234524 69348 234530
rect 69296 234466 69348 234472
rect 69768 233986 69796 240094
rect 69756 233980 69808 233986
rect 69756 233922 69808 233928
rect 70688 232626 70716 240108
rect 70676 232620 70728 232626
rect 70676 232562 70728 232568
rect 69204 220176 69256 220182
rect 69204 220118 69256 220124
rect 71332 219434 71360 240108
rect 71976 219434 72004 240108
rect 72620 235754 72648 240108
rect 73264 238754 73292 240108
rect 73172 238726 73292 238754
rect 72608 235748 72660 235754
rect 72608 235690 72660 235696
rect 70412 219406 71360 219434
rect 71792 219406 72004 219434
rect 70412 216034 70440 219406
rect 70400 216028 70452 216034
rect 70400 215970 70452 215976
rect 69112 196648 69164 196654
rect 69112 196590 69164 196596
rect 71792 192506 71820 219406
rect 71780 192500 71832 192506
rect 71780 192442 71832 192448
rect 73172 186969 73200 238726
rect 73908 219434 73936 240108
rect 74552 238754 74580 240108
rect 74552 238726 74672 238754
rect 74540 233980 74592 233986
rect 74540 233922 74592 233928
rect 73264 219406 73936 219434
rect 73264 203726 73292 219406
rect 73252 203720 73304 203726
rect 73252 203662 73304 203668
rect 73158 186960 73214 186969
rect 73158 186895 73214 186904
rect 74552 181393 74580 233922
rect 74644 193866 74672 238726
rect 75196 233986 75224 240108
rect 75184 233980 75236 233986
rect 75184 233922 75236 233928
rect 75840 230489 75868 240108
rect 76484 233102 76512 240108
rect 76564 239420 76616 239426
rect 76564 239362 76616 239368
rect 76472 233096 76524 233102
rect 76472 233038 76524 233044
rect 75826 230480 75882 230489
rect 75826 230415 75882 230424
rect 76576 214606 76604 239362
rect 77128 238134 77156 240108
rect 77772 238754 77800 240108
rect 77312 238726 77800 238754
rect 77116 238128 77168 238134
rect 77116 238070 77168 238076
rect 76564 214600 76616 214606
rect 76564 214542 76616 214548
rect 74632 193860 74684 193866
rect 74632 193802 74684 193808
rect 77312 184210 77340 238726
rect 78416 219434 78444 240108
rect 79060 237454 79088 240108
rect 79048 237448 79100 237454
rect 79048 237390 79100 237396
rect 79704 219434 79732 240108
rect 80060 233980 80112 233986
rect 80060 233922 80112 233928
rect 77404 219406 78444 219434
rect 78692 219406 79732 219434
rect 77404 217462 77432 219406
rect 77392 217456 77444 217462
rect 77392 217398 77444 217404
rect 78692 210458 78720 219406
rect 78680 210452 78732 210458
rect 78680 210394 78732 210400
rect 80072 196790 80100 233922
rect 80348 219434 80376 240108
rect 80992 233986 81020 240108
rect 81636 238678 81664 240108
rect 81624 238672 81676 238678
rect 81624 238614 81676 238620
rect 82280 238610 82308 240108
rect 82924 238610 82952 240108
rect 82268 238604 82320 238610
rect 82268 238546 82320 238552
rect 82912 238604 82964 238610
rect 82912 238546 82964 238552
rect 80980 233980 81032 233986
rect 80980 233922 81032 233928
rect 82280 231742 82308 238546
rect 82268 231736 82320 231742
rect 82268 231678 82320 231684
rect 83568 229090 83596 240108
rect 84212 238754 84240 240108
rect 84212 238726 84332 238754
rect 84200 233980 84252 233986
rect 84200 233922 84252 233928
rect 83556 229084 83608 229090
rect 83556 229026 83608 229032
rect 83568 228410 83596 229026
rect 83556 228404 83608 228410
rect 83556 228346 83608 228352
rect 80164 219406 80376 219434
rect 80164 209438 80192 219406
rect 80152 209432 80204 209438
rect 80152 209374 80204 209380
rect 80060 196784 80112 196790
rect 80060 196726 80112 196732
rect 84212 184278 84240 233922
rect 84304 191146 84332 238726
rect 84856 233986 84884 240108
rect 84844 233980 84896 233986
rect 84844 233922 84896 233928
rect 85500 219434 85528 240108
rect 86144 233170 86172 240108
rect 86788 238746 86816 240108
rect 86776 238740 86828 238746
rect 86776 238682 86828 238688
rect 86788 238542 86816 238682
rect 86776 238536 86828 238542
rect 86776 238478 86828 238484
rect 86224 237448 86276 237454
rect 86224 237390 86276 237396
rect 86132 233164 86184 233170
rect 86132 233106 86184 233112
rect 84396 219406 85528 219434
rect 84396 207738 84424 219406
rect 86236 209302 86264 237390
rect 86960 233912 87012 233918
rect 86960 233854 87012 233860
rect 86224 209296 86276 209302
rect 86224 209238 86276 209244
rect 86972 207806 87000 233854
rect 87432 221542 87460 240108
rect 88076 233918 88104 240108
rect 88064 233912 88116 233918
rect 88064 233854 88116 233860
rect 88720 231130 88748 240108
rect 89364 238406 89392 240108
rect 90008 238754 90036 240108
rect 89732 238726 90036 238754
rect 89352 238400 89404 238406
rect 89352 238342 89404 238348
rect 88984 232620 89036 232626
rect 88984 232562 89036 232568
rect 88708 231124 88760 231130
rect 88708 231066 88760 231072
rect 87420 221536 87472 221542
rect 87420 221478 87472 221484
rect 88996 211818 89024 232562
rect 88984 211812 89036 211818
rect 88984 211754 89036 211760
rect 86960 207800 87012 207806
rect 86960 207742 87012 207748
rect 84384 207732 84436 207738
rect 84384 207674 84436 207680
rect 89732 192710 89760 238726
rect 90652 219434 90680 240108
rect 91296 235686 91324 240108
rect 91284 235680 91336 235686
rect 91284 235622 91336 235628
rect 91940 231606 91968 240108
rect 92584 238754 92612 240108
rect 92492 238726 92612 238754
rect 91928 231600 91980 231606
rect 91928 231542 91980 231548
rect 89824 219406 90680 219434
rect 89824 206514 89852 219406
rect 92492 211886 92520 238726
rect 93228 219434 93256 240108
rect 92584 219406 93256 219434
rect 92584 215966 92612 219406
rect 92572 215960 92624 215966
rect 92572 215902 92624 215908
rect 92480 211880 92532 211886
rect 92480 211822 92532 211828
rect 89812 206508 89864 206514
rect 89812 206450 89864 206456
rect 89720 192704 89772 192710
rect 89720 192646 89772 192652
rect 84292 191140 84344 191146
rect 84292 191082 84344 191088
rect 84200 184272 84252 184278
rect 84200 184214 84252 184220
rect 77300 184204 77352 184210
rect 77300 184146 77352 184152
rect 93872 182986 93900 240108
rect 94516 219434 94544 240108
rect 95160 233986 95188 240108
rect 95804 234462 95832 240108
rect 95792 234456 95844 234462
rect 95792 234398 95844 234404
rect 95148 233980 95200 233986
rect 95148 233922 95200 233928
rect 96448 233918 96476 240108
rect 97092 238754 97120 240108
rect 96632 238726 97120 238754
rect 95240 233912 95292 233918
rect 95240 233854 95292 233860
rect 96436 233912 96488 233918
rect 96436 233854 96488 233860
rect 93964 219406 94544 219434
rect 93964 196722 93992 219406
rect 93952 196716 94004 196722
rect 93952 196658 94004 196664
rect 95252 186998 95280 233854
rect 95884 233844 95936 233850
rect 95884 233786 95936 233792
rect 95896 210662 95924 233786
rect 95884 210656 95936 210662
rect 95884 210598 95936 210604
rect 96632 201006 96660 238726
rect 97736 219434 97764 240108
rect 98380 238241 98408 240108
rect 98366 238232 98422 238241
rect 98366 238167 98422 238176
rect 99024 237250 99052 240108
rect 99668 238754 99696 240108
rect 99392 238726 99696 238754
rect 99012 237244 99064 237250
rect 99012 237186 99064 237192
rect 98644 236700 98696 236706
rect 98644 236642 98696 236648
rect 96724 219406 97764 219434
rect 96724 214674 96752 219406
rect 96712 214668 96764 214674
rect 96712 214610 96764 214616
rect 96620 201000 96672 201006
rect 96620 200942 96672 200948
rect 95240 186992 95292 186998
rect 95240 186934 95292 186940
rect 93860 182980 93912 182986
rect 93860 182922 93912 182928
rect 74538 181384 74594 181393
rect 74538 181319 74594 181328
rect 68928 180124 68980 180130
rect 68928 180066 68980 180072
rect 98656 178673 98684 236642
rect 99392 198014 99420 238726
rect 100312 225622 100340 240108
rect 100760 233912 100812 233918
rect 100760 233854 100812 233860
rect 100300 225616 100352 225622
rect 100300 225558 100352 225564
rect 100772 199646 100800 233854
rect 100956 219434 100984 240108
rect 101600 233918 101628 240108
rect 102244 238754 102272 240108
rect 102152 238726 102272 238754
rect 101588 233912 101640 233918
rect 101588 233854 101640 233860
rect 100864 219406 100984 219434
rect 100864 214742 100892 219406
rect 100852 214736 100904 214742
rect 100852 214678 100904 214684
rect 100760 199640 100812 199646
rect 100760 199582 100812 199588
rect 99380 198008 99432 198014
rect 99380 197950 99432 197956
rect 102048 190528 102100 190534
rect 102048 190470 102100 190476
rect 100668 187740 100720 187746
rect 100668 187682 100720 187688
rect 98642 178664 98698 178673
rect 98642 178599 98698 178608
rect 100680 177585 100708 187682
rect 102060 177721 102088 190470
rect 102152 185706 102180 238726
rect 102888 220250 102916 240108
rect 103532 237386 103560 240108
rect 104176 238754 104204 240108
rect 103624 238726 104204 238754
rect 103520 237380 103572 237386
rect 103520 237322 103572 237328
rect 102876 220244 102928 220250
rect 102876 220186 102928 220192
rect 103624 210526 103652 238726
rect 104716 237380 104768 237386
rect 104716 237322 104768 237328
rect 104728 231674 104756 237322
rect 104716 231668 104768 231674
rect 104716 231610 104768 231616
rect 104820 219434 104848 240108
rect 105464 238754 105492 240108
rect 103716 219406 104848 219434
rect 104912 238726 105492 238754
rect 103612 210520 103664 210526
rect 103612 210462 103664 210468
rect 103716 200802 103744 219406
rect 103704 200796 103756 200802
rect 103704 200738 103756 200744
rect 103428 189100 103480 189106
rect 103428 189042 103480 189048
rect 102140 185700 102192 185706
rect 102140 185642 102192 185648
rect 102046 177712 102102 177721
rect 102046 177647 102102 177656
rect 103440 177585 103468 189042
rect 104912 187134 104940 238726
rect 106108 219434 106136 240108
rect 106752 238377 106780 240108
rect 106738 238368 106794 238377
rect 106738 238303 106794 238312
rect 106924 238128 106976 238134
rect 106924 238070 106976 238076
rect 105004 219406 106136 219434
rect 105004 216102 105032 219406
rect 104992 216096 105044 216102
rect 104992 216038 105044 216044
rect 104900 187128 104952 187134
rect 104900 187070 104952 187076
rect 106936 182850 106964 238070
rect 107396 230450 107424 240108
rect 107660 233912 107712 233918
rect 107660 233854 107712 233860
rect 107384 230444 107436 230450
rect 107384 230386 107436 230392
rect 107672 205154 107700 233854
rect 108040 219434 108068 240108
rect 108684 233918 108712 240108
rect 109972 238754 110000 240108
rect 110616 238882 110644 240108
rect 111064 239420 111116 239426
rect 111064 239362 111116 239368
rect 110420 238876 110472 238882
rect 110420 238818 110472 238824
rect 110604 238876 110656 238882
rect 110604 238818 110656 238824
rect 109696 238726 110000 238754
rect 109696 237318 109724 238726
rect 109684 237312 109736 237318
rect 109684 237254 109736 237260
rect 108672 233912 108724 233918
rect 108672 233854 108724 233860
rect 107764 219406 108068 219434
rect 107764 209098 107792 219406
rect 107752 209092 107804 209098
rect 107752 209034 107804 209040
rect 107660 205148 107712 205154
rect 107660 205090 107712 205096
rect 109696 189854 109724 237254
rect 109684 189848 109736 189854
rect 109684 189790 109736 189796
rect 106924 182844 106976 182850
rect 106924 182786 106976 182792
rect 110236 179512 110288 179518
rect 110432 179489 110460 238818
rect 111076 238610 111104 239362
rect 111064 238604 111116 238610
rect 111064 238546 111116 238552
rect 111260 219434 111288 240108
rect 111904 219434 111932 240108
rect 112548 235890 112576 240108
rect 113192 237386 113220 240108
rect 113180 237380 113232 237386
rect 113180 237322 113232 237328
rect 112536 235884 112588 235890
rect 112536 235826 112588 235832
rect 113836 235618 113864 240108
rect 114480 238746 114508 240108
rect 114468 238740 114520 238746
rect 114468 238682 114520 238688
rect 115124 238513 115152 240108
rect 115110 238504 115166 238513
rect 115110 238439 115166 238448
rect 113824 235612 113876 235618
rect 113824 235554 113876 235560
rect 115768 233918 115796 240108
rect 114560 233912 114612 233918
rect 114560 233854 114612 233860
rect 115756 233912 115808 233918
rect 115756 233854 115808 233860
rect 110524 219406 111288 219434
rect 111812 219406 111932 219434
rect 110524 202230 110552 219406
rect 111812 211954 111840 219406
rect 114572 217530 114600 233854
rect 116412 219434 116440 240108
rect 117056 239737 117084 240108
rect 117042 239728 117098 239737
rect 117042 239663 117098 239672
rect 117700 238610 117728 240108
rect 117688 238604 117740 238610
rect 117688 238546 117740 238552
rect 118344 238474 118372 240108
rect 118988 238649 119016 240108
rect 118974 238640 119030 238649
rect 118974 238575 119030 238584
rect 118332 238468 118384 238474
rect 118332 238410 118384 238416
rect 117228 238060 117280 238066
rect 117228 238002 117280 238008
rect 117240 237153 117268 238002
rect 117226 237144 117282 237153
rect 117226 237079 117282 237088
rect 116584 235272 116636 235278
rect 116584 235214 116636 235220
rect 115952 219406 116440 219434
rect 114560 217524 114612 217530
rect 114560 217466 114612 217472
rect 111800 211948 111852 211954
rect 111800 211890 111852 211896
rect 110512 202224 110564 202230
rect 110512 202166 110564 202172
rect 115952 193934 115980 219406
rect 116596 199510 116624 235214
rect 117964 222896 118016 222902
rect 117964 222838 118016 222844
rect 116584 199504 116636 199510
rect 116584 199446 116636 199452
rect 115940 193928 115992 193934
rect 115940 193870 115992 193876
rect 117976 189922 118004 222838
rect 119632 219434 119660 240108
rect 119724 235822 119752 291926
rect 119988 291916 120040 291922
rect 119988 291858 120040 291864
rect 120000 291378 120028 291858
rect 119988 291372 120040 291378
rect 119988 291314 120040 291320
rect 120736 268705 120764 364346
rect 124956 347812 125008 347818
rect 124956 347754 125008 347760
rect 122104 311160 122156 311166
rect 122104 311102 122156 311108
rect 120906 294264 120962 294273
rect 120906 294199 120962 294208
rect 120814 292768 120870 292777
rect 120814 292703 120870 292712
rect 120828 283626 120856 292703
rect 120816 283620 120868 283626
rect 120816 283562 120868 283568
rect 120814 282296 120870 282305
rect 120814 282231 120870 282240
rect 120722 268696 120778 268705
rect 120722 268631 120778 268640
rect 120724 251048 120776 251054
rect 120170 251016 120226 251025
rect 120170 250951 120226 250960
rect 120722 251016 120724 251025
rect 120776 251016 120778 251025
rect 120722 250951 120778 250960
rect 120078 241496 120134 241505
rect 120078 241431 120134 241440
rect 119712 235816 119764 235822
rect 119712 235758 119764 235764
rect 120092 232558 120120 241431
rect 120080 232552 120132 232558
rect 120080 232494 120132 232500
rect 120184 221474 120212 250951
rect 120724 233980 120776 233986
rect 120724 233922 120776 233928
rect 120172 221468 120224 221474
rect 120172 221410 120224 221416
rect 118712 219406 119660 219434
rect 118712 206378 118740 219406
rect 118700 206372 118752 206378
rect 118700 206314 118752 206320
rect 120736 199442 120764 233922
rect 120724 199436 120776 199442
rect 120724 199378 120776 199384
rect 120828 192778 120856 282231
rect 120920 242282 120948 294199
rect 121000 292936 121052 292942
rect 121000 292878 121052 292884
rect 121012 282198 121040 292878
rect 121460 292528 121512 292534
rect 121460 292470 121512 292476
rect 121472 291825 121500 292470
rect 121458 291816 121514 291825
rect 121458 291751 121514 291760
rect 121458 291136 121514 291145
rect 121458 291071 121514 291080
rect 121472 289950 121500 291071
rect 121550 290456 121606 290465
rect 121550 290391 121606 290400
rect 121460 289944 121512 289950
rect 121460 289886 121512 289892
rect 121564 289882 121592 290391
rect 121552 289876 121604 289882
rect 121552 289818 121604 289824
rect 121460 289808 121512 289814
rect 121458 289776 121460 289785
rect 121512 289776 121514 289785
rect 121458 289711 121514 289720
rect 122010 289096 122066 289105
rect 122010 289031 122066 289040
rect 121550 288416 121606 288425
rect 121460 288380 121512 288386
rect 121550 288351 121606 288360
rect 121460 288322 121512 288328
rect 121472 287745 121500 288322
rect 121458 287736 121514 287745
rect 121458 287671 121514 287680
rect 121460 287632 121512 287638
rect 121460 287574 121512 287580
rect 121472 286385 121500 287574
rect 121564 287094 121592 288351
rect 121552 287088 121604 287094
rect 121552 287030 121604 287036
rect 121642 287056 121698 287065
rect 121642 286991 121698 287000
rect 121458 286376 121514 286385
rect 121458 286311 121514 286320
rect 121656 285802 121684 286991
rect 121644 285796 121696 285802
rect 121644 285738 121696 285744
rect 121460 285660 121512 285666
rect 121460 285602 121512 285608
rect 121472 284345 121500 285602
rect 121550 285016 121606 285025
rect 121550 284951 121606 284960
rect 121458 284336 121514 284345
rect 121458 284271 121514 284280
rect 121458 282976 121514 282985
rect 121458 282911 121460 282920
rect 121512 282911 121514 282920
rect 121460 282882 121512 282888
rect 121000 282192 121052 282198
rect 121000 282134 121052 282140
rect 121458 281616 121514 281625
rect 121458 281551 121460 281560
rect 121512 281551 121514 281560
rect 121460 281522 121512 281528
rect 121564 280838 121592 284951
rect 121552 280832 121604 280838
rect 121552 280774 121604 280780
rect 121458 280256 121514 280265
rect 121458 280191 121460 280200
rect 121512 280191 121514 280200
rect 121460 280162 121512 280168
rect 121550 279576 121606 279585
rect 121550 279511 121606 279520
rect 121458 278896 121514 278905
rect 121458 278831 121460 278840
rect 121512 278831 121514 278840
rect 121460 278802 121512 278808
rect 121564 278798 121592 279511
rect 121552 278792 121604 278798
rect 121552 278734 121604 278740
rect 121550 278216 121606 278225
rect 121550 278151 121606 278160
rect 121458 277536 121514 277545
rect 121564 277506 121592 278151
rect 121458 277471 121514 277480
rect 121552 277500 121604 277506
rect 121472 277438 121500 277471
rect 121552 277442 121604 277448
rect 121460 277432 121512 277438
rect 121460 277374 121512 277380
rect 122024 277394 122052 289031
rect 122116 285705 122144 311102
rect 122196 305040 122248 305046
rect 122196 304982 122248 304988
rect 122208 287638 122236 304982
rect 123484 299804 123536 299810
rect 123484 299746 123536 299752
rect 122196 287632 122248 287638
rect 122196 287574 122248 287580
rect 122102 285696 122158 285705
rect 122102 285631 122158 285640
rect 122378 280936 122434 280945
rect 122378 280871 122434 280880
rect 122024 277366 122236 277394
rect 121550 276856 121606 276865
rect 121550 276791 121606 276800
rect 121458 276176 121514 276185
rect 121564 276146 121592 276791
rect 121458 276111 121514 276120
rect 121552 276140 121604 276146
rect 121472 276078 121500 276111
rect 121552 276082 121604 276088
rect 121460 276072 121512 276078
rect 121460 276014 121512 276020
rect 121550 275496 121606 275505
rect 121550 275431 121606 275440
rect 121458 274816 121514 274825
rect 121458 274751 121460 274760
rect 121512 274751 121514 274760
rect 121460 274722 121512 274728
rect 121564 274718 121592 275431
rect 121552 274712 121604 274718
rect 121552 274654 121604 274660
rect 121460 274644 121512 274650
rect 121460 274586 121512 274592
rect 121472 274145 121500 274586
rect 121458 274136 121514 274145
rect 121458 274071 121514 274080
rect 121458 273456 121514 273465
rect 121458 273391 121514 273400
rect 121472 273290 121500 273391
rect 121460 273284 121512 273290
rect 121460 273226 121512 273232
rect 121000 272536 121052 272542
rect 121000 272478 121052 272484
rect 120908 242276 120960 242282
rect 120908 242218 120960 242224
rect 121012 237250 121040 272478
rect 121458 272096 121514 272105
rect 121458 272031 121460 272040
rect 121512 272031 121514 272040
rect 121460 272002 121512 272008
rect 121458 271416 121514 271425
rect 121458 271351 121514 271360
rect 121472 270570 121500 271351
rect 121460 270564 121512 270570
rect 121460 270506 121512 270512
rect 121550 270056 121606 270065
rect 121550 269991 121606 270000
rect 121458 269376 121514 269385
rect 121458 269311 121514 269320
rect 121472 269142 121500 269311
rect 121564 269210 121592 269991
rect 121552 269204 121604 269210
rect 121552 269146 121604 269152
rect 121460 269136 121512 269142
rect 121460 269078 121512 269084
rect 122102 267336 122158 267345
rect 122102 267271 122158 267280
rect 121458 266656 121514 266665
rect 121458 266591 121514 266600
rect 121472 266422 121500 266591
rect 121460 266416 121512 266422
rect 121460 266358 121512 266364
rect 121458 265976 121514 265985
rect 121458 265911 121514 265920
rect 121472 264994 121500 265911
rect 121460 264988 121512 264994
rect 121460 264930 121512 264936
rect 121550 264616 121606 264625
rect 121550 264551 121606 264560
rect 121458 263936 121514 263945
rect 121458 263871 121514 263880
rect 121472 263702 121500 263871
rect 121460 263696 121512 263702
rect 121460 263638 121512 263644
rect 121564 263634 121592 264551
rect 121552 263628 121604 263634
rect 121552 263570 121604 263576
rect 121460 263560 121512 263566
rect 121460 263502 121512 263508
rect 121472 263265 121500 263502
rect 121458 263256 121514 263265
rect 121458 263191 121514 263200
rect 121458 262576 121514 262585
rect 121458 262511 121514 262520
rect 121472 262274 121500 262511
rect 121460 262268 121512 262274
rect 121460 262210 121512 262216
rect 121550 261896 121606 261905
rect 121550 261831 121606 261840
rect 121460 261520 121512 261526
rect 121460 261462 121512 261468
rect 121472 261225 121500 261462
rect 121458 261216 121514 261225
rect 121458 261151 121514 261160
rect 121564 260914 121592 261831
rect 121552 260908 121604 260914
rect 121552 260850 121604 260856
rect 121550 260536 121606 260545
rect 121550 260471 121606 260480
rect 121458 259856 121514 259865
rect 121458 259791 121514 259800
rect 121472 259554 121500 259791
rect 121460 259548 121512 259554
rect 121460 259490 121512 259496
rect 121564 259486 121592 260471
rect 121552 259480 121604 259486
rect 121552 259422 121604 259428
rect 121550 259176 121606 259185
rect 121550 259111 121606 259120
rect 121458 258496 121514 258505
rect 121458 258431 121514 258440
rect 121472 258194 121500 258431
rect 121460 258188 121512 258194
rect 121460 258130 121512 258136
rect 121564 258126 121592 259111
rect 121552 258120 121604 258126
rect 121552 258062 121604 258068
rect 121550 257816 121606 257825
rect 121550 257751 121606 257760
rect 121458 257136 121514 257145
rect 121458 257071 121514 257080
rect 121472 256766 121500 257071
rect 121564 256834 121592 257751
rect 121552 256828 121604 256834
rect 121552 256770 121604 256776
rect 121460 256760 121512 256766
rect 121460 256702 121512 256708
rect 121550 256456 121606 256465
rect 121550 256391 121606 256400
rect 121458 255776 121514 255785
rect 121458 255711 121514 255720
rect 121472 255338 121500 255711
rect 121564 255406 121592 256391
rect 121552 255400 121604 255406
rect 121552 255342 121604 255348
rect 121460 255332 121512 255338
rect 121460 255274 121512 255280
rect 121458 254416 121514 254425
rect 121458 254351 121514 254360
rect 121472 253978 121500 254351
rect 121460 253972 121512 253978
rect 121460 253914 121512 253920
rect 121550 253736 121606 253745
rect 121550 253671 121606 253680
rect 121458 253056 121514 253065
rect 121458 252991 121514 253000
rect 121472 252618 121500 252991
rect 121564 252686 121592 253671
rect 121552 252680 121604 252686
rect 121552 252622 121604 252628
rect 121460 252612 121512 252618
rect 121460 252554 121512 252560
rect 121550 252376 121606 252385
rect 121550 252311 121606 252320
rect 121458 251696 121514 251705
rect 121458 251631 121514 251640
rect 121472 251326 121500 251631
rect 121460 251320 121512 251326
rect 121460 251262 121512 251268
rect 121564 251258 121592 252311
rect 121552 251252 121604 251258
rect 121552 251194 121604 251200
rect 121458 250336 121514 250345
rect 121458 250271 121514 250280
rect 121472 249830 121500 250271
rect 121460 249824 121512 249830
rect 121460 249766 121512 249772
rect 121458 248976 121514 248985
rect 121458 248911 121514 248920
rect 121472 248470 121500 248911
rect 121460 248464 121512 248470
rect 121460 248406 121512 248412
rect 121458 248296 121514 248305
rect 121458 248231 121514 248240
rect 121472 247110 121500 248231
rect 121460 247104 121512 247110
rect 121460 247046 121512 247052
rect 121550 246936 121606 246945
rect 121550 246871 121606 246880
rect 121458 246256 121514 246265
rect 121458 246191 121514 246200
rect 121472 245818 121500 246191
rect 121460 245812 121512 245818
rect 121460 245754 121512 245760
rect 121564 245750 121592 246871
rect 121552 245744 121604 245750
rect 121552 245686 121604 245692
rect 121550 245576 121606 245585
rect 121550 245511 121606 245520
rect 121458 244896 121514 244905
rect 121458 244831 121514 244840
rect 121472 244390 121500 244831
rect 121460 244384 121512 244390
rect 121460 244326 121512 244332
rect 121564 244322 121592 245511
rect 121552 244316 121604 244322
rect 121552 244258 121604 244264
rect 121460 244248 121512 244254
rect 121460 244190 121512 244196
rect 121550 244216 121606 244225
rect 121472 243545 121500 244190
rect 121550 244151 121606 244160
rect 121458 243536 121514 243545
rect 121458 243471 121514 243480
rect 121564 242962 121592 244151
rect 121552 242956 121604 242962
rect 121552 242898 121604 242904
rect 121644 242888 121696 242894
rect 121458 242856 121514 242865
rect 121644 242830 121696 242836
rect 121458 242791 121514 242800
rect 121472 242214 121500 242791
rect 121460 242208 121512 242214
rect 121656 242185 121684 242830
rect 121460 242150 121512 242156
rect 121642 242176 121698 242185
rect 121642 242111 121698 242120
rect 121458 240816 121514 240825
rect 121458 240751 121514 240760
rect 121472 240174 121500 240751
rect 121460 240168 121512 240174
rect 121460 240110 121512 240116
rect 121550 240136 121606 240145
rect 121550 240071 121606 240080
rect 121564 238950 121592 240071
rect 121552 238944 121604 238950
rect 121552 238886 121604 238892
rect 121000 237244 121052 237250
rect 121000 237186 121052 237192
rect 122116 232529 122144 267271
rect 122208 262886 122236 277366
rect 122286 272776 122342 272785
rect 122286 272711 122342 272720
rect 122196 262880 122248 262886
rect 122196 262822 122248 262828
rect 122300 247722 122328 272711
rect 122392 260166 122420 280871
rect 122380 260160 122432 260166
rect 122380 260102 122432 260108
rect 122288 247716 122340 247722
rect 122288 247658 122340 247664
rect 122102 232520 122158 232529
rect 122102 232455 122158 232464
rect 120816 192772 120868 192778
rect 120816 192714 120868 192720
rect 117964 189916 118016 189922
rect 117964 189858 118016 189864
rect 115848 185020 115900 185026
rect 115848 184962 115900 184968
rect 110696 182232 110748 182238
rect 110696 182174 110748 182180
rect 110236 179454 110288 179460
rect 110418 179480 110474 179489
rect 100666 177576 100722 177585
rect 100666 177511 100722 177520
rect 103426 177576 103482 177585
rect 103426 177511 103482 177520
rect 104624 177064 104676 177070
rect 110248 177041 110276 179454
rect 110418 179415 110474 179424
rect 104624 177006 104676 177012
rect 110234 177032 110290 177041
rect 104636 176769 104664 177006
rect 110234 176967 110290 176976
rect 108120 176860 108172 176866
rect 108120 176802 108172 176808
rect 107016 176792 107068 176798
rect 104622 176760 104678 176769
rect 104622 176695 104678 176704
rect 107014 176760 107016 176769
rect 108132 176769 108160 176802
rect 107068 176760 107070 176769
rect 107014 176695 107070 176704
rect 108118 176760 108174 176769
rect 108118 176695 108174 176704
rect 98368 176044 98420 176050
rect 98368 175986 98420 175992
rect 98380 175409 98408 175986
rect 110432 175982 110460 179415
rect 110708 177585 110736 182174
rect 112996 180940 113048 180946
rect 112996 180882 113048 180888
rect 113008 177585 113036 180882
rect 114376 179444 114428 179450
rect 114376 179386 114428 179392
rect 110694 177576 110750 177585
rect 110694 177511 110750 177520
rect 112994 177576 113050 177585
rect 112994 177511 113050 177520
rect 114388 177041 114416 179386
rect 115860 177585 115888 184962
rect 122748 184952 122800 184958
rect 122748 184894 122800 184900
rect 119988 183592 120040 183598
rect 119988 183534 120040 183540
rect 118424 178152 118476 178158
rect 118424 178094 118476 178100
rect 115846 177576 115902 177585
rect 115846 177511 115902 177520
rect 114374 177032 114430 177041
rect 114374 176967 114430 176976
rect 118436 176769 118464 178094
rect 120000 177585 120028 183534
rect 121092 181008 121144 181014
rect 121092 180950 121144 180956
rect 121104 177585 121132 180950
rect 119986 177576 120042 177585
rect 119986 177511 120042 177520
rect 121090 177576 121146 177585
rect 121090 177511 121146 177520
rect 122760 176769 122788 184894
rect 123496 182889 123524 299746
rect 124220 298784 124272 298790
rect 124220 298726 124272 298732
rect 123576 294364 123628 294370
rect 123576 294306 123628 294312
rect 123588 240825 123616 294306
rect 123668 285728 123720 285734
rect 123668 285670 123720 285676
rect 123574 240816 123630 240825
rect 123574 240751 123630 240760
rect 123680 235754 123708 285670
rect 124232 272542 124260 298726
rect 124864 298444 124916 298450
rect 124864 298386 124916 298392
rect 124220 272536 124272 272542
rect 124220 272478 124272 272484
rect 124128 245676 124180 245682
rect 124128 245618 124180 245624
rect 124140 242593 124168 245618
rect 124126 242584 124182 242593
rect 124126 242519 124182 242528
rect 123668 235748 123720 235754
rect 123668 235690 123720 235696
rect 124876 196858 124904 298386
rect 124968 251054 124996 347754
rect 125048 272060 125100 272066
rect 125048 272002 125100 272008
rect 124956 251048 125008 251054
rect 124956 250990 125008 250996
rect 124864 196852 124916 196858
rect 124864 196794 124916 196800
rect 123482 182880 123538 182889
rect 123482 182815 123538 182824
rect 125060 181665 125088 272002
rect 125140 269204 125192 269210
rect 125140 269146 125192 269152
rect 125152 222970 125180 269146
rect 125612 238746 125640 371826
rect 126624 371278 126652 371826
rect 126612 371272 126664 371278
rect 126612 371214 126664 371220
rect 144092 370524 144144 370530
rect 144092 370466 144144 370472
rect 144104 369918 144132 370466
rect 143540 369912 143592 369918
rect 143540 369854 143592 369860
rect 144092 369912 144144 369918
rect 144092 369854 144144 369860
rect 140044 368620 140096 368626
rect 140044 368562 140096 368568
rect 129004 364472 129056 364478
rect 129004 364414 129056 364420
rect 126244 360664 126296 360670
rect 126244 360606 126296 360612
rect 126256 288386 126284 360606
rect 126980 356720 127032 356726
rect 126980 356662 127032 356668
rect 126428 355020 126480 355026
rect 126428 354962 126480 354968
rect 126336 292868 126388 292874
rect 126336 292810 126388 292816
rect 126244 288380 126296 288386
rect 126244 288322 126296 288328
rect 126244 274780 126296 274786
rect 126244 274722 126296 274728
rect 125600 238740 125652 238746
rect 125600 238682 125652 238688
rect 125140 222964 125192 222970
rect 125140 222906 125192 222912
rect 126256 184414 126284 274722
rect 126348 202298 126376 292810
rect 126440 292534 126468 354962
rect 126428 292528 126480 292534
rect 126428 292470 126480 292476
rect 126428 247104 126480 247110
rect 126428 247046 126480 247052
rect 126336 202292 126388 202298
rect 126336 202234 126388 202240
rect 126440 190058 126468 247046
rect 126992 234462 127020 356662
rect 127622 295352 127678 295361
rect 127622 295287 127678 295296
rect 126980 234456 127032 234462
rect 126980 234398 127032 234404
rect 126428 190052 126480 190058
rect 126428 189994 126480 190000
rect 126888 186380 126940 186386
rect 126888 186322 126940 186328
rect 126244 184408 126296 184414
rect 126244 184350 126296 184356
rect 125046 181656 125102 181665
rect 125046 181591 125102 181600
rect 123024 178220 123076 178226
rect 123024 178162 123076 178168
rect 123036 176769 123064 178162
rect 126900 177585 126928 186322
rect 127636 184249 127664 295287
rect 127716 291304 127768 291310
rect 127716 291246 127768 291252
rect 127728 213314 127756 291246
rect 129016 235890 129044 364414
rect 130384 363044 130436 363050
rect 130384 362986 130436 362992
rect 129280 314696 129332 314702
rect 129280 314638 129332 314644
rect 129096 292800 129148 292806
rect 129096 292742 129148 292748
rect 129004 235884 129056 235890
rect 129004 235826 129056 235832
rect 127716 213308 127768 213314
rect 127716 213250 127768 213256
rect 129108 202366 129136 292742
rect 129188 291372 129240 291378
rect 129188 291314 129240 291320
rect 129200 203658 129228 291314
rect 129292 235686 129320 314638
rect 129648 297084 129700 297090
rect 129648 297026 129700 297032
rect 129660 296041 129688 297026
rect 129646 296032 129702 296041
rect 129646 295967 129702 295976
rect 129280 235680 129332 235686
rect 129280 235622 129332 235628
rect 129292 231810 129320 235622
rect 129280 231804 129332 231810
rect 129280 231746 129332 231752
rect 130396 229090 130424 362986
rect 138664 361956 138716 361962
rect 138664 361898 138716 361904
rect 134524 361888 134576 361894
rect 134524 361830 134576 361836
rect 130474 357504 130530 357513
rect 130474 357439 130530 357448
rect 130488 242894 130516 357439
rect 130568 301096 130620 301102
rect 130568 301038 130620 301044
rect 130476 242888 130528 242894
rect 130476 242830 130528 242836
rect 130384 229084 130436 229090
rect 130384 229026 130436 229032
rect 130580 213382 130608 301038
rect 131764 298240 131816 298246
rect 131764 298182 131816 298188
rect 130660 270564 130712 270570
rect 130660 270506 130712 270512
rect 130568 213376 130620 213382
rect 130568 213318 130620 213324
rect 129188 203652 129240 203658
rect 129188 203594 129240 203600
rect 129096 202360 129148 202366
rect 129096 202302 129148 202308
rect 130672 195498 130700 270506
rect 131776 204921 131804 298182
rect 133236 297016 133288 297022
rect 133236 296958 133288 296964
rect 133144 296948 133196 296954
rect 133144 296890 133196 296896
rect 131856 291236 131908 291242
rect 131856 291178 131908 291184
rect 131868 221610 131896 291178
rect 131948 249824 132000 249830
rect 131948 249766 132000 249772
rect 131856 221604 131908 221610
rect 131856 221546 131908 221552
rect 131762 204912 131818 204921
rect 131762 204847 131818 204856
rect 130660 195492 130712 195498
rect 130660 195434 130712 195440
rect 131960 185910 131988 249766
rect 133156 191049 133184 296890
rect 133248 198150 133276 296958
rect 133328 277500 133380 277506
rect 133328 277442 133380 277448
rect 133340 226234 133368 277442
rect 134536 233102 134564 361830
rect 135904 357536 135956 357542
rect 135904 357478 135956 357484
rect 134708 302456 134760 302462
rect 134708 302398 134760 302404
rect 134616 292732 134668 292738
rect 134616 292674 134668 292680
rect 134524 233096 134576 233102
rect 134524 233038 134576 233044
rect 133328 226228 133380 226234
rect 133328 226170 133380 226176
rect 133236 198144 133288 198150
rect 133236 198086 133288 198092
rect 134628 194070 134656 292674
rect 134720 204950 134748 302398
rect 135916 231606 135944 357478
rect 136088 299736 136140 299742
rect 136088 299678 136140 299684
rect 135996 294432 136048 294438
rect 135996 294374 136048 294380
rect 135904 231600 135956 231606
rect 135904 231542 135956 231548
rect 134708 204944 134760 204950
rect 134708 204886 134760 204892
rect 134616 194064 134668 194070
rect 134616 194006 134668 194012
rect 133142 191040 133198 191049
rect 133142 190975 133198 190984
rect 136008 188358 136036 294374
rect 136100 209234 136128 299678
rect 137284 298376 137336 298382
rect 137284 298318 137336 298324
rect 136180 263696 136232 263702
rect 136180 263638 136232 263644
rect 136088 209228 136140 209234
rect 136088 209170 136140 209176
rect 136192 200938 136220 263638
rect 137296 210594 137324 298318
rect 137376 295588 137428 295594
rect 137376 295530 137428 295536
rect 137388 228886 137416 295530
rect 137468 251320 137520 251326
rect 137468 251262 137520 251268
rect 137376 228880 137428 228886
rect 137376 228822 137428 228828
rect 137480 218754 137508 251262
rect 138676 238406 138704 361898
rect 138756 305176 138808 305182
rect 138756 305118 138808 305124
rect 138664 238400 138716 238406
rect 138664 238342 138716 238348
rect 137468 218748 137520 218754
rect 137468 218690 137520 218696
rect 137284 210588 137336 210594
rect 137284 210530 137336 210536
rect 136180 200932 136232 200938
rect 136180 200874 136232 200880
rect 138768 192574 138796 305118
rect 138848 294160 138900 294166
rect 138848 294102 138900 294108
rect 138756 192568 138808 192574
rect 138756 192510 138808 192516
rect 138860 188494 138888 294102
rect 138940 280220 138992 280226
rect 138940 280162 138992 280168
rect 138952 198218 138980 280162
rect 140056 244254 140084 368562
rect 142804 359032 142856 359038
rect 142804 358974 142856 358980
rect 140228 296812 140280 296818
rect 140228 296754 140280 296760
rect 140136 294296 140188 294302
rect 140136 294238 140188 294244
rect 140044 244248 140096 244254
rect 140044 244190 140096 244196
rect 140148 234054 140176 294238
rect 140240 263022 140268 296754
rect 141516 292596 141568 292602
rect 141516 292538 141568 292544
rect 141424 273284 141476 273290
rect 141424 273226 141476 273232
rect 140688 269816 140740 269822
rect 140688 269758 140740 269764
rect 140228 263016 140280 263022
rect 140228 262958 140280 262964
rect 140228 245812 140280 245818
rect 140228 245754 140280 245760
rect 140136 234048 140188 234054
rect 140136 233990 140188 233996
rect 140240 200870 140268 245754
rect 140700 237318 140728 269758
rect 140688 237312 140740 237318
rect 140688 237254 140740 237260
rect 141436 221678 141464 273226
rect 141528 240786 141556 292538
rect 141608 262268 141660 262274
rect 141608 262210 141660 262216
rect 141516 240780 141568 240786
rect 141516 240722 141568 240728
rect 141424 221672 141476 221678
rect 141424 221614 141476 221620
rect 141620 216170 141648 262210
rect 142816 238882 142844 358974
rect 142896 303680 142948 303686
rect 142896 303622 142948 303628
rect 142804 238876 142856 238882
rect 142804 238818 142856 238824
rect 141608 216164 141660 216170
rect 141608 216106 141660 216112
rect 142908 210730 142936 303622
rect 142988 282940 143040 282946
rect 142988 282882 143040 282888
rect 142896 210724 142948 210730
rect 142896 210666 142948 210672
rect 140228 200864 140280 200870
rect 140228 200806 140280 200812
rect 138940 198212 138992 198218
rect 138940 198154 138992 198160
rect 143000 191214 143028 282882
rect 143080 269136 143132 269142
rect 143080 269078 143132 269084
rect 143092 206582 143120 269078
rect 143552 261526 143580 369854
rect 146944 369164 146996 369170
rect 146944 369106 146996 369112
rect 146956 368694 146984 369106
rect 146944 368688 146996 368694
rect 146944 368630 146996 368636
rect 144184 301232 144236 301238
rect 144184 301174 144236 301180
rect 143540 261520 143592 261526
rect 143540 261462 143592 261468
rect 144196 209370 144224 301174
rect 144368 299600 144420 299606
rect 144368 299542 144420 299548
rect 144276 256828 144328 256834
rect 144276 256770 144328 256776
rect 144184 209364 144236 209370
rect 144184 209306 144236 209312
rect 143080 206576 143132 206582
rect 143080 206518 143132 206524
rect 142988 191208 143040 191214
rect 142988 191150 143040 191156
rect 138848 188488 138900 188494
rect 138848 188430 138900 188436
rect 144288 188426 144316 256770
rect 144380 233102 144408 299542
rect 145564 295520 145616 295526
rect 145564 295462 145616 295468
rect 144460 261520 144512 261526
rect 144460 261462 144512 261468
rect 144368 233096 144420 233102
rect 144368 233038 144420 233044
rect 144472 220794 144500 261462
rect 144460 220788 144512 220794
rect 144460 220730 144512 220736
rect 145576 203794 145604 295462
rect 145654 291952 145710 291961
rect 145654 291887 145710 291896
rect 145668 227633 145696 291887
rect 145748 274712 145800 274718
rect 145748 274654 145800 274660
rect 145654 227624 145710 227633
rect 145654 227559 145710 227568
rect 145760 223446 145788 274654
rect 146956 263566 146984 368630
rect 148324 302388 148376 302394
rect 148324 302330 148376 302336
rect 147036 291848 147088 291854
rect 147036 291790 147088 291796
rect 146944 263560 146996 263566
rect 146944 263502 146996 263508
rect 146956 262954 146984 263502
rect 146944 262948 146996 262954
rect 146944 262890 146996 262896
rect 146944 259548 146996 259554
rect 146944 259490 146996 259496
rect 145748 223440 145800 223446
rect 145748 223382 145800 223388
rect 145564 203788 145616 203794
rect 145564 203730 145616 203736
rect 144276 188420 144328 188426
rect 144276 188362 144328 188368
rect 135996 188352 136048 188358
rect 135996 188294 136048 188300
rect 131948 185904 132000 185910
rect 131948 185846 132000 185852
rect 127622 184240 127678 184249
rect 127622 184175 127678 184184
rect 130752 182300 130804 182306
rect 130752 182242 130804 182248
rect 128084 180872 128136 180878
rect 128084 180814 128136 180820
rect 128096 177585 128124 180814
rect 129464 178084 129516 178090
rect 129464 178026 129516 178032
rect 126886 177576 126942 177585
rect 126886 177511 126942 177520
rect 128082 177576 128138 177585
rect 128082 177511 128138 177520
rect 128176 176928 128228 176934
rect 128176 176870 128228 176876
rect 128188 176769 128216 176870
rect 129476 176769 129504 178026
rect 130764 177585 130792 182242
rect 132040 179580 132092 179586
rect 132040 179522 132092 179528
rect 130750 177576 130806 177585
rect 130750 177511 130806 177520
rect 132052 177041 132080 179522
rect 146956 178702 146984 259490
rect 147048 202434 147076 291790
rect 147220 276140 147272 276146
rect 147220 276082 147272 276088
rect 147128 245744 147180 245750
rect 147128 245686 147180 245692
rect 147036 202428 147088 202434
rect 147036 202370 147088 202376
rect 147140 194138 147168 245686
rect 147232 226273 147260 276082
rect 147218 226264 147274 226273
rect 147218 226199 147274 226208
rect 147128 194132 147180 194138
rect 147128 194074 147180 194080
rect 148336 192846 148364 302330
rect 148416 299668 148468 299674
rect 148416 299610 148468 299616
rect 148428 238882 148456 299610
rect 149716 299441 149744 700334
rect 153212 380186 153240 702406
rect 170324 700398 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 170312 700392 170364 700398
rect 170312 700334 170364 700340
rect 193220 700324 193272 700330
rect 193220 700266 193272 700272
rect 179052 697604 179104 697610
rect 179052 697546 179104 697552
rect 153200 380180 153252 380186
rect 153200 380122 153252 380128
rect 170956 368552 171008 368558
rect 170956 368494 171008 368500
rect 152462 365800 152518 365809
rect 152462 365735 152518 365744
rect 151728 325712 151780 325718
rect 151728 325654 151780 325660
rect 149796 301164 149848 301170
rect 149796 301106 149848 301112
rect 149702 299432 149758 299441
rect 149702 299367 149758 299376
rect 149704 289944 149756 289950
rect 149704 289886 149756 289892
rect 148508 258188 148560 258194
rect 148508 258130 148560 258136
rect 148416 238876 148468 238882
rect 148416 238818 148468 238824
rect 148520 224874 148548 258130
rect 148600 240168 148652 240174
rect 148600 240110 148652 240116
rect 148508 224868 148560 224874
rect 148508 224810 148560 224816
rect 148612 212022 148640 240110
rect 148968 238944 149020 238950
rect 148968 238886 149020 238892
rect 148980 233918 149008 238886
rect 148968 233912 149020 233918
rect 148968 233854 149020 233860
rect 148600 212016 148652 212022
rect 148600 211958 148652 211964
rect 149716 207874 149744 289886
rect 149704 207868 149756 207874
rect 149704 207810 149756 207816
rect 149808 203726 149836 301106
rect 151176 295724 151228 295730
rect 151176 295666 151228 295672
rect 151084 278860 151136 278866
rect 151084 278802 151136 278808
rect 149888 255400 149940 255406
rect 149888 255342 149940 255348
rect 149900 231606 149928 255342
rect 149980 242276 150032 242282
rect 149980 242218 150032 242224
rect 149888 231600 149940 231606
rect 149888 231542 149940 231548
rect 149992 224942 150020 242218
rect 149980 224936 150032 224942
rect 149980 224878 150032 224884
rect 148416 203720 148468 203726
rect 148416 203662 148468 203668
rect 149796 203720 149848 203726
rect 149796 203662 149848 203668
rect 148324 192840 148376 192846
rect 148324 192782 148376 192788
rect 148428 184346 148456 203662
rect 151096 198286 151124 278802
rect 151188 221474 151216 295666
rect 151740 230450 151768 325654
rect 152476 235618 152504 365735
rect 162308 364540 162360 364546
rect 162308 364482 162360 364488
rect 158628 357808 158680 357814
rect 158628 357750 158680 357756
rect 154488 357604 154540 357610
rect 154488 357546 154540 357552
rect 154396 307080 154448 307086
rect 154396 307022 154448 307028
rect 154408 306406 154436 307022
rect 154396 306400 154448 306406
rect 154396 306342 154448 306348
rect 152556 302320 152608 302326
rect 152556 302262 152608 302268
rect 152464 235612 152516 235618
rect 152464 235554 152516 235560
rect 151728 230444 151780 230450
rect 151728 230386 151780 230392
rect 151740 229838 151768 230386
rect 151728 229832 151780 229838
rect 151728 229774 151780 229780
rect 151176 221468 151228 221474
rect 151176 221410 151228 221416
rect 151084 198280 151136 198286
rect 151084 198222 151136 198228
rect 152568 189990 152596 302262
rect 153844 301028 153896 301034
rect 153844 300970 153896 300976
rect 153108 286340 153160 286346
rect 153108 286282 153160 286288
rect 153120 285802 153148 286282
rect 153108 285796 153160 285802
rect 153108 285738 153160 285744
rect 152648 252680 152700 252686
rect 152648 252622 152700 252628
rect 152660 196926 152688 252622
rect 153120 218006 153148 285738
rect 153856 223514 153884 300970
rect 153936 259480 153988 259486
rect 153936 259422 153988 259428
rect 153844 223508 153896 223514
rect 153844 223450 153896 223456
rect 153948 219434 153976 259422
rect 154408 235890 154436 306342
rect 154396 235884 154448 235890
rect 154396 235826 154448 235832
rect 153936 219428 153988 219434
rect 153936 219370 153988 219376
rect 153844 218816 153896 218822
rect 153844 218758 153896 218764
rect 153108 218000 153160 218006
rect 153108 217942 153160 217948
rect 152648 196920 152700 196926
rect 152648 196862 152700 196868
rect 153856 195294 153884 218758
rect 153844 195288 153896 195294
rect 153844 195230 153896 195236
rect 152556 189984 152608 189990
rect 152556 189926 152608 189932
rect 148416 184340 148468 184346
rect 148416 184282 148468 184288
rect 154500 181490 154528 357546
rect 157248 345092 157300 345098
rect 157248 345034 157300 345040
rect 155224 300960 155276 300966
rect 155224 300902 155276 300908
rect 155236 214810 155264 300902
rect 156696 296880 156748 296886
rect 156696 296822 156748 296828
rect 156604 295384 156656 295390
rect 156604 295326 156656 295332
rect 155868 283620 155920 283626
rect 155868 283562 155920 283568
rect 155880 282946 155908 283562
rect 155868 282940 155920 282946
rect 155868 282882 155920 282888
rect 155316 260908 155368 260914
rect 155316 260850 155368 260856
rect 155328 232558 155356 260850
rect 155316 232552 155368 232558
rect 155316 232494 155368 232500
rect 155880 219366 155908 282882
rect 156512 257372 156564 257378
rect 156512 257314 156564 257320
rect 156524 257281 156552 257314
rect 156510 257272 156566 257281
rect 156510 257207 156566 257216
rect 155868 219360 155920 219366
rect 155868 219302 155920 219308
rect 155224 214804 155276 214810
rect 155224 214746 155276 214752
rect 156616 188562 156644 295326
rect 156708 220726 156736 296822
rect 157156 281512 157208 281518
rect 157156 281454 157208 281460
rect 157168 280226 157196 281454
rect 157156 280220 157208 280226
rect 157156 280162 157208 280168
rect 157168 237250 157196 280162
rect 157260 237289 157288 345034
rect 158444 297424 158496 297430
rect 158444 297366 158496 297372
rect 158456 297090 158484 297366
rect 158444 297084 158496 297090
rect 158444 297026 158496 297032
rect 158456 296857 158484 297026
rect 158442 296848 158498 296857
rect 158442 296783 158498 296792
rect 157340 296744 157392 296750
rect 157340 296686 157392 296692
rect 157352 281518 157380 296686
rect 157984 281580 158036 281586
rect 157984 281522 158036 281528
rect 157340 281512 157392 281518
rect 157340 281454 157392 281460
rect 157338 254280 157394 254289
rect 157338 254215 157394 254224
rect 157352 254046 157380 254215
rect 157340 254040 157392 254046
rect 157340 253982 157392 253988
rect 157246 237280 157302 237289
rect 157156 237244 157208 237250
rect 157246 237215 157302 237224
rect 157156 237186 157208 237192
rect 157260 233170 157288 237215
rect 157248 233164 157300 233170
rect 157248 233106 157300 233112
rect 156696 220720 156748 220726
rect 156696 220662 156748 220668
rect 156604 188556 156656 188562
rect 156604 188498 156656 188504
rect 154488 181484 154540 181490
rect 154488 181426 154540 181432
rect 146944 178696 146996 178702
rect 146944 178638 146996 178644
rect 148232 178288 148284 178294
rect 148232 178230 148284 178236
rect 132038 177032 132094 177041
rect 132038 176967 132094 176976
rect 133144 176996 133196 177002
rect 133144 176938 133196 176944
rect 133156 176769 133184 176938
rect 148244 176769 148272 178230
rect 157996 177313 158024 281522
rect 158536 278860 158588 278866
rect 158536 278802 158588 278808
rect 158444 254040 158496 254046
rect 158444 253982 158496 253988
rect 158456 230382 158484 253982
rect 158444 230376 158496 230382
rect 158444 230318 158496 230324
rect 158548 226166 158576 278802
rect 158536 226160 158588 226166
rect 158536 226102 158588 226108
rect 158640 180266 158668 357750
rect 160744 340944 160796 340950
rect 160744 340886 160796 340892
rect 160560 312588 160612 312594
rect 160560 312530 160612 312536
rect 160572 311953 160600 312530
rect 160558 311944 160614 311953
rect 160558 311879 160560 311888
rect 160612 311879 160614 311888
rect 160560 311850 160612 311856
rect 160572 311819 160600 311850
rect 160756 311166 160784 340886
rect 160744 311160 160796 311166
rect 160744 311102 160796 311108
rect 162124 305108 162176 305114
rect 162124 305050 162176 305056
rect 160008 300960 160060 300966
rect 160008 300902 160060 300908
rect 159364 298172 159416 298178
rect 159364 298114 159416 298120
rect 158720 282192 158772 282198
rect 158720 282134 158772 282140
rect 158732 281586 158760 282134
rect 158720 281580 158772 281586
rect 158720 281522 158772 281528
rect 159376 202162 159404 298114
rect 159916 281580 159968 281586
rect 159916 281522 159968 281528
rect 159456 255332 159508 255338
rect 159456 255274 159508 255280
rect 159468 231849 159496 255274
rect 159928 240106 159956 281522
rect 159916 240100 159968 240106
rect 159916 240042 159968 240048
rect 159454 231840 159510 231849
rect 159454 231775 159510 231784
rect 159364 202156 159416 202162
rect 159364 202098 159416 202104
rect 160020 184482 160048 300902
rect 160744 291848 160796 291854
rect 160744 291790 160796 291796
rect 160100 272536 160152 272542
rect 160100 272478 160152 272484
rect 160112 271930 160140 272478
rect 160100 271924 160152 271930
rect 160100 271866 160152 271872
rect 160098 244896 160154 244905
rect 160098 244831 160154 244840
rect 160112 244390 160140 244831
rect 160100 244384 160152 244390
rect 160100 244326 160152 244332
rect 160756 242214 160784 291790
rect 161204 271924 161256 271930
rect 161204 271866 161256 271872
rect 160744 242208 160796 242214
rect 160744 242150 160796 242156
rect 160756 227662 160784 242150
rect 161216 241466 161244 271866
rect 161388 267776 161440 267782
rect 161388 267718 161440 267724
rect 161294 244896 161350 244905
rect 161294 244831 161350 244840
rect 161204 241460 161256 241466
rect 161204 241402 161256 241408
rect 160744 227656 160796 227662
rect 160744 227598 160796 227604
rect 160744 225684 160796 225690
rect 160744 225626 160796 225632
rect 160756 218822 160784 225626
rect 160744 218816 160796 218822
rect 160744 218758 160796 218764
rect 161308 213897 161336 244831
rect 161294 213888 161350 213897
rect 161294 213823 161350 213832
rect 160100 201000 160152 201006
rect 160100 200942 160152 200948
rect 160112 195430 160140 200942
rect 160100 195424 160152 195430
rect 160100 195366 160152 195372
rect 160744 193996 160796 194002
rect 160744 193938 160796 193944
rect 160008 184476 160060 184482
rect 160008 184418 160060 184424
rect 158628 180260 158680 180266
rect 158628 180202 158680 180208
rect 157982 177304 158038 177313
rect 157982 177239 158038 177248
rect 118422 176760 118478 176769
rect 118422 176695 118478 176704
rect 122746 176760 122802 176769
rect 122746 176695 122802 176704
rect 123022 176760 123078 176769
rect 123022 176695 123078 176704
rect 128174 176760 128230 176769
rect 128174 176695 128230 176704
rect 129462 176760 129518 176769
rect 129462 176695 129518 176704
rect 133142 176760 133198 176769
rect 133142 176695 133198 176704
rect 135718 176760 135774 176769
rect 135718 176695 135774 176704
rect 148230 176760 148286 176769
rect 148230 176695 148286 176704
rect 158994 176760 159050 176769
rect 158994 176695 158996 176704
rect 135732 176662 135760 176695
rect 159048 176695 159050 176704
rect 158996 176666 159048 176672
rect 135720 176656 135772 176662
rect 135720 176598 135772 176604
rect 134432 176248 134484 176254
rect 134432 176190 134484 176196
rect 124496 176180 124548 176186
rect 124496 176122 124548 176128
rect 116952 176112 117004 176118
rect 116952 176054 117004 176060
rect 110420 175976 110472 175982
rect 110420 175918 110472 175924
rect 116964 175681 116992 176054
rect 124508 175681 124536 176122
rect 134444 175681 134472 176190
rect 160756 175982 160784 193938
rect 161400 187202 161428 267718
rect 162136 205222 162164 305050
rect 162216 292664 162268 292670
rect 162216 292606 162268 292612
rect 162124 205216 162176 205222
rect 162124 205158 162176 205164
rect 162228 199578 162256 292606
rect 162320 289814 162348 364482
rect 166264 363112 166316 363118
rect 166264 363054 166316 363060
rect 164148 357740 164200 357746
rect 164148 357682 164200 357688
rect 162308 289808 162360 289814
rect 162308 289750 162360 289756
rect 162768 285728 162820 285734
rect 162768 285670 162820 285676
rect 162308 263016 162360 263022
rect 162308 262958 162360 262964
rect 162320 261526 162348 262958
rect 162308 261520 162360 261526
rect 162308 261462 162360 261468
rect 162676 261520 162728 261526
rect 162676 261462 162728 261468
rect 162306 229800 162362 229809
rect 162306 229735 162362 229744
rect 162320 222086 162348 229735
rect 162688 229090 162716 261462
rect 162780 235754 162808 285670
rect 163504 277432 163556 277438
rect 163504 277374 163556 277380
rect 162768 235748 162820 235754
rect 162768 235690 162820 235696
rect 162676 229084 162728 229090
rect 162676 229026 162728 229032
rect 162308 222080 162360 222086
rect 162308 222022 162360 222028
rect 162768 218884 162820 218890
rect 162768 218826 162820 218832
rect 162780 215286 162808 218826
rect 162768 215280 162820 215286
rect 162768 215222 162820 215228
rect 162308 209432 162360 209438
rect 162308 209374 162360 209380
rect 162216 199572 162268 199578
rect 162216 199514 162268 199520
rect 161388 187196 161440 187202
rect 161388 187138 161440 187144
rect 162320 187066 162348 209374
rect 163516 191350 163544 277374
rect 163596 263628 163648 263634
rect 163596 263570 163648 263576
rect 163608 230246 163636 263570
rect 163596 230240 163648 230246
rect 163596 230182 163648 230188
rect 163504 191344 163556 191350
rect 163504 191286 163556 191292
rect 162308 187060 162360 187066
rect 162308 187002 162360 187008
rect 164160 180033 164188 357682
rect 165068 300892 165120 300898
rect 165068 300834 165120 300840
rect 164976 295656 165028 295662
rect 164976 295598 165028 295604
rect 164884 289876 164936 289882
rect 164884 289818 164936 289824
rect 164146 180024 164202 180033
rect 164146 179959 164202 179968
rect 164896 177410 164924 289818
rect 164988 189689 165016 295598
rect 165080 241233 165108 300834
rect 166276 274650 166304 363054
rect 169116 298308 169168 298314
rect 169116 298250 169168 298256
rect 169024 289876 169076 289882
rect 169024 289818 169076 289824
rect 167736 287088 167788 287094
rect 167736 287030 167788 287036
rect 166264 274644 166316 274650
rect 166264 274586 166316 274592
rect 166448 266416 166500 266422
rect 165618 266384 165674 266393
rect 166448 266358 166500 266364
rect 165618 266319 165620 266328
rect 165672 266319 165674 266328
rect 165620 266290 165672 266296
rect 166264 264988 166316 264994
rect 166264 264930 166316 264936
rect 165160 260160 165212 260166
rect 165160 260102 165212 260108
rect 165066 241224 165122 241233
rect 165066 241159 165122 241168
rect 165172 222902 165200 260102
rect 165160 222896 165212 222902
rect 165160 222838 165212 222844
rect 166172 210656 166224 210662
rect 166172 210598 166224 210604
rect 166184 205086 166212 210598
rect 166172 205080 166224 205086
rect 166172 205022 166224 205028
rect 164974 189680 165030 189689
rect 164974 189615 165030 189624
rect 165344 179580 165396 179586
rect 165344 179522 165396 179528
rect 164884 177404 164936 177410
rect 164884 177346 164936 177352
rect 164516 176996 164568 177002
rect 164516 176938 164568 176944
rect 160744 175976 160796 175982
rect 160744 175918 160796 175924
rect 116950 175672 117006 175681
rect 116950 175607 117006 175616
rect 124494 175672 124550 175681
rect 124494 175607 124550 175616
rect 134430 175672 134486 175681
rect 134430 175607 134486 175616
rect 98366 175400 98422 175409
rect 98366 175335 98422 175344
rect 164528 175234 164556 176938
rect 164516 175228 164568 175234
rect 164516 175170 164568 175176
rect 67638 128072 67694 128081
rect 67638 128007 67694 128016
rect 67454 120864 67510 120873
rect 67454 120799 67510 120808
rect 67468 90953 67496 120799
rect 67652 93838 67680 128007
rect 67730 100736 67786 100745
rect 67730 100671 67786 100680
rect 67640 93832 67692 93838
rect 67640 93774 67692 93780
rect 67454 90944 67510 90953
rect 67454 90879 67510 90888
rect 67744 86970 67772 100671
rect 165356 173874 165384 179522
rect 166276 178809 166304 264930
rect 166356 242956 166408 242962
rect 166356 242898 166408 242904
rect 166262 178800 166318 178809
rect 166262 178735 166318 178744
rect 166368 177342 166396 242898
rect 166460 229906 166488 266358
rect 166908 259480 166960 259486
rect 166908 259422 166960 259428
rect 166448 229900 166500 229906
rect 166448 229842 166500 229848
rect 166540 181008 166592 181014
rect 166540 180950 166592 180956
rect 166448 178288 166500 178294
rect 166448 178230 166500 178236
rect 166356 177336 166408 177342
rect 166356 177278 166408 177284
rect 165436 176928 165488 176934
rect 165436 176870 165488 176876
rect 165448 174554 165476 176870
rect 166264 176724 166316 176730
rect 166264 176666 166316 176672
rect 165528 176248 165580 176254
rect 165528 176190 165580 176196
rect 165540 175166 165568 176190
rect 165528 175160 165580 175166
rect 165528 175102 165580 175108
rect 165436 174548 165488 174554
rect 165436 174490 165488 174496
rect 165344 173868 165396 173874
rect 165344 173810 165396 173816
rect 166276 149054 166304 176666
rect 166460 150414 166488 178230
rect 166552 168366 166580 180950
rect 166920 180334 166948 259422
rect 167644 258120 167696 258126
rect 167644 258062 167696 258068
rect 167000 247716 167052 247722
rect 167000 247658 167052 247664
rect 167012 239970 167040 247658
rect 167000 239964 167052 239970
rect 167000 239906 167052 239912
rect 167656 182918 167684 258062
rect 167748 228954 167776 287030
rect 167828 280832 167880 280838
rect 167828 280774 167880 280780
rect 167840 236706 167868 280774
rect 169036 269822 169064 289818
rect 169128 280838 169156 298250
rect 170968 298110 170996 368494
rect 175096 367124 175148 367130
rect 175096 367066 175148 367072
rect 171784 366444 171836 366450
rect 171784 366386 171836 366392
rect 171048 356380 171100 356386
rect 171048 356322 171100 356328
rect 169760 298104 169812 298110
rect 169760 298046 169812 298052
rect 170956 298104 171008 298110
rect 170956 298046 171008 298052
rect 169772 297401 169800 298046
rect 169758 297392 169814 297401
rect 169758 297327 169814 297336
rect 170494 293992 170550 294001
rect 170494 293927 170550 293936
rect 169116 280832 169168 280838
rect 169116 280774 169168 280780
rect 169024 269816 169076 269822
rect 169024 269758 169076 269764
rect 169116 262948 169168 262954
rect 169116 262890 169168 262896
rect 169024 262880 169076 262886
rect 169024 262822 169076 262828
rect 168378 242176 168434 242185
rect 168378 242111 168434 242120
rect 168392 241534 168420 242111
rect 168380 241528 168432 241534
rect 168380 241470 168432 241476
rect 167828 236700 167880 236706
rect 167828 236642 167880 236648
rect 167736 228948 167788 228954
rect 167736 228890 167788 228896
rect 169036 217326 169064 262822
rect 169128 236774 169156 262890
rect 170404 252612 170456 252618
rect 170404 252554 170456 252560
rect 169668 241528 169720 241534
rect 169668 241470 169720 241476
rect 169116 236768 169168 236774
rect 169116 236710 169168 236716
rect 169680 230450 169708 241470
rect 169668 230444 169720 230450
rect 169668 230386 169720 230392
rect 169024 217320 169076 217326
rect 169024 217262 169076 217268
rect 167736 205148 167788 205154
rect 167736 205090 167788 205096
rect 167748 184385 167776 205090
rect 169116 186380 169168 186386
rect 169116 186322 169168 186328
rect 167734 184376 167790 184385
rect 167734 184311 167790 184320
rect 167644 182912 167696 182918
rect 167644 182854 167696 182860
rect 167736 180940 167788 180946
rect 167736 180882 167788 180888
rect 166908 180328 166960 180334
rect 166908 180270 166960 180276
rect 166632 178152 166684 178158
rect 166632 178094 166684 178100
rect 166540 168360 166592 168366
rect 166540 168302 166592 168308
rect 166644 167006 166672 178094
rect 166998 176896 167054 176905
rect 166998 176831 167054 176840
rect 167012 171834 167040 176831
rect 167000 171828 167052 171834
rect 167000 171770 167052 171776
rect 167642 171592 167698 171601
rect 167642 171527 167698 171536
rect 166632 167000 166684 167006
rect 166632 166942 166684 166948
rect 167656 151094 167684 171527
rect 167748 164218 167776 180882
rect 167828 179512 167880 179518
rect 167828 179454 167880 179460
rect 167736 164212 167788 164218
rect 167736 164154 167788 164160
rect 167840 162858 167868 179454
rect 169024 176860 169076 176866
rect 169024 176802 169076 176808
rect 167920 176180 167972 176186
rect 167920 176122 167972 176128
rect 167932 169726 167960 176122
rect 167920 169720 167972 169726
rect 167920 169662 167972 169668
rect 167828 162852 167880 162858
rect 167828 162794 167880 162800
rect 169036 161430 169064 176802
rect 169128 171086 169156 186322
rect 170416 185842 170444 252554
rect 170508 232626 170536 293927
rect 170588 276072 170640 276078
rect 170588 276014 170640 276020
rect 170496 232620 170548 232626
rect 170496 232562 170548 232568
rect 170600 225690 170628 276014
rect 170588 225684 170640 225690
rect 170588 225626 170640 225632
rect 170404 185836 170456 185842
rect 170404 185778 170456 185784
rect 170496 185020 170548 185026
rect 170496 184962 170548 184968
rect 169300 178220 169352 178226
rect 169300 178162 169352 178168
rect 169208 176112 169260 176118
rect 169208 176054 169260 176060
rect 169116 171080 169168 171086
rect 169116 171022 169168 171028
rect 169220 166938 169248 176054
rect 169312 169658 169340 178162
rect 170404 176044 170456 176050
rect 170404 175986 170456 175992
rect 169300 169652 169352 169658
rect 169300 169594 169352 169600
rect 169208 166932 169260 166938
rect 169208 166874 169260 166880
rect 169024 161424 169076 161430
rect 169024 161366 169076 161372
rect 170416 155922 170444 175986
rect 170508 165578 170536 184962
rect 170680 183592 170732 183598
rect 170680 183534 170732 183540
rect 170588 177064 170640 177070
rect 170588 177006 170640 177012
rect 170496 165572 170548 165578
rect 170496 165514 170548 165520
rect 170600 160070 170628 177006
rect 170692 166870 170720 183534
rect 171060 177546 171088 356322
rect 171140 295452 171192 295458
rect 171140 295394 171192 295400
rect 171152 278866 171180 295394
rect 171796 286346 171824 366386
rect 172428 359168 172480 359174
rect 172428 359110 172480 359116
rect 171784 286340 171836 286346
rect 171784 286282 171836 286288
rect 171140 278860 171192 278866
rect 171140 278802 171192 278808
rect 171784 278792 171836 278798
rect 171784 278734 171836 278740
rect 171796 189854 171824 278734
rect 172336 276072 172388 276078
rect 172336 276014 172388 276020
rect 171876 253972 171928 253978
rect 171876 253914 171928 253920
rect 171784 189848 171836 189854
rect 171784 189790 171836 189796
rect 171784 187740 171836 187746
rect 171784 187682 171836 187688
rect 171048 177540 171100 177546
rect 171048 177482 171100 177488
rect 170680 166864 170732 166870
rect 170680 166806 170732 166812
rect 170588 160064 170640 160070
rect 170588 160006 170640 160012
rect 171796 157350 171824 187682
rect 171888 181558 171916 253914
rect 172348 238746 172376 276014
rect 172336 238740 172388 238746
rect 172336 238682 172388 238688
rect 171968 189100 172020 189106
rect 171968 189042 172020 189048
rect 171876 181552 171928 181558
rect 171876 181494 171928 181500
rect 171876 176792 171928 176798
rect 171876 176734 171928 176740
rect 171888 161362 171916 176734
rect 171876 161356 171928 161362
rect 171876 161298 171928 161304
rect 171980 158710 172008 189042
rect 172334 160168 172390 160177
rect 172334 160103 172390 160112
rect 171968 158704 172020 158710
rect 171968 158646 172020 158652
rect 171784 157344 171836 157350
rect 171784 157286 171836 157292
rect 170404 155916 170456 155922
rect 170404 155858 170456 155864
rect 171784 151836 171836 151842
rect 171784 151778 171836 151784
rect 167644 151088 167696 151094
rect 167644 151030 167696 151036
rect 166448 150408 166500 150414
rect 166448 150350 166500 150356
rect 166264 149048 166316 149054
rect 166264 148990 166316 148996
rect 166264 146328 166316 146334
rect 166264 146270 166316 146276
rect 165528 95940 165580 95946
rect 165528 95882 165580 95888
rect 112350 94752 112406 94761
rect 112350 94687 112406 94696
rect 113178 94752 113234 94761
rect 113178 94687 113234 94696
rect 123206 94752 123262 94761
rect 123206 94687 123262 94696
rect 151910 94752 151966 94761
rect 151910 94687 151966 94696
rect 112364 93974 112392 94687
rect 112352 93968 112404 93974
rect 112352 93910 112404 93916
rect 113192 93906 113220 94687
rect 123220 94042 123248 94687
rect 126888 94512 126940 94518
rect 125598 94480 125654 94489
rect 126888 94454 126940 94460
rect 125598 94415 125654 94424
rect 123208 94036 123260 94042
rect 123208 93978 123260 93984
rect 113180 93900 113232 93906
rect 113180 93842 113232 93848
rect 121734 93664 121790 93673
rect 121734 93599 121790 93608
rect 93950 93528 94006 93537
rect 93950 93463 94006 93472
rect 107750 93528 107806 93537
rect 107750 93463 107806 93472
rect 93964 93226 93992 93463
rect 93952 93220 94004 93226
rect 93952 93162 94004 93168
rect 107764 93158 107792 93463
rect 121748 93362 121776 93599
rect 121736 93356 121788 93362
rect 121736 93298 121788 93304
rect 110142 93256 110198 93265
rect 110142 93191 110198 93200
rect 107752 93152 107804 93158
rect 107752 93094 107804 93100
rect 88984 92472 89036 92478
rect 85762 92440 85818 92449
rect 85762 92375 85818 92384
rect 87234 92440 87290 92449
rect 87234 92375 87290 92384
rect 88982 92440 88984 92449
rect 89036 92440 89038 92449
rect 88982 92375 89038 92384
rect 100482 92440 100538 92449
rect 100482 92375 100538 92384
rect 107474 92440 107530 92449
rect 107474 92375 107530 92384
rect 109682 92440 109738 92449
rect 109682 92375 109738 92384
rect 75826 91216 75882 91225
rect 75826 91151 75882 91160
rect 85486 91216 85542 91225
rect 85486 91151 85542 91160
rect 67732 86964 67784 86970
rect 67732 86906 67784 86912
rect 67272 82816 67324 82822
rect 67272 82758 67324 82764
rect 66904 77240 66956 77246
rect 66904 77182 66956 77188
rect 75840 77178 75868 91151
rect 75828 77172 75880 77178
rect 75828 77114 75880 77120
rect 49700 75200 49752 75206
rect 49700 75142 49752 75148
rect 49608 48272 49660 48278
rect 49608 48214 49660 48220
rect 49620 47938 49648 48214
rect 48964 47932 49016 47938
rect 48964 47874 49016 47880
rect 49608 47932 49660 47938
rect 49608 47874 49660 47880
rect 48320 32428 48372 32434
rect 48320 32370 48372 32376
rect 48332 16574 48360 32370
rect 45572 16546 46704 16574
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 45100 3528 45152 3534
rect 45100 3470 45152 3476
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45112 354 45140 3470
rect 46676 480 46704 16546
rect 45438 354 45550 480
rect 45112 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 48976 8974 49004 47874
rect 49712 16574 49740 75142
rect 52460 73908 52512 73914
rect 52460 73850 52512 73856
rect 51080 61396 51132 61402
rect 51080 61338 51132 61344
rect 49712 16546 50200 16574
rect 48964 8968 49016 8974
rect 48964 8910 49016 8916
rect 50172 480 50200 16546
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51092 354 51120 61338
rect 52472 6914 52500 73850
rect 85500 73166 85528 91151
rect 85776 91118 85804 92375
rect 87248 92342 87276 92375
rect 87236 92336 87288 92342
rect 87236 92278 87288 92284
rect 99286 91488 99342 91497
rect 99286 91423 99342 91432
rect 99102 91352 99158 91361
rect 99102 91287 99158 91296
rect 86866 91216 86922 91225
rect 86866 91151 86922 91160
rect 90730 91216 90786 91225
rect 90730 91151 90786 91160
rect 92386 91216 92442 91225
rect 92386 91151 92442 91160
rect 93766 91216 93822 91225
rect 93766 91151 93822 91160
rect 95146 91216 95202 91225
rect 95146 91151 95202 91160
rect 96526 91216 96582 91225
rect 96526 91151 96582 91160
rect 97078 91216 97134 91225
rect 97078 91151 97134 91160
rect 97906 91216 97962 91225
rect 97906 91151 97962 91160
rect 85764 91112 85816 91118
rect 85764 91054 85816 91060
rect 86880 79830 86908 91151
rect 90744 88262 90772 91151
rect 90732 88256 90784 88262
rect 90732 88198 90784 88204
rect 92400 81326 92428 91151
rect 92388 81320 92440 81326
rect 92388 81262 92440 81268
rect 86868 79824 86920 79830
rect 86868 79766 86920 79772
rect 93780 78402 93808 91151
rect 95160 80034 95188 91151
rect 96540 84046 96568 91151
rect 97092 86873 97120 91151
rect 97078 86864 97134 86873
rect 97078 86799 97134 86808
rect 96528 84040 96580 84046
rect 96528 83982 96580 83988
rect 97920 82754 97948 91151
rect 99116 84182 99144 91287
rect 99194 91216 99250 91225
rect 99194 91151 99250 91160
rect 99104 84176 99156 84182
rect 99104 84118 99156 84124
rect 97908 82748 97960 82754
rect 97908 82690 97960 82696
rect 95148 80028 95200 80034
rect 95148 79970 95200 79976
rect 99208 79762 99236 91151
rect 99196 79756 99248 79762
rect 99196 79698 99248 79704
rect 99300 78538 99328 91423
rect 100496 90914 100524 92375
rect 107488 92274 107516 92375
rect 107476 92268 107528 92274
rect 107476 92210 107528 92216
rect 104254 91624 104310 91633
rect 104254 91559 104310 91568
rect 101862 91488 101918 91497
rect 101862 91423 101918 91432
rect 100574 91216 100630 91225
rect 100574 91151 100630 91160
rect 100484 90908 100536 90914
rect 100484 90850 100536 90856
rect 99288 78532 99340 78538
rect 99288 78474 99340 78480
rect 93768 78396 93820 78402
rect 93768 78338 93820 78344
rect 100588 75886 100616 91151
rect 101876 85474 101904 91423
rect 102046 91352 102102 91361
rect 102046 91287 102102 91296
rect 103334 91352 103390 91361
rect 103334 91287 103390 91296
rect 101954 91216 102010 91225
rect 101954 91151 102010 91160
rect 101864 85468 101916 85474
rect 101864 85410 101916 85416
rect 101968 82793 101996 91151
rect 101954 82784 102010 82793
rect 101954 82719 102010 82728
rect 102060 78606 102088 91287
rect 103348 82618 103376 91287
rect 103426 91216 103482 91225
rect 103426 91151 103482 91160
rect 103336 82612 103388 82618
rect 103336 82554 103388 82560
rect 103440 81433 103468 91151
rect 104268 89486 104296 91559
rect 106186 91352 106242 91361
rect 106186 91287 106242 91296
rect 104806 91216 104862 91225
rect 104806 91151 104862 91160
rect 106094 91216 106150 91225
rect 106094 91151 106150 91160
rect 104256 89480 104308 89486
rect 104256 89422 104308 89428
rect 103426 81424 103482 81433
rect 103426 81359 103482 81368
rect 102048 78600 102100 78606
rect 102048 78542 102100 78548
rect 100576 75880 100628 75886
rect 100576 75822 100628 75828
rect 104820 74458 104848 91151
rect 106108 84153 106136 91151
rect 106094 84144 106150 84153
rect 106094 84079 106150 84088
rect 106200 77110 106228 91287
rect 107566 91216 107622 91225
rect 107566 91151 107622 91160
rect 108486 91216 108542 91225
rect 109696 91186 109724 92375
rect 108486 91151 108542 91160
rect 109684 91180 109736 91186
rect 107580 84114 107608 91151
rect 108500 85406 108528 91151
rect 109684 91122 109736 91128
rect 110156 86834 110184 93191
rect 111614 92440 111670 92449
rect 111614 92375 111670 92384
rect 114190 92440 114246 92449
rect 114190 92375 114246 92384
rect 118054 92440 118110 92449
rect 118054 92375 118056 92384
rect 110234 91216 110290 91225
rect 110234 91151 110290 91160
rect 110248 88233 110276 91151
rect 111628 90982 111656 92375
rect 114204 92206 114232 92375
rect 118108 92375 118110 92384
rect 124494 92440 124550 92449
rect 124494 92375 124550 92384
rect 125414 92440 125470 92449
rect 125414 92375 125470 92384
rect 118056 92346 118108 92352
rect 114192 92200 114244 92206
rect 114192 92142 114244 92148
rect 115386 91760 115442 91769
rect 115386 91695 115442 91704
rect 111706 91216 111762 91225
rect 111706 91151 111762 91160
rect 113086 91216 113142 91225
rect 113086 91151 113142 91160
rect 113914 91216 113970 91225
rect 113914 91151 113970 91160
rect 111616 90976 111668 90982
rect 111616 90918 111668 90924
rect 110234 88224 110290 88233
rect 110234 88159 110290 88168
rect 110144 86828 110196 86834
rect 110144 86770 110196 86776
rect 108488 85400 108540 85406
rect 108488 85342 108540 85348
rect 107568 84108 107620 84114
rect 107568 84050 107620 84056
rect 111720 82686 111748 91151
rect 111708 82680 111760 82686
rect 111708 82622 111760 82628
rect 106188 77104 106240 77110
rect 106188 77046 106240 77052
rect 113100 75818 113128 91151
rect 113928 85542 113956 91151
rect 115400 89622 115428 91695
rect 124126 91488 124182 91497
rect 124126 91423 124182 91432
rect 119894 91352 119950 91361
rect 119894 91287 119950 91296
rect 120722 91352 120778 91361
rect 120722 91287 120778 91296
rect 115846 91216 115902 91225
rect 117134 91216 117190 91225
rect 115846 91151 115902 91160
rect 116676 91180 116728 91186
rect 115388 89616 115440 89622
rect 115388 89558 115440 89564
rect 113916 85536 113968 85542
rect 113916 85478 113968 85484
rect 115860 83978 115888 91151
rect 117134 91151 117190 91160
rect 118238 91216 118294 91225
rect 118238 91151 118294 91160
rect 116676 91122 116728 91128
rect 116584 91112 116636 91118
rect 116584 91054 116636 91060
rect 115848 83972 115900 83978
rect 115848 83914 115900 83920
rect 113088 75812 113140 75818
rect 113088 75754 113140 75760
rect 116596 74526 116624 91054
rect 116688 78674 116716 91122
rect 117148 88194 117176 91151
rect 117136 88188 117188 88194
rect 117136 88130 117188 88136
rect 118252 86766 118280 91151
rect 118240 86760 118292 86766
rect 118240 86702 118292 86708
rect 119908 85338 119936 91287
rect 119986 91216 120042 91225
rect 119986 91151 120042 91160
rect 119896 85332 119948 85338
rect 119896 85274 119948 85280
rect 120000 79898 120028 91151
rect 120736 88058 120764 91287
rect 121366 91216 121422 91225
rect 121366 91151 121422 91160
rect 122746 91216 122802 91225
rect 122746 91151 122802 91160
rect 124034 91216 124090 91225
rect 124034 91151 124090 91160
rect 120724 88052 120776 88058
rect 120724 87994 120776 88000
rect 121380 79966 121408 91151
rect 121368 79960 121420 79966
rect 121368 79902 121420 79908
rect 119988 79892 120040 79898
rect 119988 79834 120040 79840
rect 116676 78668 116728 78674
rect 116676 78610 116728 78616
rect 122760 78470 122788 91151
rect 124048 85270 124076 91151
rect 124036 85264 124088 85270
rect 124036 85206 124088 85212
rect 124140 83910 124168 91423
rect 124508 90846 124536 92375
rect 124496 90840 124548 90846
rect 124496 90782 124548 90788
rect 125428 90778 125456 92375
rect 125416 90772 125468 90778
rect 125416 90714 125468 90720
rect 124128 83904 124180 83910
rect 124128 83846 124180 83852
rect 122748 78464 122800 78470
rect 122748 78406 122800 78412
rect 120080 76560 120132 76566
rect 120080 76502 120132 76508
rect 116584 74520 116636 74526
rect 116584 74462 116636 74468
rect 104808 74452 104860 74458
rect 104808 74394 104860 74400
rect 85488 73160 85540 73166
rect 85488 73102 85540 73108
rect 114560 72548 114612 72554
rect 114560 72490 114612 72496
rect 66260 72480 66312 72486
rect 66260 72422 66312 72428
rect 62120 68332 62172 68338
rect 62120 68274 62172 68280
rect 60740 64184 60792 64190
rect 60740 64126 60792 64132
rect 53840 60036 53892 60042
rect 53840 59978 53892 59984
rect 52552 54528 52604 54534
rect 52552 54470 52604 54476
rect 52564 16574 52592 54470
rect 53852 16574 53880 59978
rect 57980 57248 58032 57254
rect 57980 57190 58032 57196
rect 55218 36544 55274 36553
rect 55218 36479 55274 36488
rect 55232 16574 55260 36479
rect 56600 24200 56652 24206
rect 56600 24142 56652 24148
rect 56612 16574 56640 24142
rect 57992 16574 58020 57190
rect 60752 16574 60780 64126
rect 62132 16574 62160 68274
rect 63500 62892 63552 62898
rect 63500 62834 63552 62840
rect 63512 16574 63540 62834
rect 64880 55888 64932 55894
rect 64880 55830 64932 55836
rect 64892 16574 64920 55830
rect 66272 16574 66300 72422
rect 103520 71120 103572 71126
rect 103520 71062 103572 71068
rect 89720 69692 89772 69698
rect 89720 69634 89772 69640
rect 80060 65612 80112 65618
rect 80060 65554 80112 65560
rect 70400 61464 70452 61470
rect 70400 61406 70452 61412
rect 67638 59936 67694 59945
rect 67638 59871 67694 59880
rect 52564 16546 53328 16574
rect 53852 16546 54984 16574
rect 55232 16546 56088 16574
rect 56612 16546 56824 16574
rect 57992 16546 58480 16574
rect 60752 16546 60872 16574
rect 62132 16546 63264 16574
rect 63512 16546 64368 16574
rect 64892 16546 65104 16574
rect 66272 16546 66760 16574
rect 52472 6886 52592 6914
rect 52564 480 52592 6886
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53300 354 53328 16546
rect 54956 480 54984 16546
rect 56060 480 56088 16546
rect 53718 354 53830 480
rect 53300 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 58452 480 58480 16546
rect 59360 13116 59412 13122
rect 59360 13058 59412 13064
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 13058
rect 60844 480 60872 16546
rect 62028 8968 62080 8974
rect 62028 8910 62080 8916
rect 62040 480 62068 8910
rect 63236 480 63264 16546
rect 64340 480 64368 16546
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66732 480 66760 16546
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 59871
rect 69018 54496 69074 54505
rect 69018 54431 69074 54440
rect 69032 16574 69060 54431
rect 70412 16574 70440 61406
rect 74540 58676 74592 58682
rect 74540 58618 74592 58624
rect 71780 33856 71832 33862
rect 71780 33798 71832 33804
rect 71792 16574 71820 33798
rect 73160 31136 73212 31142
rect 73160 31078 73212 31084
rect 73172 16574 73200 31078
rect 74552 16574 74580 58618
rect 78680 44940 78732 44946
rect 78680 44882 78732 44888
rect 75920 42084 75972 42090
rect 75920 42026 75972 42032
rect 69032 16546 69152 16574
rect 70412 16546 71544 16574
rect 71792 16546 72648 16574
rect 73172 16546 73384 16574
rect 74552 16546 75040 16574
rect 69124 480 69152 16546
rect 70308 6180 70360 6186
rect 70308 6122 70360 6128
rect 70320 480 70348 6122
rect 71516 480 71544 16546
rect 72620 480 72648 16546
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 16546
rect 75012 480 75040 16546
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 75932 354 75960 42026
rect 77300 39364 77352 39370
rect 77300 39306 77352 39312
rect 77312 6914 77340 39306
rect 77390 17232 77446 17241
rect 77390 17167 77446 17176
rect 77404 16574 77432 17167
rect 78692 16574 78720 44882
rect 80072 16574 80100 65554
rect 81440 57316 81492 57322
rect 81440 57258 81492 57264
rect 81452 16574 81480 57258
rect 85580 55956 85632 55962
rect 85580 55898 85632 55904
rect 82820 49088 82872 49094
rect 82820 49030 82872 49036
rect 82832 16574 82860 49030
rect 77404 16546 78168 16574
rect 78692 16546 79272 16574
rect 80072 16546 80928 16574
rect 81452 16546 81664 16574
rect 82832 16546 83320 16574
rect 77312 6886 77432 6914
rect 77404 480 77432 6886
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78140 354 78168 16546
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 79244 354 79272 16546
rect 80900 480 80928 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83292 480 83320 16546
rect 84200 15904 84252 15910
rect 84200 15846 84252 15852
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 15846
rect 85592 6914 85620 55898
rect 85672 50448 85724 50454
rect 85672 50390 85724 50396
rect 85684 16574 85712 50390
rect 88340 46232 88392 46238
rect 88340 46174 88392 46180
rect 86960 22840 87012 22846
rect 86960 22782 87012 22788
rect 86972 16574 87000 22782
rect 88352 16574 88380 46174
rect 89732 16574 89760 69634
rect 93860 68400 93912 68406
rect 93860 68342 93912 68348
rect 91100 25628 91152 25634
rect 91100 25570 91152 25576
rect 91112 16574 91140 25570
rect 85684 16546 86448 16574
rect 86972 16546 87552 16574
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 91112 16546 91600 16574
rect 85592 6886 85712 6914
rect 85684 480 85712 6886
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86420 354 86448 16546
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 87524 354 87552 16546
rect 89180 480 89208 16546
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 92480 10328 92532 10334
rect 92480 10270 92532 10276
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 10270
rect 93872 6914 93900 68342
rect 96620 66904 96672 66910
rect 96620 66846 96672 66852
rect 93952 38004 94004 38010
rect 93952 37946 94004 37952
rect 93964 16574 93992 37946
rect 96632 16574 96660 66846
rect 98000 33788 98052 33794
rect 98000 33730 98052 33736
rect 98012 16574 98040 33730
rect 102140 28348 102192 28354
rect 102140 28290 102192 28296
rect 100760 26920 100812 26926
rect 100760 26862 100812 26868
rect 93964 16546 94728 16574
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 93872 6886 93992 6914
rect 93964 480 93992 6886
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94700 354 94728 16546
rect 96252 9036 96304 9042
rect 96252 8978 96304 8984
rect 96264 480 96292 8978
rect 97460 480 97488 16546
rect 95118 354 95230 480
rect 94700 326 95230 354
rect 95118 -960 95230 326
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99840 7676 99892 7682
rect 99840 7618 99892 7624
rect 99852 480 99880 7618
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 26862
rect 102152 16574 102180 28290
rect 103532 16574 103560 71062
rect 110420 51808 110472 51814
rect 110420 51750 110472 51756
rect 104900 42152 104952 42158
rect 104900 42094 104952 42100
rect 104912 16574 104940 42094
rect 107660 39432 107712 39438
rect 107660 39374 107712 39380
rect 106280 32496 106332 32502
rect 106280 32438 106332 32444
rect 106292 16574 106320 32438
rect 107672 16574 107700 39374
rect 109040 18692 109092 18698
rect 109040 18634 109092 18640
rect 102152 16546 102272 16574
rect 103532 16546 104112 16574
rect 104912 16546 105768 16574
rect 106292 16546 106504 16574
rect 107672 16546 108160 16574
rect 102244 480 102272 16546
rect 103336 3528 103388 3534
rect 103336 3470 103388 3476
rect 103348 480 103376 3470
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105740 480 105768 16546
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108132 480 108160 16546
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109052 354 109080 18634
rect 110432 3602 110460 51750
rect 110512 17332 110564 17338
rect 110512 17274 110564 17280
rect 110420 3596 110472 3602
rect 110420 3538 110472 3544
rect 110524 480 110552 17274
rect 114572 16574 114600 72490
rect 118700 29708 118752 29714
rect 118700 29650 118752 29656
rect 117318 26888 117374 26897
rect 117318 26823 117374 26832
rect 115940 20052 115992 20058
rect 115940 19994 115992 20000
rect 115952 16574 115980 19994
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 112352 11824 112404 11830
rect 112352 11766 112404 11772
rect 111616 3596 111668 3602
rect 111616 3538 111668 3544
rect 111628 480 111656 3538
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 11766
rect 114008 3664 114060 3670
rect 114008 3606 114060 3612
rect 114020 480 114048 3606
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 26823
rect 118712 3602 118740 29650
rect 120092 16574 120120 76502
rect 124220 69760 124272 69766
rect 124220 69702 124272 69708
rect 121460 53168 121512 53174
rect 121460 53110 121512 53116
rect 121472 16574 121500 53110
rect 122840 40724 122892 40730
rect 122840 40666 122892 40672
rect 122852 16574 122880 40666
rect 124232 16574 124260 69702
rect 120092 16546 120672 16574
rect 121472 16546 122328 16574
rect 122852 16546 123064 16574
rect 124232 16546 124720 16574
rect 118700 3596 118752 3602
rect 118700 3538 118752 3544
rect 119896 3596 119948 3602
rect 119896 3538 119948 3544
rect 118792 2168 118844 2174
rect 118792 2110 118844 2116
rect 118804 480 118832 2110
rect 119908 480 119936 3538
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 122300 480 122328 16546
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 124692 480 124720 16546
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125612 354 125640 94415
rect 125782 92440 125838 92449
rect 125782 92375 125838 92384
rect 125796 92138 125824 92375
rect 126900 92342 126928 94454
rect 151924 94110 151952 94687
rect 151912 94104 151964 94110
rect 151912 94046 151964 94052
rect 151542 93528 151598 93537
rect 151542 93463 151598 93472
rect 151556 93294 151584 93463
rect 151544 93288 151596 93294
rect 128174 93256 128230 93265
rect 151544 93230 151596 93236
rect 128174 93191 128230 93200
rect 126888 92336 126940 92342
rect 126888 92278 126940 92284
rect 125784 92132 125836 92138
rect 125784 92074 125836 92080
rect 126886 91352 126942 91361
rect 126886 91287 126942 91296
rect 126794 91216 126850 91225
rect 126794 91151 126850 91160
rect 126808 81190 126836 91151
rect 126900 81258 126928 91287
rect 128188 89554 128216 93191
rect 128358 93120 128414 93129
rect 128358 93055 128414 93064
rect 128372 92274 128400 93055
rect 165540 92478 165568 95882
rect 165528 92472 165580 92478
rect 129462 92440 129518 92449
rect 129462 92375 129518 92384
rect 135718 92440 135774 92449
rect 165528 92414 165580 92420
rect 135718 92375 135774 92384
rect 129476 92342 129504 92375
rect 129464 92336 129516 92342
rect 129464 92278 129516 92284
rect 135732 92274 135760 92375
rect 128360 92268 128412 92274
rect 128360 92210 128412 92216
rect 135720 92268 135772 92274
rect 135720 92210 135772 92216
rect 151726 92168 151782 92177
rect 151726 92103 151782 92112
rect 132222 91624 132278 91633
rect 132222 91559 132278 91568
rect 151358 91624 151414 91633
rect 151358 91559 151414 91568
rect 130750 91216 130806 91225
rect 130750 91151 130806 91160
rect 128176 89548 128228 89554
rect 128176 89490 128228 89496
rect 130764 86698 130792 91151
rect 132236 89350 132264 91559
rect 133142 91216 133198 91225
rect 133142 91151 133198 91160
rect 134706 91216 134762 91225
rect 134706 91151 134762 91160
rect 132224 89344 132276 89350
rect 132224 89286 132276 89292
rect 133156 88126 133184 91151
rect 133144 88120 133196 88126
rect 133144 88062 133196 88068
rect 130752 86692 130804 86698
rect 130752 86634 130804 86640
rect 134720 85202 134748 91151
rect 151372 89418 151400 91559
rect 151740 90710 151768 92103
rect 151728 90704 151780 90710
rect 151728 90646 151780 90652
rect 151360 89412 151412 89418
rect 151360 89354 151412 89360
rect 166276 85202 166304 146270
rect 167644 144968 167696 144974
rect 167644 144910 167696 144916
rect 166356 124228 166408 124234
rect 166356 124170 166408 124176
rect 166368 85270 166396 124170
rect 166448 118720 166500 118726
rect 166448 118662 166500 118668
rect 166460 93974 166488 118662
rect 166540 100020 166592 100026
rect 166540 99962 166592 99968
rect 166448 93968 166500 93974
rect 166448 93910 166500 93916
rect 166552 92138 166580 99962
rect 166540 92132 166592 92138
rect 166540 92074 166592 92080
rect 167000 91860 167052 91866
rect 167000 91802 167052 91808
rect 167012 89350 167040 91802
rect 167000 89344 167052 89350
rect 167000 89286 167052 89292
rect 167656 86698 167684 144910
rect 167828 140072 167880 140078
rect 167828 140014 167880 140020
rect 167736 122868 167788 122874
rect 167736 122810 167788 122816
rect 167748 93362 167776 122810
rect 167840 110129 167868 140014
rect 170404 135380 170456 135386
rect 170404 135322 170456 135328
rect 169116 135312 169168 135318
rect 169116 135254 169168 135260
rect 169024 128376 169076 128382
rect 169024 128318 169076 128324
rect 167920 122120 167972 122126
rect 167920 122062 167972 122068
rect 167932 111761 167960 122062
rect 167918 111752 167974 111761
rect 167918 111687 167974 111696
rect 167826 110120 167882 110129
rect 167826 110055 167882 110064
rect 167920 109064 167972 109070
rect 167920 109006 167972 109012
rect 167828 98048 167880 98054
rect 167828 97990 167880 97996
rect 167736 93356 167788 93362
rect 167736 93298 167788 93304
rect 167644 86692 167696 86698
rect 167644 86634 167696 86640
rect 166356 85264 166408 85270
rect 166356 85206 166408 85212
rect 134708 85196 134760 85202
rect 134708 85138 134760 85144
rect 166264 85196 166316 85202
rect 166264 85138 166316 85144
rect 126888 81252 126940 81258
rect 126888 81194 126940 81200
rect 126796 81184 126848 81190
rect 126796 81126 126848 81132
rect 167840 79830 167868 97990
rect 167932 84046 167960 109006
rect 168104 108996 168156 109002
rect 168104 108938 168156 108944
rect 168116 108769 168144 108938
rect 168102 108760 168158 108769
rect 168102 108695 168158 108704
rect 167920 84040 167972 84046
rect 167920 83982 167972 83988
rect 167828 79824 167880 79830
rect 167828 79766 167880 79772
rect 169036 79762 169064 128318
rect 169128 93906 169156 135254
rect 169208 110492 169260 110498
rect 169208 110434 169260 110440
rect 169116 93900 169168 93906
rect 169116 93842 169168 93848
rect 169220 90914 169248 110434
rect 169300 100088 169352 100094
rect 169300 100030 169352 100036
rect 169312 92206 169340 100030
rect 169300 92200 169352 92206
rect 169300 92142 169352 92148
rect 169208 90908 169260 90914
rect 169208 90850 169260 90856
rect 169024 79756 169076 79762
rect 169024 79698 169076 79704
rect 170416 75818 170444 135322
rect 170496 124296 170548 124302
rect 170496 124238 170548 124244
rect 170508 83910 170536 124238
rect 170588 122936 170640 122942
rect 170588 122878 170640 122884
rect 170600 88058 170628 122878
rect 170680 106344 170732 106350
rect 170680 106286 170732 106292
rect 170588 88052 170640 88058
rect 170588 87994 170640 88000
rect 170496 83904 170548 83910
rect 170496 83846 170548 83852
rect 170692 78402 170720 106286
rect 171796 94110 171824 151778
rect 171876 138032 171928 138038
rect 171876 137974 171928 137980
rect 171784 94104 171836 94110
rect 171784 94046 171836 94052
rect 171888 85338 171916 137974
rect 172348 127634 172376 160103
rect 172336 127628 172388 127634
rect 172336 127570 172388 127576
rect 171968 113212 172020 113218
rect 171968 113154 172020 113160
rect 171980 89486 172008 113154
rect 172440 99346 172468 359110
rect 173164 359100 173216 359106
rect 173164 359042 173216 359048
rect 173176 310486 173204 359042
rect 175108 333742 175136 367066
rect 178684 362976 178736 362982
rect 178684 362918 178736 362924
rect 176108 360528 176160 360534
rect 176108 360470 176160 360476
rect 176016 360460 176068 360466
rect 176016 360402 176068 360408
rect 175924 356312 175976 356318
rect 175924 356254 175976 356260
rect 175188 342304 175240 342310
rect 175188 342246 175240 342252
rect 175096 333736 175148 333742
rect 175096 333678 175148 333684
rect 175108 333266 175136 333678
rect 175096 333260 175148 333266
rect 175096 333202 175148 333208
rect 175096 327140 175148 327146
rect 175096 327082 175148 327088
rect 173164 310480 173216 310486
rect 173164 310422 173216 310428
rect 173808 305040 173860 305046
rect 173808 304982 173860 304988
rect 173164 294024 173216 294030
rect 173164 293966 173216 293972
rect 172428 99340 172480 99346
rect 172428 99282 172480 99288
rect 172060 95260 172112 95266
rect 172060 95202 172112 95208
rect 171968 89480 172020 89486
rect 171968 89422 172020 89428
rect 171876 85332 171928 85338
rect 171876 85274 171928 85280
rect 170680 78396 170732 78402
rect 170680 78338 170732 78344
rect 172072 77178 172100 95202
rect 173176 95169 173204 293966
rect 173256 244316 173308 244322
rect 173256 244258 173308 244264
rect 173268 231198 173296 244258
rect 173820 240650 173848 304982
rect 174636 251252 174688 251258
rect 174636 251194 174688 251200
rect 174544 248464 174596 248470
rect 174544 248406 174596 248412
rect 173808 240644 173860 240650
rect 173808 240586 173860 240592
rect 173256 231192 173308 231198
rect 173256 231134 173308 231140
rect 173348 140820 173400 140826
rect 173348 140762 173400 140768
rect 173256 132524 173308 132530
rect 173256 132466 173308 132472
rect 173162 95160 173218 95169
rect 173162 95095 173218 95104
rect 173268 85406 173296 132466
rect 173360 94042 173388 140762
rect 173440 125656 173492 125662
rect 173440 125598 173492 125604
rect 173348 94036 173400 94042
rect 173348 93978 173400 93984
rect 173452 90778 173480 125598
rect 174556 95198 174584 248406
rect 174648 235686 174676 251194
rect 174636 235680 174688 235686
rect 174636 235622 174688 235628
rect 174544 95192 174596 95198
rect 174544 95134 174596 95140
rect 173440 90772 173492 90778
rect 173440 90714 173492 90720
rect 173256 85400 173308 85406
rect 173256 85342 173308 85348
rect 172060 77172 172112 77178
rect 172060 77114 172112 77120
rect 170404 75812 170456 75818
rect 170404 75754 170456 75760
rect 175108 75274 175136 327082
rect 175096 75268 175148 75274
rect 175096 75210 175148 75216
rect 175200 15978 175228 342246
rect 175936 285666 175964 356254
rect 176028 351218 176056 360402
rect 176120 352578 176148 360470
rect 176658 354376 176714 354385
rect 176658 354311 176714 354320
rect 176672 354006 176700 354311
rect 176660 354000 176712 354006
rect 176660 353942 176712 353948
rect 176108 352572 176160 352578
rect 176108 352514 176160 352520
rect 176566 352200 176622 352209
rect 176566 352135 176622 352144
rect 176016 351212 176068 351218
rect 176016 351154 176068 351160
rect 176474 310040 176530 310049
rect 176474 309975 176530 309984
rect 176488 307086 176516 309975
rect 176476 307080 176528 307086
rect 176476 307022 176528 307028
rect 176382 292360 176438 292369
rect 176382 292295 176438 292304
rect 175924 285660 175976 285666
rect 175924 285602 175976 285608
rect 175280 280832 175332 280838
rect 175280 280774 175332 280780
rect 175292 276078 175320 280774
rect 175280 276072 175332 276078
rect 175280 276014 175332 276020
rect 175924 256760 175976 256766
rect 175924 256702 175976 256708
rect 175936 237182 175964 256702
rect 175924 237176 175976 237182
rect 175924 237118 175976 237124
rect 176396 84862 176424 292295
rect 176474 252920 176530 252929
rect 176474 252855 176530 252864
rect 176384 84856 176436 84862
rect 176384 84798 176436 84804
rect 175188 15972 175240 15978
rect 175188 15914 175240 15920
rect 135260 14544 135312 14550
rect 135260 14486 135312 14492
rect 128912 11892 128964 11898
rect 128912 11834 128964 11840
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 11834
rect 135272 3398 135300 14486
rect 176488 10402 176516 252855
rect 176580 29782 176608 352135
rect 176658 345400 176714 345409
rect 176658 345335 176714 345344
rect 176672 345098 176700 345335
rect 176660 345092 176712 345098
rect 176660 345034 176712 345040
rect 176842 343360 176898 343369
rect 176842 343295 176898 343304
rect 176856 342310 176884 343295
rect 176844 342304 176896 342310
rect 176844 342246 176896 342252
rect 176842 334520 176898 334529
rect 176842 334455 176898 334464
rect 176856 334014 176884 334455
rect 176844 334008 176896 334014
rect 176844 333950 176896 333956
rect 176660 333736 176712 333742
rect 176660 333678 176712 333684
rect 176672 332625 176700 333678
rect 176658 332616 176714 332625
rect 176658 332551 176714 332560
rect 176658 327720 176714 327729
rect 176658 327655 176714 327664
rect 176672 327146 176700 327655
rect 176660 327140 176712 327146
rect 176660 327082 176712 327088
rect 176658 325816 176714 325825
rect 176658 325751 176714 325760
rect 176672 325718 176700 325751
rect 176660 325712 176712 325718
rect 176660 325654 176712 325660
rect 177946 321600 178002 321609
rect 177946 321535 178002 321544
rect 177854 318880 177910 318889
rect 177854 318815 177910 318824
rect 176658 314800 176714 314809
rect 176658 314735 176714 314744
rect 176672 314702 176700 314735
rect 176660 314696 176712 314702
rect 176660 314638 176712 314644
rect 176658 312760 176714 312769
rect 176658 312695 176714 312704
rect 176672 312594 176700 312695
rect 176660 312588 176712 312594
rect 176660 312530 176712 312536
rect 176658 305960 176714 305969
rect 176658 305895 176714 305904
rect 176672 305046 176700 305895
rect 176660 305040 176712 305046
rect 176660 304982 176712 304988
rect 176658 301200 176714 301209
rect 176658 301135 176714 301144
rect 176672 300966 176700 301135
rect 176660 300960 176712 300966
rect 176660 300902 176712 300908
rect 176658 299160 176714 299169
rect 176658 299095 176714 299104
rect 176672 298110 176700 299095
rect 176660 298104 176712 298110
rect 176660 298046 176712 298052
rect 176660 297424 176712 297430
rect 176660 297366 176712 297372
rect 176672 297265 176700 297366
rect 176658 297256 176714 297265
rect 176658 297191 176714 297200
rect 176658 295080 176714 295089
rect 176658 295015 176714 295024
rect 176672 291854 176700 295015
rect 176660 291848 176712 291854
rect 176660 291790 176712 291796
rect 176658 290320 176714 290329
rect 176658 290255 176714 290264
rect 176672 289882 176700 290255
rect 176660 289876 176712 289882
rect 176660 289818 176712 289824
rect 176658 286240 176714 286249
rect 176658 286175 176714 286184
rect 176672 285734 176700 286175
rect 176660 285728 176712 285734
rect 176660 285670 176712 285676
rect 176658 283520 176714 283529
rect 176658 283455 176714 283464
rect 176672 282946 176700 283455
rect 176660 282940 176712 282946
rect 176660 282882 176712 282888
rect 176658 281616 176714 281625
rect 176658 281551 176660 281560
rect 176712 281551 176714 281560
rect 176660 281522 176712 281528
rect 176660 280152 176712 280158
rect 176660 280094 176712 280100
rect 176672 279585 176700 280094
rect 176658 279576 176714 279585
rect 176658 279511 176714 279520
rect 176660 278724 176712 278730
rect 176660 278666 176712 278672
rect 176672 277545 176700 278666
rect 176658 277536 176714 277545
rect 176658 277471 176714 277480
rect 177488 276004 177540 276010
rect 177488 275946 177540 275952
rect 177500 274825 177528 275946
rect 177486 274816 177542 274825
rect 177486 274751 177542 274760
rect 176658 272640 176714 272649
rect 176658 272575 176714 272584
rect 176672 271930 176700 272575
rect 176660 271924 176712 271930
rect 176660 271866 176712 271872
rect 177762 270600 177818 270609
rect 177762 270535 177818 270544
rect 176658 268560 176714 268569
rect 176658 268495 176714 268504
rect 176672 267782 176700 268495
rect 176660 267776 176712 267782
rect 176660 267718 176712 267724
rect 176660 266348 176712 266354
rect 176660 266290 176712 266296
rect 176672 265985 176700 266290
rect 176658 265976 176714 265985
rect 176658 265911 176714 265920
rect 176658 261760 176714 261769
rect 176658 261695 176714 261704
rect 176672 261526 176700 261695
rect 176660 261520 176712 261526
rect 176660 261462 176712 261468
rect 176658 259720 176714 259729
rect 176658 259655 176714 259664
rect 176672 259486 176700 259655
rect 176660 259480 176712 259486
rect 176660 259422 176712 259428
rect 176658 254960 176714 254969
rect 176658 254895 176714 254904
rect 176672 254046 176700 254895
rect 176660 254040 176712 254046
rect 176660 253982 176712 253988
rect 177670 250880 177726 250889
rect 177670 250815 177726 250824
rect 176658 246120 176714 246129
rect 176658 246055 176714 246064
rect 176672 245682 176700 246055
rect 176660 245676 176712 245682
rect 176660 245618 176712 245624
rect 177578 242040 177634 242049
rect 177578 241975 177634 241984
rect 177592 241534 177620 241975
rect 177580 241528 177632 241534
rect 177580 241470 177632 241476
rect 177684 227322 177712 250815
rect 177672 227316 177724 227322
rect 177672 227258 177724 227264
rect 177776 160750 177804 270535
rect 177764 160744 177816 160750
rect 177764 160686 177816 160692
rect 177304 153264 177356 153270
rect 177304 153206 177356 153212
rect 177316 90710 177344 153206
rect 177868 148374 177896 318815
rect 177856 148368 177908 148374
rect 177856 148310 177908 148316
rect 177488 137284 177540 137290
rect 177488 137226 177540 137232
rect 177396 114572 177448 114578
rect 177396 114514 177448 114520
rect 177304 90704 177356 90710
rect 177304 90646 177356 90652
rect 177408 77110 177436 114514
rect 177500 109002 177528 137226
rect 177488 108996 177540 109002
rect 177488 108938 177540 108944
rect 177396 77104 177448 77110
rect 177396 77046 177448 77052
rect 177960 35358 177988 321535
rect 178696 302258 178724 362918
rect 178684 302252 178736 302258
rect 178684 302194 178736 302200
rect 178696 288425 178724 302194
rect 178682 288416 178738 288425
rect 178682 288351 178738 288360
rect 179064 257378 179092 697546
rect 189080 365832 189132 365838
rect 189080 365774 189132 365780
rect 189092 364334 189120 365774
rect 189092 364306 189304 364334
rect 181628 361820 181680 361826
rect 181628 361762 181680 361768
rect 179512 361684 179564 361690
rect 179512 361626 179564 361632
rect 179236 358828 179288 358834
rect 179236 358770 179288 358776
rect 179248 345014 179276 358770
rect 179524 348197 179552 361626
rect 179786 357776 179842 357785
rect 179786 357711 179842 357720
rect 179800 354074 179828 357711
rect 179880 357672 179932 357678
rect 179880 357614 179932 357620
rect 179788 354068 179840 354074
rect 179788 354010 179840 354016
rect 179892 351286 179920 357614
rect 181640 355042 181668 361762
rect 182916 357808 182968 357814
rect 182916 357750 182968 357756
rect 181332 355014 181668 355042
rect 182928 355042 182956 357750
rect 186780 357740 186832 357746
rect 186780 357682 186832 357688
rect 184940 357604 184992 357610
rect 184940 357546 184992 357552
rect 184952 355042 184980 357546
rect 186792 355042 186820 357682
rect 189276 355042 189304 364306
rect 193232 361962 193260 700266
rect 195244 374672 195296 374678
rect 195244 374614 195296 374620
rect 193220 361956 193272 361962
rect 193220 361898 193272 361904
rect 193232 357649 193260 361898
rect 195256 361622 195284 374614
rect 198740 369912 198792 369918
rect 198740 369854 198792 369860
rect 198752 364334 198780 369854
rect 201512 366450 201540 702986
rect 206284 702500 206336 702506
rect 206284 702442 206336 702448
rect 202880 368688 202932 368694
rect 202880 368630 202932 368636
rect 201500 366444 201552 366450
rect 201500 366386 201552 366392
rect 202892 364334 202920 368630
rect 198752 364306 199608 364334
rect 202892 364306 203472 364334
rect 195244 361616 195296 361622
rect 195244 361558 195296 361564
rect 195256 357746 195284 361558
rect 195244 357740 195296 357746
rect 195244 357682 195296 357688
rect 193218 357640 193274 357649
rect 191748 357604 191800 357610
rect 193218 357575 193274 357584
rect 193862 357640 193918 357649
rect 193862 357575 193918 357584
rect 191748 357546 191800 357552
rect 191760 355042 191788 357546
rect 193876 355042 193904 357575
rect 182928 355014 183264 355042
rect 184952 355014 185196 355042
rect 186792 355014 187128 355042
rect 189276 355014 189704 355042
rect 191636 355014 191788 355042
rect 193568 355014 193904 355042
rect 195256 355042 195284 357682
rect 197728 356380 197780 356386
rect 197728 356322 197780 356328
rect 197740 355042 197768 356322
rect 199580 355042 199608 364306
rect 201592 359032 201644 359038
rect 201592 358974 201644 358980
rect 200028 357740 200080 357746
rect 200028 357682 200080 357688
rect 200040 357406 200068 357682
rect 200028 357400 200080 357406
rect 200028 357342 200080 357348
rect 201500 357400 201552 357406
rect 201500 357342 201552 357348
rect 201512 355337 201540 357342
rect 201498 355328 201554 355337
rect 201498 355263 201554 355272
rect 201604 355042 201632 358974
rect 203444 355042 203472 364306
rect 206296 357513 206324 702442
rect 218992 700398 219020 703520
rect 218980 700392 219032 700398
rect 218980 700334 219032 700340
rect 235184 700330 235212 703520
rect 235172 700324 235224 700330
rect 235172 700266 235224 700272
rect 267660 697610 267688 703520
rect 283852 702434 283880 703520
rect 282932 702406 283880 702434
rect 267648 697604 267700 697610
rect 267648 697546 267700 697552
rect 212448 696244 212500 696250
rect 212448 696186 212500 696192
rect 209044 376780 209096 376786
rect 209044 376722 209096 376728
rect 209056 365702 209084 376722
rect 212460 369918 212488 696186
rect 274548 470620 274600 470626
rect 274548 470562 274600 470568
rect 247040 381540 247092 381546
rect 247040 381482 247092 381488
rect 232504 371340 232556 371346
rect 232504 371282 232556 371288
rect 211804 369912 211856 369918
rect 211804 369854 211856 369860
rect 212448 369912 212500 369918
rect 212448 369854 212500 369860
rect 208400 365696 208452 365702
rect 208400 365638 208452 365644
rect 209044 365696 209096 365702
rect 209044 365638 209096 365644
rect 208412 364546 208440 365638
rect 208400 364540 208452 364546
rect 208400 364482 208452 364488
rect 206282 357504 206338 357513
rect 206282 357439 206338 357448
rect 206296 355042 206324 357439
rect 208412 355314 208440 364482
rect 211816 357785 211844 369854
rect 226340 367328 226392 367334
rect 226340 367270 226392 367276
rect 219440 365764 219492 365770
rect 219440 365706 219492 365712
rect 213918 364440 213974 364449
rect 213918 364375 213974 364384
rect 213932 358766 213960 364375
rect 219452 360466 219480 365706
rect 226352 364334 226380 367270
rect 226352 364306 226656 364334
rect 219440 360460 219492 360466
rect 219440 360402 219492 360408
rect 220268 360460 220320 360466
rect 220268 360402 220320 360408
rect 218336 359168 218388 359174
rect 218336 359110 218388 359116
rect 213920 358760 213972 358766
rect 213920 358702 213972 358708
rect 214472 358760 214524 358766
rect 214472 358702 214524 358708
rect 211802 357776 211858 357785
rect 211802 357711 211858 357720
rect 208366 355286 208440 355314
rect 195256 355014 195500 355042
rect 197740 355014 198076 355042
rect 199580 355014 200008 355042
rect 201604 355014 201940 355042
rect 203444 355014 203872 355042
rect 206296 355014 206448 355042
rect 208366 355028 208394 355286
rect 211816 355042 211844 357711
rect 214484 357678 214512 358702
rect 217048 358148 217100 358154
rect 217048 358090 217100 358096
rect 214564 358080 214616 358086
rect 214564 358022 214616 358028
rect 214472 357672 214524 357678
rect 214472 357614 214524 357620
rect 214484 355042 214512 357614
rect 214576 356726 214604 358022
rect 214564 356720 214616 356726
rect 214564 356662 214616 356668
rect 217060 355042 217088 358090
rect 211816 355014 212244 355042
rect 214484 355014 214820 355042
rect 216752 355014 217088 355042
rect 218348 355042 218376 359110
rect 220280 355042 220308 360402
rect 223488 357672 223540 357678
rect 223488 357614 223540 357620
rect 223500 355042 223528 357614
rect 225420 356380 225472 356386
rect 225420 356322 225472 356328
rect 225432 355042 225460 356322
rect 218348 355014 218684 355042
rect 220280 355014 220616 355042
rect 223192 355014 223528 355042
rect 225124 355014 225460 355042
rect 226628 355042 226656 364306
rect 228824 363180 228876 363186
rect 228824 363122 228876 363128
rect 226628 355014 227056 355042
rect 209962 354920 210018 354929
rect 210018 354878 210312 354906
rect 209962 354855 210018 354864
rect 228836 354770 228864 363122
rect 231676 361888 231728 361894
rect 231676 361830 231728 361836
rect 231688 354770 231716 361830
rect 232516 358154 232544 371282
rect 234620 366376 234672 366382
rect 234620 366318 234672 366324
rect 233792 360460 233844 360466
rect 233792 360402 233844 360408
rect 232504 358148 232556 358154
rect 232504 358090 232556 358096
rect 233804 355042 233832 360402
rect 234632 359038 234660 366318
rect 238760 364608 238812 364614
rect 238760 364550 238812 364556
rect 238772 364334 238800 364550
rect 238772 364306 239536 364334
rect 237472 360528 237524 360534
rect 237472 360470 237524 360476
rect 234620 359032 234672 359038
rect 234620 358974 234672 358980
rect 235540 359032 235592 359038
rect 235540 358974 235592 358980
rect 233496 355014 233832 355042
rect 235080 355020 235132 355026
rect 235080 354962 235132 354968
rect 235092 354906 235120 354962
rect 235552 354906 235580 358974
rect 237484 354906 237512 360470
rect 239508 355042 239536 364306
rect 243634 363080 243690 363089
rect 243634 363015 243690 363024
rect 243648 361622 243676 363015
rect 243636 361616 243688 361622
rect 243636 361558 243688 361564
rect 242162 357504 242218 357513
rect 242162 357439 242218 357448
rect 242176 355042 242204 357439
rect 239508 355014 239936 355042
rect 241716 355014 242204 355042
rect 243648 355042 243676 361558
rect 245844 360256 245896 360262
rect 245844 360198 245896 360204
rect 243648 355014 243800 355042
rect 235092 354878 235580 354906
rect 237360 354878 237512 354906
rect 228836 354742 228988 354770
rect 231564 354742 231716 354770
rect 241716 354754 241744 355014
rect 245856 354770 245884 360198
rect 247052 354793 247080 381482
rect 270500 380180 270552 380186
rect 270500 380122 270552 380128
rect 267004 371272 267056 371278
rect 267004 371214 267056 371220
rect 264244 367192 264296 367198
rect 264244 367134 264296 367140
rect 251180 364540 251232 364546
rect 251180 364482 251232 364488
rect 251192 364334 251220 364482
rect 251192 364306 251772 364334
rect 250536 360596 250588 360602
rect 250536 360538 250588 360544
rect 250548 355042 250576 360538
rect 250240 355014 250576 355042
rect 251744 355042 251772 364306
rect 264256 358970 264284 367134
rect 253940 358964 253992 358970
rect 253940 358906 253992 358912
rect 264244 358964 264296 358970
rect 264244 358906 264296 358912
rect 264888 358964 264940 358970
rect 264888 358906 264940 358912
rect 253952 356454 253980 358906
rect 258906 358864 258962 358873
rect 258906 358799 258962 358808
rect 256792 357536 256844 357542
rect 256792 357478 256844 357484
rect 253940 356448 253992 356454
rect 253940 356390 253992 356396
rect 253952 355042 253980 356390
rect 251744 355014 252172 355042
rect 253952 355014 254104 355042
rect 256804 354929 256832 357478
rect 258920 355042 258948 358799
rect 264900 357490 264928 358906
rect 267016 357746 267044 371214
rect 269026 357776 269082 357785
rect 267004 357740 267056 357746
rect 269026 357711 269082 357720
rect 267004 357682 267056 357688
rect 264900 357462 265020 357490
rect 262772 356108 262824 356114
rect 262772 356050 262824 356056
rect 258612 355014 258948 355042
rect 256790 354920 256846 354929
rect 262784 354906 262812 356050
rect 264992 355314 265020 357462
rect 267016 355314 267044 357682
rect 264992 355286 265066 355314
rect 265038 355028 265066 355286
rect 266970 355286 267044 355314
rect 266970 355028 266998 355286
rect 269040 355042 269068 357711
rect 270512 356250 270540 380122
rect 274560 356794 274588 470562
rect 282932 368626 282960 702406
rect 300136 700466 300164 703520
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 300124 700460 300176 700466
rect 300124 700402 300176 700408
rect 310520 700460 310572 700466
rect 310520 700402 310572 700408
rect 309140 700392 309192 700398
rect 309140 700334 309192 700340
rect 299480 700324 299532 700330
rect 299480 700266 299532 700272
rect 302056 700324 302108 700330
rect 302056 700266 302108 700272
rect 295340 378820 295392 378826
rect 295340 378762 295392 378768
rect 291844 372632 291896 372638
rect 291844 372574 291896 372580
rect 282920 368620 282972 368626
rect 282920 368562 282972 368568
rect 282932 367810 282960 368562
rect 282920 367804 282972 367810
rect 282920 367746 282972 367752
rect 282920 364472 282972 364478
rect 282920 364414 282972 364420
rect 279332 360664 279384 360670
rect 279332 360606 279384 360612
rect 280068 360664 280120 360670
rect 280068 360606 280120 360612
rect 275008 360324 275060 360330
rect 275008 360266 275060 360272
rect 275020 358086 275048 360266
rect 275008 358080 275060 358086
rect 275008 358022 275060 358028
rect 276940 358080 276992 358086
rect 276940 358022 276992 358028
rect 275652 357808 275704 357814
rect 275652 357750 275704 357756
rect 273536 356788 273588 356794
rect 273536 356730 273588 356736
rect 274548 356788 274600 356794
rect 274548 356730 274600 356736
rect 273548 356318 273576 356730
rect 273536 356312 273588 356318
rect 273536 356254 273588 356260
rect 270500 356244 270552 356250
rect 270500 356186 270552 356192
rect 268916 355014 269068 355042
rect 270512 355042 270540 356186
rect 270512 355014 270848 355042
rect 273548 354906 273576 356254
rect 274560 356153 274588 356730
rect 274546 356144 274602 356153
rect 274546 356079 274602 356088
rect 275664 355042 275692 357750
rect 275356 355014 275692 355042
rect 276952 355042 276980 358022
rect 276952 355014 277288 355042
rect 262476 354878 262812 354906
rect 273424 354878 273576 354906
rect 256790 354855 256846 354864
rect 241704 354748 241756 354754
rect 245732 354742 245884 354770
rect 247038 354784 247094 354793
rect 247038 354719 247094 354728
rect 248142 354784 248198 354793
rect 256804 354770 256832 354855
rect 279344 354770 279372 360606
rect 280080 360262 280108 360606
rect 280068 360256 280120 360262
rect 280068 360198 280120 360204
rect 282932 358766 282960 364414
rect 287428 363112 287480 363118
rect 287428 363054 287480 363060
rect 282920 358760 282972 358766
rect 282920 358702 282972 358708
rect 283564 358760 283616 358766
rect 283564 358702 283616 358708
rect 283576 357542 283604 358702
rect 287440 357610 287468 363054
rect 285680 357604 285732 357610
rect 285680 357546 285732 357552
rect 287428 357604 287480 357610
rect 287428 357546 287480 357552
rect 283564 357536 283616 357542
rect 283564 357478 283616 357484
rect 282090 356280 282146 356289
rect 282090 356215 282146 356224
rect 282104 355042 282132 356215
rect 281796 355014 282132 355042
rect 283576 354906 283604 357478
rect 285692 356726 285720 357546
rect 285680 356720 285732 356726
rect 285680 356662 285732 356668
rect 287440 354906 287468 357546
rect 283576 354878 283728 354906
rect 287440 354878 287592 354906
rect 290168 354890 290504 354906
rect 290168 354884 290516 354890
rect 290168 354878 290464 354884
rect 290464 354826 290516 354832
rect 285956 354816 286008 354822
rect 248198 354742 248308 354770
rect 256680 354742 256832 354770
rect 260544 354754 260788 354770
rect 260544 354748 260800 354754
rect 260544 354742 260748 354748
rect 248142 354719 248198 354728
rect 241704 354690 241756 354696
rect 279220 354742 279372 354770
rect 285660 354764 285956 354770
rect 285660 354758 286008 354764
rect 285660 354742 285996 354758
rect 260748 354690 260800 354696
rect 291856 354674 291884 372574
rect 293960 367804 294012 367810
rect 293960 367746 294012 367752
rect 293132 358896 293184 358902
rect 293132 358838 293184 358844
rect 292132 357734 292344 357762
rect 292132 355314 292160 357734
rect 292316 357610 292344 357734
rect 292212 357604 292264 357610
rect 292212 357546 292264 357552
rect 292304 357604 292356 357610
rect 292304 357546 292356 357552
rect 292086 355286 292160 355314
rect 292086 355028 292114 355286
rect 292224 355178 292252 357546
rect 292224 355150 292344 355178
rect 292316 354674 292344 355150
rect 293040 355088 293092 355094
rect 293040 355030 293092 355036
rect 291764 354657 291884 354674
rect 292224 354657 292344 354674
rect 291750 354648 291884 354657
rect 291806 354646 291884 354648
rect 292210 354648 292344 354657
rect 291750 354583 291806 354592
rect 292266 354646 292344 354648
rect 292210 354583 292266 354592
rect 179880 351280 179932 351286
rect 179880 351222 179932 351228
rect 179510 348188 179566 348197
rect 179510 348123 179566 348132
rect 179524 347818 179552 348123
rect 179512 347812 179564 347818
rect 179512 347754 179564 347760
rect 179248 344986 179368 345014
rect 179340 341374 179368 344986
rect 179510 341388 179566 341397
rect 179340 341346 179510 341374
rect 179340 340950 179368 341346
rect 179510 341323 179566 341332
rect 179328 340944 179380 340950
rect 179328 340886 179380 340892
rect 179142 336560 179198 336569
rect 179142 336495 179198 336504
rect 179052 257372 179104 257378
rect 179052 257314 179104 257320
rect 179064 257145 179092 257314
rect 179050 257136 179106 257145
rect 179050 257071 179106 257080
rect 179050 246120 179106 246129
rect 179050 246055 179106 246064
rect 179064 224641 179092 246055
rect 179050 224632 179106 224641
rect 179050 224567 179106 224576
rect 179156 71194 179184 336495
rect 293052 328409 293080 355030
rect 293144 338745 293172 358838
rect 293224 357740 293276 357746
rect 293224 357682 293276 357688
rect 293130 338736 293186 338745
rect 293130 338671 293186 338680
rect 293236 337414 293264 357682
rect 293866 338736 293922 338745
rect 293866 338671 293922 338680
rect 293880 338162 293908 338671
rect 293868 338156 293920 338162
rect 293868 338098 293920 338104
rect 293224 337408 293276 337414
rect 293224 337350 293276 337356
rect 293972 334665 294000 367746
rect 294052 355156 294104 355162
rect 294052 355098 294104 355104
rect 293958 334656 294014 334665
rect 293958 334591 294014 334600
rect 293972 334014 294000 334591
rect 293960 334008 294012 334014
rect 293960 333950 294012 333956
rect 294064 329905 294092 355098
rect 295352 349858 295380 378762
rect 295984 367260 296036 367266
rect 295984 367202 296036 367208
rect 295340 349852 295392 349858
rect 295340 349794 295392 349800
rect 295352 349625 295380 349794
rect 295338 349616 295394 349625
rect 295338 349551 295394 349560
rect 295996 346458 296024 367202
rect 296904 364404 296956 364410
rect 296904 364346 296956 364352
rect 296812 360392 296864 360398
rect 296812 360334 296864 360340
rect 296720 359100 296772 359106
rect 296720 359042 296772 359048
rect 296166 357640 296222 357649
rect 296166 357575 296222 357584
rect 296074 354376 296130 354385
rect 296074 354311 296130 354320
rect 295984 346452 296036 346458
rect 295984 346394 296036 346400
rect 295996 345545 296024 346394
rect 295982 345536 296038 345545
rect 295982 345471 296038 345480
rect 296088 342922 296116 354311
rect 296180 352578 296208 357575
rect 296168 352572 296220 352578
rect 296168 352514 296220 352520
rect 296076 342916 296128 342922
rect 296076 342858 296128 342864
rect 295338 340776 295394 340785
rect 295338 340711 295394 340720
rect 295352 339522 295380 340711
rect 295340 339516 295392 339522
rect 295340 339458 295392 339464
rect 295340 336728 295392 336734
rect 295338 336696 295340 336705
rect 295392 336696 295394 336705
rect 295338 336631 295394 336640
rect 295338 331936 295394 331945
rect 295338 331871 295340 331880
rect 295392 331871 295394 331880
rect 295340 331842 295392 331848
rect 294050 329896 294106 329905
rect 294050 329831 294106 329840
rect 294326 329896 294382 329905
rect 294326 329831 294328 329840
rect 294380 329831 294382 329840
rect 294328 329802 294380 329808
rect 293038 328400 293094 328409
rect 293038 328335 293094 328344
rect 293052 327146 293080 328335
rect 293040 327140 293092 327146
rect 293040 327082 293092 327088
rect 294142 325816 294198 325825
rect 294142 325751 294198 325760
rect 179510 308068 179566 308077
rect 179510 308003 179566 308012
rect 179234 303920 179290 303929
rect 179234 303855 179290 303864
rect 179144 71188 179196 71194
rect 179144 71130 179196 71136
rect 177948 35352 178000 35358
rect 177948 35294 178000 35300
rect 176568 29776 176620 29782
rect 176568 29718 176620 29724
rect 179248 21554 179276 303855
rect 179326 263800 179382 263809
rect 179326 263735 179382 263744
rect 179340 79354 179368 263735
rect 179418 248160 179474 248169
rect 179418 248095 179474 248104
rect 179328 79348 179380 79354
rect 179328 79290 179380 79296
rect 179432 33930 179460 248095
rect 179524 243001 179552 308003
rect 293222 301336 293278 301345
rect 293222 301271 293278 301280
rect 293236 300898 293264 301271
rect 293224 300892 293276 300898
rect 293224 300834 293276 300840
rect 293130 287736 293186 287745
rect 293130 287671 293186 287680
rect 293038 268152 293094 268161
rect 293038 268087 293094 268096
rect 179786 244148 179842 244157
rect 179786 244083 179842 244092
rect 179510 242992 179566 243001
rect 179510 242927 179566 242936
rect 179800 241514 179828 244083
rect 179616 241486 179828 241514
rect 179512 239896 179564 239902
rect 179512 239838 179564 239844
rect 179524 38078 179552 239838
rect 179616 47598 179644 241486
rect 204258 240680 204314 240689
rect 180432 240644 180484 240650
rect 180432 240586 180484 240592
rect 184020 240644 184072 240650
rect 276294 240680 276350 240689
rect 204314 240638 204852 240666
rect 204258 240615 204314 240624
rect 184020 240586 184072 240592
rect 180030 239902 180058 240108
rect 180444 240038 180472 240586
rect 180812 240094 181976 240122
rect 183572 240094 183908 240122
rect 180432 240032 180484 240038
rect 180432 239974 180484 239980
rect 180018 239896 180070 239902
rect 180018 239838 180070 239844
rect 179604 47592 179656 47598
rect 179604 47534 179656 47540
rect 179512 38072 179564 38078
rect 179512 38014 179564 38020
rect 179420 33924 179472 33930
rect 179420 33866 179472 33872
rect 179236 21548 179288 21554
rect 179236 21490 179288 21496
rect 176476 10396 176528 10402
rect 176476 10338 176528 10344
rect 180812 6390 180840 240094
rect 180892 238808 180944 238814
rect 180892 238750 180944 238756
rect 180904 234433 180932 238750
rect 180890 234424 180946 234433
rect 180890 234359 180946 234368
rect 182824 180328 182876 180334
rect 182824 180270 182876 180276
rect 180800 6384 180852 6390
rect 180800 6326 180852 6332
rect 182836 6254 182864 180270
rect 182916 120148 182968 120154
rect 182916 120090 182968 120096
rect 182928 88194 182956 120090
rect 182916 88188 182968 88194
rect 182916 88130 182968 88136
rect 183572 13258 183600 240094
rect 184032 233170 184060 240586
rect 184952 240094 185840 240122
rect 184020 233164 184072 233170
rect 184020 233106 184072 233112
rect 184204 180260 184256 180266
rect 184204 180202 184256 180208
rect 184216 87650 184244 180202
rect 184296 121508 184348 121514
rect 184296 121450 184348 121456
rect 184204 87644 184256 87650
rect 184204 87586 184256 87592
rect 184308 86766 184336 121450
rect 184388 113280 184440 113286
rect 184388 113222 184440 113228
rect 184296 86760 184348 86766
rect 184296 86702 184348 86708
rect 184400 82618 184428 113222
rect 184388 82612 184440 82618
rect 184388 82554 184440 82560
rect 184952 68474 184980 240094
rect 187758 239850 187786 240108
rect 187712 239822 187786 239850
rect 189092 240094 190348 240122
rect 186964 232620 187016 232626
rect 186964 232562 187016 232568
rect 186976 187241 187004 232562
rect 186962 187232 187018 187241
rect 186962 187167 187018 187176
rect 185584 146396 185636 146402
rect 185584 146338 185636 146344
rect 185596 88126 185624 146338
rect 186964 140888 187016 140894
rect 186964 140830 187016 140836
rect 185676 106412 185728 106418
rect 185676 106354 185728 106360
rect 185584 88120 185636 88126
rect 185584 88062 185636 88068
rect 185688 81326 185716 106354
rect 186976 90846 187004 140830
rect 187056 120216 187108 120222
rect 187056 120158 187108 120164
rect 186964 90840 187016 90846
rect 186964 90782 187016 90788
rect 187068 83978 187096 120158
rect 187056 83972 187108 83978
rect 187056 83914 187108 83920
rect 185676 81320 185728 81326
rect 185676 81262 185728 81268
rect 184940 68468 184992 68474
rect 184940 68410 184992 68416
rect 187712 43654 187740 239822
rect 189092 231606 189120 240094
rect 192266 239850 192294 240108
rect 192220 239822 192294 239850
rect 193232 240094 194212 240122
rect 195992 240094 196144 240122
rect 192220 237153 192248 239822
rect 192206 237144 192262 237153
rect 192206 237079 192262 237088
rect 192484 236768 192536 236774
rect 192484 236710 192536 236716
rect 189080 231600 189132 231606
rect 189080 231542 189132 231548
rect 189724 231600 189776 231606
rect 189724 231542 189776 231548
rect 189736 192642 189764 231542
rect 191104 213376 191156 213382
rect 191104 213318 191156 213324
rect 189724 192636 189776 192642
rect 189724 192578 189776 192584
rect 188344 187128 188396 187134
rect 188344 187070 188396 187076
rect 188356 98666 188384 187070
rect 189724 184476 189776 184482
rect 189724 184418 189776 184424
rect 188436 138100 188488 138106
rect 188436 138042 188488 138048
rect 188344 98660 188396 98666
rect 188344 98602 188396 98608
rect 188448 92410 188476 138042
rect 188528 107704 188580 107710
rect 188528 107646 188580 107652
rect 188436 92404 188488 92410
rect 188436 92346 188488 92352
rect 188540 80034 188568 107646
rect 188528 80028 188580 80034
rect 188528 79970 188580 79976
rect 187700 43648 187752 43654
rect 187700 43590 187752 43596
rect 183560 13252 183612 13258
rect 183560 13194 183612 13200
rect 189736 9110 189764 184418
rect 189816 143608 189868 143614
rect 189816 143550 189868 143556
rect 189828 92342 189856 143550
rect 189908 110560 189960 110566
rect 189908 110502 189960 110508
rect 189816 92336 189868 92342
rect 189816 92278 189868 92284
rect 189920 78538 189948 110502
rect 191116 98734 191144 213318
rect 192496 195362 192524 236710
rect 192484 195356 192536 195362
rect 192484 195298 192536 195304
rect 192484 190528 192536 190534
rect 192484 190470 192536 190476
rect 192496 157282 192524 190470
rect 192484 157276 192536 157282
rect 192484 157218 192536 157224
rect 192484 153332 192536 153338
rect 192484 153274 192536 153280
rect 191196 104916 191248 104922
rect 191196 104858 191248 104864
rect 191104 98728 191156 98734
rect 191104 98670 191156 98676
rect 191208 94897 191236 104858
rect 191194 94888 191250 94897
rect 191194 94823 191250 94832
rect 192496 89418 192524 153274
rect 192576 131164 192628 131170
rect 192576 131106 192628 131112
rect 192484 89412 192536 89418
rect 192484 89354 192536 89360
rect 192482 84824 192538 84833
rect 192482 84759 192538 84768
rect 189908 78532 189960 78538
rect 189908 78474 189960 78480
rect 189724 9104 189776 9110
rect 189724 9046 189776 9052
rect 182824 6248 182876 6254
rect 182824 6190 182876 6196
rect 192496 3466 192524 84759
rect 192588 74458 192616 131106
rect 192668 111852 192720 111858
rect 192668 111794 192720 111800
rect 192680 85474 192708 111794
rect 192668 85468 192720 85474
rect 192668 85410 192720 85416
rect 192576 74452 192628 74458
rect 192576 74394 192628 74400
rect 193232 24274 193260 240094
rect 195992 238882 196020 240094
rect 198706 239850 198734 240108
rect 200132 240094 200652 240122
rect 201512 240094 202584 240122
rect 198706 239822 198780 239850
rect 195980 238876 196032 238882
rect 195980 238818 196032 238824
rect 195992 227186 196020 238818
rect 196624 227316 196676 227322
rect 196624 227258 196676 227264
rect 195980 227180 196032 227186
rect 195980 227122 196032 227128
rect 195244 187196 195296 187202
rect 195244 187138 195296 187144
rect 193864 145580 193916 145586
rect 193864 145522 193916 145528
rect 193876 92274 193904 145522
rect 193956 116000 194008 116006
rect 193956 115942 194008 115948
rect 193968 93158 193996 115942
rect 194048 103556 194100 103562
rect 194048 103498 194100 103504
rect 193956 93152 194008 93158
rect 193956 93094 194008 93100
rect 193864 92268 193916 92274
rect 193864 92210 193916 92216
rect 194060 89729 194088 103498
rect 194046 89720 194102 89729
rect 194046 89655 194102 89664
rect 193220 24268 193272 24274
rect 193220 24210 193272 24216
rect 195256 20126 195284 187138
rect 195336 117360 195388 117366
rect 195336 117302 195388 117308
rect 195348 90982 195376 117302
rect 195336 90976 195388 90982
rect 195336 90918 195388 90924
rect 195244 20120 195296 20126
rect 195244 20062 195296 20068
rect 196636 3466 196664 227258
rect 198004 227248 198056 227254
rect 198004 227190 198056 227196
rect 196716 195492 196768 195498
rect 196716 195434 196768 195440
rect 196728 177478 196756 195434
rect 198016 191185 198044 227190
rect 198002 191176 198058 191185
rect 198002 191111 198058 191120
rect 198004 181484 198056 181490
rect 198004 181426 198056 181432
rect 196716 177472 196768 177478
rect 196716 177414 196768 177420
rect 196716 128444 196768 128450
rect 196716 128386 196768 128392
rect 196728 78606 196756 128386
rect 196808 125724 196860 125730
rect 196808 125666 196860 125672
rect 196820 81190 196848 125666
rect 196808 81184 196860 81190
rect 196808 81126 196860 81132
rect 196716 78600 196768 78606
rect 196716 78542 196768 78548
rect 198016 4894 198044 181426
rect 198096 127628 198148 127634
rect 198096 127570 198148 127576
rect 198108 96626 198136 127570
rect 198280 103624 198332 103630
rect 198280 103566 198332 103572
rect 198188 102196 198240 102202
rect 198188 102138 198240 102144
rect 198096 96620 198148 96626
rect 198096 96562 198148 96568
rect 198200 86902 198228 102138
rect 198292 91050 198320 103566
rect 198752 91798 198780 239822
rect 199384 111920 199436 111926
rect 199384 111862 199436 111868
rect 198740 91792 198792 91798
rect 198740 91734 198792 91740
rect 198280 91044 198332 91050
rect 198280 90986 198332 90992
rect 198188 86896 198240 86902
rect 198188 86838 198240 86844
rect 199396 75886 199424 111862
rect 200132 77994 200160 240094
rect 200764 102264 200816 102270
rect 200764 102206 200816 102212
rect 200776 89690 200804 102206
rect 200764 89684 200816 89690
rect 200764 89626 200816 89632
rect 200120 77988 200172 77994
rect 200120 77930 200172 77936
rect 199384 75880 199436 75886
rect 199384 75822 199436 75828
rect 201512 43586 201540 240094
rect 204824 238406 204852 240638
rect 276294 240615 276350 240624
rect 291936 240644 291988 240650
rect 276308 240530 276336 240615
rect 291936 240586 291988 240592
rect 276000 240502 276336 240530
rect 207092 240094 207428 240122
rect 204812 238400 204864 238406
rect 204812 238342 204864 238348
rect 207400 237425 207428 240094
rect 208412 240094 209024 240122
rect 210436 240094 210956 240122
rect 212552 240094 212888 240122
rect 215220 240094 215464 240122
rect 216692 240094 217396 240122
rect 207386 237416 207442 237425
rect 207386 237351 207442 237360
rect 202142 235240 202198 235249
rect 202142 235175 202198 235184
rect 202156 213382 202184 235175
rect 206282 232656 206338 232665
rect 206282 232591 206338 232600
rect 203616 229900 203668 229906
rect 203616 229842 203668 229848
rect 202144 213376 202196 213382
rect 202144 213318 202196 213324
rect 203524 210656 203576 210662
rect 203524 210598 203576 210604
rect 202236 151904 202288 151910
rect 202236 151846 202288 151852
rect 202144 139460 202196 139466
rect 202144 139402 202196 139408
rect 202156 78470 202184 139402
rect 202248 93294 202276 151846
rect 202236 93288 202288 93294
rect 202236 93230 202288 93236
rect 202144 78464 202196 78470
rect 202144 78406 202196 78412
rect 201500 43580 201552 43586
rect 201500 43522 201552 43528
rect 203536 14550 203564 210598
rect 203628 181490 203656 229842
rect 203616 181484 203668 181490
rect 203616 181426 203668 181432
rect 205640 151088 205692 151094
rect 205640 151030 205692 151036
rect 203616 150476 203668 150482
rect 203616 150418 203668 150424
rect 203628 122126 203656 150418
rect 205652 150346 205680 151030
rect 205640 150340 205692 150346
rect 205640 150282 205692 150288
rect 204904 145036 204956 145042
rect 204904 144978 204956 144984
rect 203616 122120 203668 122126
rect 203616 122062 203668 122068
rect 203616 117428 203668 117434
rect 203616 117370 203668 117376
rect 203628 86834 203656 117370
rect 203708 104984 203760 104990
rect 203708 104926 203760 104932
rect 203720 88262 203748 104926
rect 204916 91866 204944 144978
rect 205088 105052 205140 105058
rect 205088 104994 205140 105000
rect 204996 100768 205048 100774
rect 204996 100710 205048 100716
rect 204904 91860 204956 91866
rect 204904 91802 204956 91808
rect 203708 88256 203760 88262
rect 203708 88198 203760 88204
rect 203616 86828 203668 86834
rect 203616 86770 203668 86776
rect 205008 73166 205036 100710
rect 205100 93838 205128 104994
rect 205088 93832 205140 93838
rect 205088 93774 205140 93780
rect 206296 88330 206324 232591
rect 207664 221536 207716 221542
rect 207664 221478 207716 221484
rect 206376 182300 206428 182306
rect 206376 182242 206428 182248
rect 206388 173806 206416 182242
rect 206376 173800 206428 173806
rect 206376 173742 206428 173748
rect 206374 171728 206430 171737
rect 206374 171663 206430 171672
rect 206388 93158 206416 171663
rect 206468 127016 206520 127022
rect 206468 126958 206520 126964
rect 206376 93152 206428 93158
rect 206376 93094 206428 93100
rect 206284 88324 206336 88330
rect 206284 88266 206336 88272
rect 206480 84182 206508 126958
rect 206560 121576 206612 121582
rect 206560 121518 206612 121524
rect 206468 84176 206520 84182
rect 206468 84118 206520 84124
rect 206572 79898 206600 121518
rect 207676 95130 207704 221478
rect 207756 133952 207808 133958
rect 207756 133894 207808 133900
rect 207664 95124 207716 95130
rect 207664 95066 207716 95072
rect 207768 82686 207796 133894
rect 207848 107772 207900 107778
rect 207848 107714 207900 107720
rect 207860 93226 207888 107714
rect 207940 96688 207992 96694
rect 207940 96630 207992 96636
rect 207848 93220 207900 93226
rect 207848 93162 207900 93168
rect 207952 87990 207980 96630
rect 207940 87984 207992 87990
rect 207940 87926 207992 87932
rect 207756 82680 207808 82686
rect 207756 82622 207808 82628
rect 206560 79892 206612 79898
rect 206560 79834 206612 79840
rect 204996 73160 205048 73166
rect 204996 73102 205048 73108
rect 208412 32570 208440 240094
rect 210436 238542 210464 240094
rect 210424 238536 210476 238542
rect 210424 238478 210476 238484
rect 210436 189922 210464 238478
rect 211896 221672 211948 221678
rect 211896 221614 211948 221620
rect 209044 189916 209096 189922
rect 209044 189858 209096 189864
rect 210424 189916 210476 189922
rect 210424 189858 210476 189864
rect 209056 180266 209084 189858
rect 211068 181620 211120 181626
rect 211068 181562 211120 181568
rect 209044 180260 209096 180266
rect 209044 180202 209096 180208
rect 210424 179444 210476 179450
rect 210424 179386 210476 179392
rect 210436 164150 210464 179386
rect 210424 164144 210476 164150
rect 210424 164086 210476 164092
rect 210516 142724 210568 142730
rect 210516 142666 210568 142672
rect 210424 114640 210476 114646
rect 210424 114582 210476 114588
rect 209044 109132 209096 109138
rect 209044 109074 209096 109080
rect 209056 82754 209084 109074
rect 210436 84114 210464 114582
rect 210424 84108 210476 84114
rect 210424 84050 210476 84056
rect 209044 82748 209096 82754
rect 209044 82690 209096 82696
rect 210528 81258 210556 142666
rect 210608 118856 210660 118862
rect 210608 118798 210660 118804
rect 210620 89622 210648 118798
rect 210608 89616 210660 89622
rect 210608 89558 210660 89564
rect 210516 81252 210568 81258
rect 210516 81194 210568 81200
rect 210424 80708 210476 80714
rect 210424 80650 210476 80656
rect 208400 32564 208452 32570
rect 208400 32506 208452 32512
rect 203524 14544 203576 14550
rect 203524 14486 203576 14492
rect 198004 4888 198056 4894
rect 198004 4830 198056 4836
rect 210436 3602 210464 80650
rect 211080 3670 211108 181562
rect 211802 180024 211858 180033
rect 211802 179959 211858 179968
rect 211816 6322 211844 179959
rect 211908 178770 211936 221614
rect 211988 184952 212040 184958
rect 211988 184894 212040 184900
rect 211896 178764 211948 178770
rect 211896 178706 211948 178712
rect 212000 168298 212028 184894
rect 211988 168292 212040 168298
rect 211988 168234 212040 168240
rect 211896 150544 211948 150550
rect 211896 150486 211948 150492
rect 211908 140078 211936 150486
rect 212080 143676 212132 143682
rect 212080 143618 212132 143624
rect 211896 140072 211948 140078
rect 211896 140014 211948 140020
rect 211988 139528 212040 139534
rect 211988 139470 212040 139476
rect 211896 89004 211948 89010
rect 211896 88946 211948 88952
rect 211804 6316 211856 6322
rect 211804 6258 211856 6264
rect 211068 3664 211120 3670
rect 211068 3606 211120 3612
rect 210424 3596 210476 3602
rect 210424 3538 210476 3544
rect 211908 3534 211936 88946
rect 212000 79966 212028 139470
rect 212092 89554 212120 143618
rect 212172 118788 212224 118794
rect 212172 118730 212224 118736
rect 212080 89548 212132 89554
rect 212080 89490 212132 89496
rect 212184 85542 212212 118730
rect 212172 85536 212224 85542
rect 212172 85478 212224 85484
rect 212552 83502 212580 240094
rect 215220 239465 215248 240094
rect 215206 239456 215262 239465
rect 215206 239391 215262 239400
rect 215220 231606 215248 239391
rect 215208 231600 215260 231606
rect 215208 231542 215260 231548
rect 214564 182232 214616 182238
rect 214564 182174 214616 182180
rect 214196 178084 214248 178090
rect 214196 178026 214248 178032
rect 213920 176656 213972 176662
rect 213920 176598 213972 176604
rect 213932 175681 213960 176598
rect 213918 175672 213974 175681
rect 213918 175607 213974 175616
rect 214012 175228 214064 175234
rect 214012 175170 214064 175176
rect 213920 175160 213972 175166
rect 213920 175102 213972 175108
rect 213932 175001 213960 175102
rect 213918 174992 213974 175001
rect 213918 174927 213974 174936
rect 214024 174321 214052 175170
rect 214104 174548 214156 174554
rect 214104 174490 214156 174496
rect 214010 174312 214066 174321
rect 214010 174247 214066 174256
rect 213920 173868 213972 173874
rect 213920 173810 213972 173816
rect 213932 173641 213960 173810
rect 214012 173800 214064 173806
rect 214012 173742 214064 173748
rect 213918 173632 213974 173641
rect 213918 173567 213974 173576
rect 214024 172961 214052 173742
rect 214010 172952 214066 172961
rect 214010 172887 214066 172896
rect 214116 171601 214144 174490
rect 214208 172281 214236 178026
rect 214194 172272 214250 172281
rect 214194 172207 214250 172216
rect 214102 171592 214158 171601
rect 214102 171527 214158 171536
rect 213920 171080 213972 171086
rect 213920 171022 213972 171028
rect 213932 170377 213960 171022
rect 213918 170368 213974 170377
rect 213918 170303 213974 170312
rect 213920 169720 213972 169726
rect 213918 169688 213920 169697
rect 213972 169688 213974 169697
rect 213918 169623 213974 169632
rect 214012 169652 214064 169658
rect 214012 169594 214064 169600
rect 214024 169017 214052 169594
rect 214010 169008 214066 169017
rect 214010 168943 214066 168952
rect 213920 168360 213972 168366
rect 213920 168302 213972 168308
rect 214010 168328 214066 168337
rect 213932 167657 213960 168302
rect 214010 168263 214012 168272
rect 214064 168263 214066 168272
rect 214012 168234 214064 168240
rect 213918 167648 213974 167657
rect 213918 167583 213974 167592
rect 214104 167000 214156 167006
rect 213918 166968 213974 166977
rect 214104 166942 214156 166948
rect 213918 166903 213974 166912
rect 214012 166932 214064 166938
rect 213932 166870 213960 166903
rect 214012 166874 214064 166880
rect 213920 166864 213972 166870
rect 213920 166806 213972 166812
rect 214024 165753 214052 166874
rect 214116 166433 214144 166942
rect 214102 166424 214158 166433
rect 214102 166359 214158 166368
rect 214010 165744 214066 165753
rect 214010 165679 214066 165688
rect 213920 165572 213972 165578
rect 213920 165514 213972 165520
rect 213932 165073 213960 165514
rect 213918 165064 213974 165073
rect 213918 164999 213974 165008
rect 213920 164212 213972 164218
rect 213920 164154 213972 164160
rect 213932 163033 213960 164154
rect 214012 164144 214064 164150
rect 214012 164086 214064 164092
rect 214024 163713 214052 164086
rect 214010 163704 214066 163713
rect 214010 163639 214066 163648
rect 213918 163024 213974 163033
rect 213918 162959 213974 162968
rect 213920 162852 213972 162858
rect 213920 162794 213972 162800
rect 213932 161809 213960 162794
rect 214576 162353 214604 182174
rect 214656 180872 214708 180878
rect 214656 180814 214708 180820
rect 214668 175930 214696 180814
rect 215944 177540 215996 177546
rect 215944 177482 215996 177488
rect 214668 175902 214788 175930
rect 214656 171828 214708 171834
rect 214656 171770 214708 171776
rect 214562 162344 214618 162353
rect 214562 162279 214618 162288
rect 213918 161800 213974 161809
rect 213918 161735 213974 161744
rect 214668 161474 214696 171770
rect 214760 171057 214788 175902
rect 214746 171048 214802 171057
rect 214746 170983 214802 170992
rect 214668 161446 214972 161474
rect 213920 161424 213972 161430
rect 213920 161366 213972 161372
rect 213932 161129 213960 161366
rect 214012 161356 214064 161362
rect 214012 161298 214064 161304
rect 213918 161120 213974 161129
rect 213918 161055 213974 161064
rect 214024 160449 214052 161298
rect 214010 160440 214066 160449
rect 214010 160375 214066 160384
rect 213920 160064 213972 160070
rect 213920 160006 213972 160012
rect 213932 159089 213960 160006
rect 213918 159080 213974 159089
rect 213918 159015 213974 159024
rect 213920 158704 213972 158710
rect 213920 158646 213972 158652
rect 213932 158409 213960 158646
rect 213918 158400 213974 158409
rect 213918 158335 213974 158344
rect 214944 157729 214972 161446
rect 214930 157720 214986 157729
rect 214930 157655 214986 157664
rect 214012 157344 214064 157350
rect 214012 157286 214064 157292
rect 213920 157276 213972 157282
rect 213920 157218 213972 157224
rect 213932 157185 213960 157218
rect 213918 157176 213974 157185
rect 213918 157111 213974 157120
rect 214024 156505 214052 157286
rect 214010 156496 214066 156505
rect 214010 156431 214066 156440
rect 213920 155916 213972 155922
rect 213920 155858 213972 155864
rect 213932 155825 213960 155858
rect 213918 155816 213974 155825
rect 213918 155751 213974 155760
rect 214010 154456 214066 154465
rect 214010 154391 214066 154400
rect 213918 153776 213974 153785
rect 213918 153711 213974 153720
rect 213932 153338 213960 153711
rect 213920 153332 213972 153338
rect 213920 153274 213972 153280
rect 214024 153270 214052 154391
rect 214012 153264 214064 153270
rect 214012 153206 214064 153212
rect 213918 153096 213974 153105
rect 213918 153031 213974 153040
rect 213932 151910 213960 153031
rect 214010 152552 214066 152561
rect 214010 152487 214066 152496
rect 213920 151904 213972 151910
rect 213920 151846 213972 151852
rect 214024 151842 214052 152487
rect 214654 151872 214710 151881
rect 214012 151836 214064 151842
rect 214654 151814 214710 151816
rect 214654 151807 214788 151814
rect 214668 151786 214788 151807
rect 214012 151778 214064 151784
rect 214010 151192 214066 151201
rect 214010 151127 214066 151136
rect 214024 150550 214052 151127
rect 214012 150544 214064 150550
rect 213918 150512 213974 150521
rect 214012 150486 214064 150492
rect 213918 150447 213920 150456
rect 213972 150447 213974 150456
rect 213920 150418 213972 150424
rect 214012 150408 214064 150414
rect 214012 150350 214064 150356
rect 213920 150340 213972 150346
rect 213920 150282 213972 150288
rect 213932 149161 213960 150282
rect 214024 149841 214052 150350
rect 214010 149832 214066 149841
rect 214010 149767 214066 149776
rect 213918 149152 213974 149161
rect 213918 149087 213974 149096
rect 213920 149048 213972 149054
rect 213920 148990 213972 148996
rect 213932 148481 213960 148990
rect 213918 148472 213974 148481
rect 213918 148407 213974 148416
rect 214102 147928 214158 147937
rect 214102 147863 214158 147872
rect 214010 147248 214066 147257
rect 214010 147183 214066 147192
rect 213918 146568 213974 146577
rect 213918 146503 213974 146512
rect 213932 146402 213960 146503
rect 213920 146396 213972 146402
rect 213920 146338 213972 146344
rect 214024 146334 214052 147183
rect 214012 146328 214064 146334
rect 214012 146270 214064 146276
rect 214010 145888 214066 145897
rect 214010 145823 214066 145832
rect 213918 145208 213974 145217
rect 213918 145143 213974 145152
rect 213932 144974 213960 145143
rect 214024 145042 214052 145823
rect 214116 145586 214144 147863
rect 214104 145580 214156 145586
rect 214104 145522 214156 145528
rect 214012 145036 214064 145042
rect 214012 144978 214064 144984
rect 213920 144968 213972 144974
rect 213920 144910 213972 144916
rect 213918 144528 213974 144537
rect 213918 144463 213974 144472
rect 213932 143614 213960 144463
rect 214654 143848 214710 143857
rect 214654 143783 214710 143792
rect 214668 143682 214696 143783
rect 214656 143676 214708 143682
rect 214656 143618 214708 143624
rect 213920 143608 213972 143614
rect 213920 143550 213972 143556
rect 213918 143304 213974 143313
rect 213918 143239 213974 143248
rect 213932 142730 213960 143239
rect 213920 142724 213972 142730
rect 213920 142666 213972 142672
rect 214562 142624 214618 142633
rect 214562 142559 214618 142568
rect 214010 141944 214066 141953
rect 214010 141879 214066 141888
rect 213918 141264 213974 141273
rect 213918 141199 213974 141208
rect 213932 140826 213960 141199
rect 214024 140894 214052 141879
rect 214012 140888 214064 140894
rect 214012 140830 214064 140836
rect 213920 140820 213972 140826
rect 213920 140762 213972 140768
rect 213918 140584 213974 140593
rect 213918 140519 213974 140528
rect 213932 139466 213960 140519
rect 213920 139460 213972 139466
rect 213920 139402 213972 139408
rect 214010 139224 214066 139233
rect 214010 139159 214066 139168
rect 213918 138680 213974 138689
rect 213918 138615 213974 138624
rect 213932 138106 213960 138615
rect 213920 138100 213972 138106
rect 213920 138042 213972 138048
rect 214024 138038 214052 139159
rect 214012 138032 214064 138038
rect 214012 137974 214064 137980
rect 214010 135960 214066 135969
rect 214010 135895 214066 135904
rect 213920 135380 213972 135386
rect 213920 135322 213972 135328
rect 213932 135289 213960 135322
rect 214024 135318 214052 135895
rect 214012 135312 214064 135318
rect 213918 135280 213974 135289
rect 214012 135254 214064 135260
rect 213918 135215 213974 135224
rect 213918 134600 213974 134609
rect 213918 134535 213974 134544
rect 213932 133958 213960 134535
rect 213920 133952 213972 133958
rect 213920 133894 213972 133900
rect 213918 133376 213974 133385
rect 213918 133311 213974 133320
rect 213932 132530 213960 133311
rect 213920 132524 213972 132530
rect 213920 132466 213972 132472
rect 213918 131336 213974 131345
rect 213918 131271 213974 131280
rect 213932 131170 213960 131271
rect 213920 131164 213972 131170
rect 213920 131106 213972 131112
rect 214010 129296 214066 129305
rect 214010 129231 214066 129240
rect 213918 128752 213974 128761
rect 213918 128687 213974 128696
rect 213932 128382 213960 128687
rect 214024 128450 214052 129231
rect 214012 128444 214064 128450
rect 214012 128386 214064 128392
rect 213920 128376 213972 128382
rect 213920 128318 213972 128324
rect 213918 128072 213974 128081
rect 213918 128007 213974 128016
rect 213932 127022 213960 128007
rect 213920 127016 213972 127022
rect 213920 126958 213972 126964
rect 214010 126712 214066 126721
rect 214010 126647 214066 126656
rect 213918 126032 213974 126041
rect 213918 125967 213974 125976
rect 213932 125662 213960 125967
rect 214024 125730 214052 126647
rect 214012 125724 214064 125730
rect 214012 125666 214064 125672
rect 213920 125656 213972 125662
rect 213920 125598 213972 125604
rect 214010 125352 214066 125361
rect 214010 125287 214066 125296
rect 213918 124672 213974 124681
rect 213918 124607 213974 124616
rect 213932 124302 213960 124607
rect 213920 124296 213972 124302
rect 213920 124238 213972 124244
rect 214024 124234 214052 125287
rect 214012 124228 214064 124234
rect 214012 124170 214064 124176
rect 214010 124128 214066 124137
rect 214010 124063 214066 124072
rect 213918 123448 213974 123457
rect 213918 123383 213974 123392
rect 213932 122942 213960 123383
rect 213920 122936 213972 122942
rect 213920 122878 213972 122884
rect 214024 122874 214052 124063
rect 214012 122868 214064 122874
rect 214012 122810 214064 122816
rect 214010 122768 214066 122777
rect 214010 122703 214066 122712
rect 213918 122088 213974 122097
rect 213918 122023 213974 122032
rect 213932 121514 213960 122023
rect 214024 121582 214052 122703
rect 214012 121576 214064 121582
rect 214012 121518 214064 121524
rect 213920 121508 213972 121514
rect 213920 121450 213972 121456
rect 214010 121408 214066 121417
rect 214010 121343 214066 121352
rect 213918 120728 213974 120737
rect 213918 120663 213974 120672
rect 213932 120222 213960 120663
rect 213920 120216 213972 120222
rect 213920 120158 213972 120164
rect 214024 120154 214052 121343
rect 214012 120148 214064 120154
rect 214012 120090 214064 120096
rect 214102 120048 214158 120057
rect 214102 119983 214158 119992
rect 214010 119504 214066 119513
rect 214010 119439 214066 119448
rect 213918 118824 213974 118833
rect 214024 118794 214052 119439
rect 214116 118862 214144 119983
rect 214104 118856 214156 118862
rect 214104 118798 214156 118804
rect 213918 118759 213974 118768
rect 214012 118788 214064 118794
rect 213932 118726 213960 118759
rect 214012 118730 214064 118736
rect 213920 118720 213972 118726
rect 213920 118662 213972 118668
rect 214010 118144 214066 118153
rect 214010 118079 214066 118088
rect 213918 117464 213974 117473
rect 213918 117399 213920 117408
rect 213972 117399 213974 117408
rect 213920 117370 213972 117376
rect 214024 117366 214052 118079
rect 214012 117360 214064 117366
rect 214012 117302 214064 117308
rect 213182 116784 213238 116793
rect 213182 116719 213238 116728
rect 212540 83496 212592 83502
rect 212540 83438 212592 83444
rect 211988 79960 212040 79966
rect 211988 79902 212040 79908
rect 213196 78674 213224 116719
rect 213918 116104 213974 116113
rect 213918 116039 213974 116048
rect 213932 116006 213960 116039
rect 213920 116000 213972 116006
rect 213920 115942 213972 115948
rect 214010 115424 214066 115433
rect 214010 115359 214066 115368
rect 213918 114880 213974 114889
rect 213918 114815 213974 114824
rect 213932 114578 213960 114815
rect 214024 114646 214052 115359
rect 214012 114640 214064 114646
rect 214012 114582 214064 114588
rect 213920 114572 213972 114578
rect 213920 114514 213972 114520
rect 214010 114200 214066 114209
rect 214010 114135 214066 114144
rect 213918 113520 213974 113529
rect 213918 113455 213974 113464
rect 213932 113286 213960 113455
rect 213920 113280 213972 113286
rect 213920 113222 213972 113228
rect 214024 113218 214052 114135
rect 214012 113212 214064 113218
rect 214012 113154 214064 113160
rect 214010 112840 214066 112849
rect 214010 112775 214066 112784
rect 213918 112160 213974 112169
rect 213918 112095 213974 112104
rect 213932 111926 213960 112095
rect 213920 111920 213972 111926
rect 213920 111862 213972 111868
rect 214024 111858 214052 112775
rect 214012 111852 214064 111858
rect 214012 111794 214064 111800
rect 214010 111480 214066 111489
rect 214010 111415 214066 111424
rect 213918 110800 213974 110809
rect 213918 110735 213974 110744
rect 213932 110566 213960 110735
rect 213920 110560 213972 110566
rect 213920 110502 213972 110508
rect 214024 110498 214052 111415
rect 214012 110492 214064 110498
rect 214012 110434 214064 110440
rect 214010 110256 214066 110265
rect 214010 110191 214066 110200
rect 213918 109576 213974 109585
rect 213918 109511 213974 109520
rect 213932 109070 213960 109511
rect 214024 109138 214052 110191
rect 214012 109132 214064 109138
rect 214012 109074 214064 109080
rect 213920 109064 213972 109070
rect 213920 109006 213972 109012
rect 214010 108896 214066 108905
rect 214010 108831 214066 108840
rect 213918 108216 213974 108225
rect 213918 108151 213974 108160
rect 213932 107778 213960 108151
rect 213920 107772 213972 107778
rect 213920 107714 213972 107720
rect 214024 107710 214052 108831
rect 214012 107704 214064 107710
rect 214012 107646 214064 107652
rect 214010 107536 214066 107545
rect 214010 107471 214066 107480
rect 213918 106856 213974 106865
rect 213918 106791 213974 106800
rect 213932 106418 213960 106791
rect 213920 106412 213972 106418
rect 213920 106354 213972 106360
rect 214024 106350 214052 107471
rect 214012 106344 214064 106350
rect 214012 106286 214064 106292
rect 214010 106176 214066 106185
rect 214010 106111 214066 106120
rect 213920 105052 213972 105058
rect 213920 104994 213972 105000
rect 213932 104961 213960 104994
rect 214024 104990 214052 106111
rect 214102 105632 214158 105641
rect 214102 105567 214158 105576
rect 214012 104984 214064 104990
rect 213918 104952 213974 104961
rect 214012 104926 214064 104932
rect 214116 104922 214144 105567
rect 213918 104887 213974 104896
rect 214104 104916 214156 104922
rect 214104 104858 214156 104864
rect 214010 104272 214066 104281
rect 214010 104207 214066 104216
rect 213920 103624 213972 103630
rect 213918 103592 213920 103601
rect 213972 103592 213974 103601
rect 214024 103562 214052 104207
rect 213918 103527 213974 103536
rect 214012 103556 214064 103562
rect 214576 103514 214604 142559
rect 214654 139904 214710 139913
rect 214654 139839 214710 139848
rect 214668 139534 214696 139839
rect 214656 139528 214708 139534
rect 214656 139470 214708 139476
rect 214654 137320 214710 137329
rect 214760 137290 214788 151786
rect 214654 137255 214710 137264
rect 214748 137284 214800 137290
rect 214668 108338 214696 137255
rect 214748 137226 214800 137232
rect 214746 136640 214802 136649
rect 214746 136575 214802 136584
rect 214760 108458 214788 136575
rect 214748 108452 214800 108458
rect 214748 108394 214800 108400
rect 214668 108310 214880 108338
rect 214656 108248 214708 108254
rect 214656 108190 214708 108196
rect 214012 103498 214064 103504
rect 214392 103486 214604 103514
rect 214010 102912 214066 102921
rect 214010 102847 214066 102856
rect 214024 102270 214052 102847
rect 214012 102264 214064 102270
rect 213918 102232 213974 102241
rect 214012 102206 214064 102212
rect 213918 102167 213920 102176
rect 213972 102167 213974 102176
rect 213920 102138 213972 102144
rect 213918 101008 213974 101017
rect 213918 100943 213974 100952
rect 213932 100774 213960 100943
rect 213920 100768 213972 100774
rect 213920 100710 213972 100716
rect 214010 100328 214066 100337
rect 214010 100263 214066 100272
rect 213918 98968 213974 98977
rect 213918 98903 213974 98912
rect 213932 98054 213960 98903
rect 213920 98048 213972 98054
rect 213920 97990 213972 97996
rect 213918 97608 213974 97617
rect 213918 97543 213974 97552
rect 213932 96694 213960 97543
rect 213920 96688 213972 96694
rect 213920 96630 213972 96636
rect 213918 96384 213974 96393
rect 213918 96319 213974 96328
rect 213932 95266 213960 96319
rect 214024 95946 214052 100263
rect 214392 100026 214420 103486
rect 214668 100094 214696 108190
rect 214852 103514 214880 108310
rect 214852 103486 214972 103514
rect 214656 100088 214708 100094
rect 214656 100030 214708 100036
rect 214380 100020 214432 100026
rect 214380 99962 214432 99968
rect 214102 99648 214158 99657
rect 214102 99583 214158 99592
rect 214012 95940 214064 95946
rect 214012 95882 214064 95888
rect 213920 95260 213972 95266
rect 213920 95202 213972 95208
rect 214116 94518 214144 99583
rect 214562 98288 214618 98297
rect 214562 98223 214618 98232
rect 214104 94512 214156 94518
rect 214104 94454 214156 94460
rect 213184 78668 213236 78674
rect 213184 78610 213236 78616
rect 214576 74526 214604 98223
rect 214944 97209 214972 103486
rect 214930 97200 214986 97209
rect 214930 97135 214986 97144
rect 214838 96928 214894 96937
rect 214838 96863 214894 96872
rect 214852 86970 214880 96863
rect 214840 86964 214892 86970
rect 214840 86906 214892 86912
rect 214564 74520 214616 74526
rect 214564 74462 214616 74468
rect 215956 3534 215984 177482
rect 216036 160744 216088 160750
rect 216036 160686 216088 160692
rect 216048 3602 216076 160686
rect 216128 148368 216180 148374
rect 216128 148310 216180 148316
rect 216140 3738 216168 148310
rect 216692 11898 216720 240094
rect 219314 239850 219342 240108
rect 219268 239822 219342 239850
rect 220832 240094 221260 240122
rect 223592 240094 223836 240122
rect 224972 240094 225768 240122
rect 219268 234530 219296 239822
rect 219256 234524 219308 234530
rect 219256 234466 219308 234472
rect 220084 222964 220136 222970
rect 220084 222906 220136 222912
rect 220096 178838 220124 222906
rect 220832 181626 220860 240094
rect 223592 228886 223620 240094
rect 223580 228880 223632 228886
rect 223580 228822 223632 228828
rect 222844 225616 222896 225622
rect 222844 225558 222896 225564
rect 222856 181694 222884 225558
rect 224972 205154 225000 240094
rect 227686 239850 227714 240108
rect 229112 240094 229632 240122
rect 231872 240094 232208 240122
rect 233896 240094 234140 240122
rect 236072 240094 236316 240122
rect 227686 239822 227760 239850
rect 225604 205216 225656 205222
rect 225604 205158 225656 205164
rect 224960 205148 225012 205154
rect 224960 205090 225012 205096
rect 222844 181688 222896 181694
rect 222844 181630 222896 181636
rect 225616 181626 225644 205158
rect 227732 194002 227760 239822
rect 227720 193996 227772 194002
rect 227720 193938 227772 193944
rect 229112 189825 229140 240094
rect 229744 210724 229796 210730
rect 229744 210666 229796 210672
rect 229098 189816 229154 189825
rect 229098 189751 229154 189760
rect 229756 183025 229784 210666
rect 231872 191418 231900 240094
rect 233896 238241 233924 240094
rect 236288 238513 236316 240094
rect 237392 240094 238004 240122
rect 236274 238504 236330 238513
rect 236274 238439 236330 238448
rect 233882 238232 233938 238241
rect 233882 238167 233938 238176
rect 233896 230314 233924 238167
rect 236288 238066 236316 238439
rect 236276 238060 236328 238066
rect 236276 238002 236328 238008
rect 233884 230308 233936 230314
rect 233884 230250 233936 230256
rect 233884 217388 233936 217394
rect 233884 217330 233936 217336
rect 232504 202360 232556 202366
rect 232504 202302 232556 202308
rect 231860 191412 231912 191418
rect 231860 191354 231912 191360
rect 229742 183016 229798 183025
rect 229742 182951 229798 182960
rect 220820 181620 220872 181626
rect 220820 181562 220872 181568
rect 225604 181620 225656 181626
rect 225604 181562 225656 181568
rect 220084 178832 220136 178838
rect 220084 178774 220136 178780
rect 232516 175953 232544 202302
rect 233896 177585 233924 217330
rect 235264 203788 235316 203794
rect 235264 203730 235316 203736
rect 233976 198280 234028 198286
rect 233976 198222 234028 198228
rect 233988 178906 234016 198222
rect 233976 178900 234028 178906
rect 233976 178842 234028 178848
rect 233882 177576 233938 177585
rect 233882 177511 233938 177520
rect 235276 176662 235304 203730
rect 237392 183054 237420 240094
rect 240566 239850 240594 240108
rect 240520 239822 240594 239850
rect 242268 240094 242512 240122
rect 244292 240094 244444 240122
rect 245672 240094 246376 240122
rect 248432 240094 248952 240122
rect 240520 238649 240548 239822
rect 240506 238640 240562 238649
rect 240506 238575 240562 238584
rect 240520 238474 240548 238575
rect 240508 238468 240560 238474
rect 240508 238410 240560 238416
rect 242268 233986 242296 240094
rect 242256 233980 242308 233986
rect 242256 233922 242308 233928
rect 242164 229832 242216 229838
rect 242164 229774 242216 229780
rect 242176 216646 242204 229774
rect 242268 229022 242296 233922
rect 242256 229016 242308 229022
rect 242256 228958 242308 228964
rect 243544 225684 243596 225690
rect 243544 225626 243596 225632
rect 242164 216640 242216 216646
rect 242164 216582 242216 216588
rect 238024 213240 238076 213246
rect 238024 213182 238076 213188
rect 237380 183048 237432 183054
rect 237380 182990 237432 182996
rect 238036 181665 238064 213182
rect 242164 212016 242216 212022
rect 242164 211958 242216 211964
rect 240784 209296 240836 209302
rect 240784 209238 240836 209244
rect 238116 205012 238168 205018
rect 238116 204954 238168 204960
rect 238022 181656 238078 181665
rect 238022 181591 238078 181600
rect 238128 180334 238156 204954
rect 239404 202428 239456 202434
rect 239404 202370 239456 202376
rect 238116 180328 238168 180334
rect 238116 180270 238168 180276
rect 239416 177546 239444 202370
rect 240796 180402 240824 209238
rect 242176 180470 242204 211958
rect 242256 191276 242308 191282
rect 242256 191218 242308 191224
rect 242164 180464 242216 180470
rect 242164 180406 242216 180412
rect 240784 180396 240836 180402
rect 240784 180338 240836 180344
rect 242268 177614 242296 191218
rect 243556 188630 243584 225626
rect 243544 188624 243596 188630
rect 243544 188566 243596 188572
rect 243544 185904 243596 185910
rect 243544 185846 243596 185852
rect 242256 177608 242308 177614
rect 242256 177550 242308 177556
rect 239404 177540 239456 177546
rect 239404 177482 239456 177488
rect 235264 176656 235316 176662
rect 235264 176598 235316 176604
rect 232502 175944 232558 175953
rect 232502 175879 232558 175888
rect 243556 175846 243584 185846
rect 244292 177449 244320 240094
rect 245672 202366 245700 240094
rect 246304 231192 246356 231198
rect 246304 231134 246356 231140
rect 245660 202360 245712 202366
rect 245660 202302 245712 202308
rect 246316 192914 246344 231134
rect 247684 221604 247736 221610
rect 247684 221546 247736 221552
rect 246304 192908 246356 192914
rect 246304 192850 246356 192856
rect 246396 192772 246448 192778
rect 246396 192714 246448 192720
rect 246304 188556 246356 188562
rect 246304 188498 246356 188504
rect 244278 177440 244334 177449
rect 244278 177375 244334 177384
rect 246316 176594 246344 188498
rect 246408 179217 246436 192714
rect 246488 190052 246540 190058
rect 246488 189994 246540 190000
rect 246394 179208 246450 179217
rect 246394 179143 246450 179152
rect 246500 179042 246528 189994
rect 246488 179036 246540 179042
rect 246488 178978 246540 178984
rect 246304 176588 246356 176594
rect 246304 176530 246356 176536
rect 247696 176089 247724 221546
rect 248432 217394 248460 240094
rect 250870 239850 250898 240108
rect 252816 240094 253152 240122
rect 250824 239822 250898 239850
rect 250824 238610 250852 239822
rect 250812 238604 250864 238610
rect 250812 238546 250864 238552
rect 250824 238474 250852 238546
rect 250812 238468 250864 238474
rect 250812 238410 250864 238416
rect 253124 238134 253152 240094
rect 254734 239850 254762 240108
rect 254688 239822 254762 239850
rect 256712 240094 257324 240122
rect 258092 240094 259256 240122
rect 260852 240094 261188 240122
rect 254688 238513 254716 239822
rect 255228 238808 255280 238814
rect 255228 238750 255280 238756
rect 254674 238504 254730 238513
rect 254674 238439 254730 238448
rect 253112 238128 253164 238134
rect 253112 238070 253164 238076
rect 254688 233102 254716 238439
rect 255240 238406 255268 238750
rect 255228 238400 255280 238406
rect 255228 238342 255280 238348
rect 254676 233096 254728 233102
rect 254676 233038 254728 233044
rect 256712 225622 256740 240094
rect 256700 225616 256752 225622
rect 256700 225558 256752 225564
rect 252744 220244 252796 220250
rect 252744 220186 252796 220192
rect 251180 220176 251232 220182
rect 251180 220118 251232 220124
rect 248420 217388 248472 217394
rect 248420 217330 248472 217336
rect 249800 216028 249852 216034
rect 249800 215970 249852 215976
rect 249064 193928 249116 193934
rect 249064 193870 249116 193876
rect 247776 188488 247828 188494
rect 247776 188430 247828 188436
rect 247788 178974 247816 188430
rect 247776 178968 247828 178974
rect 247776 178910 247828 178916
rect 248052 176656 248104 176662
rect 248052 176598 248104 176604
rect 247682 176080 247738 176089
rect 247682 176015 247738 176024
rect 243544 175840 243596 175846
rect 248064 175817 248092 176598
rect 243544 175782 243596 175788
rect 248050 175808 248106 175817
rect 248050 175743 248106 175752
rect 249076 160562 249104 193870
rect 249340 178968 249392 178974
rect 249340 178910 249392 178916
rect 249248 177472 249300 177478
rect 249248 177414 249300 177420
rect 249156 175840 249208 175846
rect 249156 175782 249208 175788
rect 249168 175273 249196 175782
rect 249154 175264 249210 175273
rect 249154 175199 249210 175208
rect 249260 171873 249288 177414
rect 249352 173369 249380 178910
rect 249432 178900 249484 178906
rect 249432 178842 249484 178848
rect 249338 173360 249394 173369
rect 249338 173295 249394 173304
rect 249444 172825 249472 178842
rect 249430 172816 249486 172825
rect 249430 172751 249486 172760
rect 249246 171864 249302 171873
rect 249246 171799 249302 171808
rect 249154 160576 249210 160585
rect 249076 160534 249154 160562
rect 249154 160511 249210 160520
rect 249812 153513 249840 215970
rect 249892 206508 249944 206514
rect 249892 206450 249944 206456
rect 249798 153504 249854 153513
rect 249798 153439 249854 153448
rect 249904 151201 249932 206450
rect 249984 192704 250036 192710
rect 249984 192646 250036 192652
rect 249996 190454 250024 192646
rect 249996 190426 250208 190454
rect 250180 164393 250208 190426
rect 250166 164384 250222 164393
rect 250166 164319 250222 164328
rect 251192 157865 251220 220118
rect 252652 207800 252704 207806
rect 252652 207742 252704 207748
rect 251272 181552 251324 181558
rect 251272 181494 251324 181500
rect 251178 157856 251234 157865
rect 251178 157791 251234 157800
rect 251180 157140 251232 157146
rect 251180 157082 251232 157088
rect 251192 156369 251220 157082
rect 251178 156360 251234 156369
rect 251178 156295 251234 156304
rect 249890 151192 249946 151201
rect 249890 151127 249946 151136
rect 250628 151088 250680 151094
rect 250628 151030 250680 151036
rect 250640 143177 250668 151030
rect 251180 150204 251232 150210
rect 251180 150146 251232 150152
rect 251192 149841 251220 150146
rect 251178 149832 251234 149841
rect 251178 149767 251234 149776
rect 251284 149297 251312 181494
rect 251364 180192 251416 180198
rect 251364 180134 251416 180140
rect 251376 158817 251404 180134
rect 252560 179036 252612 179042
rect 252560 178978 252612 178984
rect 251456 177404 251508 177410
rect 251456 177346 251508 177352
rect 251468 159225 251496 177346
rect 251822 172408 251878 172417
rect 251822 172343 251878 172352
rect 251836 171902 251864 172343
rect 251824 171896 251876 171902
rect 251824 171838 251876 171844
rect 252572 171465 252600 178978
rect 252558 171456 252614 171465
rect 252558 171391 252614 171400
rect 251732 171080 251784 171086
rect 251732 171022 251784 171028
rect 251744 170921 251772 171022
rect 251730 170912 251786 170921
rect 251730 170847 251786 170856
rect 251822 170504 251878 170513
rect 251822 170439 251878 170448
rect 251836 169862 251864 170439
rect 251824 169856 251876 169862
rect 251824 169798 251876 169804
rect 252468 169652 252520 169658
rect 252468 169594 252520 169600
rect 252480 169153 252508 169594
rect 252466 169144 252522 169153
rect 252466 169079 252522 169088
rect 252376 168360 252428 168366
rect 252376 168302 252428 168308
rect 252388 167249 252416 168302
rect 252468 168224 252520 168230
rect 252466 168192 252468 168201
rect 252520 168192 252522 168201
rect 252466 168127 252522 168136
rect 252466 167648 252522 167657
rect 252466 167583 252522 167592
rect 252480 167278 252508 167583
rect 252468 167272 252520 167278
rect 252374 167240 252430 167249
rect 252468 167214 252520 167220
rect 252374 167175 252430 167184
rect 252468 167000 252520 167006
rect 252468 166942 252520 166948
rect 252376 166864 252428 166870
rect 252376 166806 252428 166812
rect 252388 166705 252416 166806
rect 252374 166696 252430 166705
rect 252374 166631 252430 166640
rect 252284 166320 252336 166326
rect 252480 166297 252508 166942
rect 252284 166262 252336 166268
rect 252466 166288 252522 166297
rect 252296 165753 252324 166262
rect 252466 166223 252522 166232
rect 252282 165744 252338 165753
rect 252282 165679 252338 165688
rect 252468 165572 252520 165578
rect 252468 165514 252520 165520
rect 252480 165345 252508 165514
rect 252466 165336 252522 165345
rect 252466 165271 252522 165280
rect 252468 165028 252520 165034
rect 252468 164970 252520 164976
rect 252480 164801 252508 164970
rect 252466 164792 252522 164801
rect 252466 164727 252522 164736
rect 252192 164212 252244 164218
rect 252192 164154 252244 164160
rect 252204 163033 252232 164154
rect 252190 163024 252246 163033
rect 252190 162959 252246 162968
rect 252100 162852 252152 162858
rect 252100 162794 252152 162800
rect 252112 162489 252140 162794
rect 252468 162784 252520 162790
rect 252468 162726 252520 162732
rect 252098 162480 252154 162489
rect 252098 162415 252154 162424
rect 251548 162104 251600 162110
rect 252480 162081 252508 162726
rect 251548 162046 251600 162052
rect 252466 162072 252522 162081
rect 251560 161537 251588 162046
rect 252466 162007 252522 162016
rect 251546 161528 251602 161537
rect 251546 161463 251602 161472
rect 251548 160268 251600 160274
rect 251548 160210 251600 160216
rect 251560 160177 251588 160210
rect 251546 160168 251602 160177
rect 251546 160103 251602 160112
rect 251454 159216 251510 159225
rect 251454 159151 251510 159160
rect 251362 158808 251418 158817
rect 251362 158743 251418 158752
rect 252468 158704 252520 158710
rect 252468 158646 252520 158652
rect 252480 158273 252508 158646
rect 252466 158264 252522 158273
rect 252466 158199 252522 158208
rect 251914 157992 251970 158001
rect 251914 157927 251970 157936
rect 251364 157072 251416 157078
rect 251364 157014 251416 157020
rect 251376 156913 251404 157014
rect 251362 156904 251418 156913
rect 251362 156839 251418 156848
rect 251824 155916 251876 155922
rect 251824 155858 251876 155864
rect 251836 155009 251864 155858
rect 251822 155000 251878 155009
rect 251822 154935 251878 154944
rect 251928 151814 251956 157927
rect 252374 155952 252430 155961
rect 252374 155887 252430 155896
rect 252388 155786 252416 155887
rect 252468 155848 252520 155854
rect 252468 155790 252520 155796
rect 252376 155780 252428 155786
rect 252376 155722 252428 155728
rect 252480 155417 252508 155790
rect 252466 155408 252522 155417
rect 252466 155343 252522 155352
rect 252284 155304 252336 155310
rect 252284 155246 252336 155252
rect 252100 154352 252152 154358
rect 252100 154294 252152 154300
rect 252112 151814 252140 154294
rect 252296 152153 252324 155246
rect 252468 154556 252520 154562
rect 252468 154498 252520 154504
rect 252480 154057 252508 154498
rect 252664 154465 252692 207742
rect 252756 169561 252784 220186
rect 252836 217456 252888 217462
rect 252836 217398 252888 217404
rect 252742 169552 252798 169561
rect 252742 169487 252798 169496
rect 252848 162110 252876 217398
rect 256700 214804 256752 214810
rect 256700 214746 256752 214752
rect 255412 206440 255464 206446
rect 255412 206382 255464 206388
rect 254032 185768 254084 185774
rect 254032 185710 254084 185716
rect 253940 182980 253992 182986
rect 253940 182922 253992 182928
rect 253202 163976 253258 163985
rect 253202 163911 253258 163920
rect 253216 163033 253244 163911
rect 253202 163024 253258 163033
rect 253202 162959 253258 162968
rect 252836 162104 252888 162110
rect 252836 162046 252888 162052
rect 253296 158772 253348 158778
rect 253296 158714 253348 158720
rect 252650 154456 252706 154465
rect 252650 154391 252706 154400
rect 252466 154048 252522 154057
rect 252466 153983 252522 153992
rect 252376 153196 252428 153202
rect 252376 153138 252428 153144
rect 252388 152697 252416 153138
rect 252468 153128 252520 153134
rect 252466 153096 252468 153105
rect 252520 153096 252522 153105
rect 252466 153031 252522 153040
rect 252374 152688 252430 152697
rect 252374 152623 252430 152632
rect 252282 152144 252338 152153
rect 252282 152079 252338 152088
rect 251836 151786 251956 151814
rect 252020 151786 252140 151814
rect 251270 149288 251326 149297
rect 251270 149223 251326 149232
rect 251836 148889 251864 151786
rect 251916 151700 251968 151706
rect 251916 151642 251968 151648
rect 251928 150793 251956 151642
rect 251914 150784 251970 150793
rect 251914 150719 251970 150728
rect 251822 148880 251878 148889
rect 251822 148815 251878 148824
rect 251732 147484 251784 147490
rect 251732 147426 251784 147432
rect 251548 147008 251600 147014
rect 251744 146985 251772 147426
rect 251548 146950 251600 146956
rect 251730 146976 251786 146985
rect 251560 144673 251588 146950
rect 251730 146911 251786 146920
rect 251916 144900 251968 144906
rect 251916 144842 251968 144848
rect 251546 144664 251602 144673
rect 251546 144599 251602 144608
rect 251928 144129 251956 144842
rect 251914 144120 251970 144129
rect 251914 144055 251970 144064
rect 250626 143168 250682 143177
rect 250626 143103 250682 143112
rect 251824 142860 251876 142866
rect 251824 142802 251876 142808
rect 251086 142624 251142 142633
rect 251086 142559 251142 142568
rect 250536 138032 250588 138038
rect 250536 137974 250588 137980
rect 250444 136672 250496 136678
rect 250444 136614 250496 136620
rect 249156 114572 249208 114578
rect 249156 114514 249208 114520
rect 217968 99340 218020 99346
rect 217968 99282 218020 99288
rect 217980 99226 218008 99282
rect 217980 99198 218100 99226
rect 217324 98728 217376 98734
rect 217324 98670 217376 98676
rect 217336 89690 217364 98670
rect 217416 98660 217468 98666
rect 217416 98602 217468 98608
rect 217428 93838 217456 98602
rect 218072 95985 218100 99198
rect 218058 95976 218114 95985
rect 218058 95911 218114 95920
rect 249064 95260 249116 95266
rect 249064 95202 249116 95208
rect 246304 94512 246356 94518
rect 246304 94454 246356 94460
rect 217416 93832 217468 93838
rect 217416 93774 217468 93780
rect 238024 91928 238076 91934
rect 238024 91870 238076 91876
rect 228364 91860 228416 91866
rect 228364 91802 228416 91808
rect 217324 89684 217376 89690
rect 217324 89626 217376 89632
rect 228376 29714 228404 91802
rect 233884 87644 233936 87650
rect 233884 87586 233936 87592
rect 228364 29708 228416 29714
rect 228364 29650 228416 29656
rect 233896 14550 233924 87586
rect 233884 14544 233936 14550
rect 233884 14486 233936 14492
rect 216680 11892 216732 11898
rect 216680 11834 216732 11840
rect 216128 3732 216180 3738
rect 216128 3674 216180 3680
rect 216036 3596 216088 3602
rect 216036 3538 216088 3544
rect 211896 3528 211948 3534
rect 211896 3470 211948 3476
rect 215944 3528 215996 3534
rect 215944 3470 215996 3476
rect 192484 3460 192536 3466
rect 192484 3402 192536 3408
rect 196624 3460 196676 3466
rect 196624 3402 196676 3408
rect 238036 3398 238064 91870
rect 242900 86284 242952 86290
rect 242900 86226 242952 86232
rect 238760 79416 238812 79422
rect 238760 79358 238812 79364
rect 238772 16574 238800 79358
rect 242164 24268 242216 24274
rect 242164 24210 242216 24216
rect 238772 16546 239352 16574
rect 135260 3392 135312 3398
rect 135260 3334 135312 3340
rect 136456 3392 136508 3398
rect 136456 3334 136508 3340
rect 235816 3392 235868 3398
rect 235816 3334 235868 3340
rect 238024 3392 238076 3398
rect 238024 3334 238076 3340
rect 136468 480 136496 3334
rect 235828 480 235856 3334
rect 239324 480 239352 16546
rect 242176 3738 242204 24210
rect 240508 3732 240560 3738
rect 240508 3674 240560 3680
rect 242164 3732 242216 3738
rect 242164 3674 242216 3680
rect 240520 480 240548 3674
rect 242912 3398 242940 86226
rect 245660 79348 245712 79354
rect 245660 79290 245712 79296
rect 245672 16574 245700 79290
rect 245672 16546 245976 16574
rect 245200 9104 245252 9110
rect 245200 9046 245252 9052
rect 242900 3392 242952 3398
rect 242900 3334 242952 3340
rect 244096 3392 244148 3398
rect 244096 3334 244148 3340
rect 241704 3324 241756 3330
rect 241704 3266 241756 3272
rect 241716 480 241744 3266
rect 242898 3224 242954 3233
rect 242898 3159 242954 3168
rect 242912 480 242940 3159
rect 244108 480 244136 3334
rect 245212 480 245240 9046
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 16546
rect 246316 3330 246344 94454
rect 249076 43518 249104 95202
rect 249168 71058 249196 114514
rect 249246 97064 249302 97073
rect 249246 96999 249302 97008
rect 249156 71052 249208 71058
rect 249156 70994 249208 71000
rect 249260 48278 249288 96999
rect 249248 48272 249300 48278
rect 249248 48214 249300 48220
rect 249064 43512 249116 43518
rect 249064 43454 249116 43460
rect 250456 32502 250484 136614
rect 250548 76566 250576 137974
rect 250994 95704 251050 95713
rect 250994 95639 251050 95648
rect 251008 91934 251036 95639
rect 250996 91928 251048 91934
rect 250996 91870 251048 91876
rect 250536 76560 250588 76566
rect 250536 76502 250588 76508
rect 250444 32496 250496 32502
rect 250444 32438 250496 32444
rect 247592 3732 247644 3738
rect 247592 3674 247644 3680
rect 246304 3324 246356 3330
rect 246304 3266 246356 3272
rect 247604 480 247632 3674
rect 248788 3664 248840 3670
rect 248788 3606 248840 3612
rect 248800 480 248828 3606
rect 251100 3602 251128 142559
rect 251732 140684 251784 140690
rect 251732 140626 251784 140632
rect 251744 139913 251772 140626
rect 251730 139904 251786 139913
rect 251730 139839 251786 139848
rect 251732 139800 251784 139806
rect 251732 139742 251784 139748
rect 251744 139505 251772 139742
rect 251730 139496 251786 139505
rect 251730 139431 251786 139440
rect 251364 138780 251416 138786
rect 251364 138722 251416 138728
rect 251376 138553 251404 138722
rect 251362 138544 251418 138553
rect 251362 138479 251418 138488
rect 251732 136468 251784 136474
rect 251732 136410 251784 136416
rect 251744 135697 251772 136410
rect 251730 135688 251786 135697
rect 251730 135623 251786 135632
rect 251732 133816 251784 133822
rect 251732 133758 251784 133764
rect 251744 132841 251772 133758
rect 251730 132832 251786 132841
rect 251730 132767 251786 132776
rect 251730 129160 251786 129169
rect 251730 129095 251786 129104
rect 251744 128518 251772 129095
rect 251732 128512 251784 128518
rect 251732 128454 251784 128460
rect 251180 125384 251232 125390
rect 251178 125352 251180 125361
rect 251232 125352 251234 125361
rect 251178 125287 251234 125296
rect 251548 121304 251600 121310
rect 251548 121246 251600 121252
rect 251560 120601 251588 121246
rect 251546 120592 251602 120601
rect 251546 120527 251602 120536
rect 251732 119400 251784 119406
rect 251732 119342 251784 119348
rect 251548 114504 251600 114510
rect 251548 114446 251600 114452
rect 251560 114073 251588 114446
rect 251546 114064 251602 114073
rect 251546 113999 251602 114008
rect 251548 113144 251600 113150
rect 251548 113086 251600 113092
rect 251560 112169 251588 113086
rect 251546 112160 251602 112169
rect 251546 112095 251602 112104
rect 251548 107092 251600 107098
rect 251548 107034 251600 107040
rect 251560 107001 251588 107034
rect 251546 106992 251602 107001
rect 251546 106927 251602 106936
rect 251640 106208 251692 106214
rect 251640 106150 251692 106156
rect 251652 106049 251680 106150
rect 251638 106040 251694 106049
rect 251638 105975 251694 105984
rect 251270 104136 251326 104145
rect 251270 104071 251326 104080
rect 251180 99000 251232 99006
rect 251178 98968 251180 98977
rect 251232 98968 251234 98977
rect 251178 98903 251234 98912
rect 251178 96656 251234 96665
rect 251178 96591 251234 96600
rect 251192 11014 251220 96591
rect 251180 11008 251232 11014
rect 251180 10950 251232 10956
rect 251284 6914 251312 104071
rect 251744 103514 251772 119342
rect 251836 117881 251864 142802
rect 252020 142154 252048 151786
rect 252468 151768 252520 151774
rect 252466 151736 252468 151745
rect 252520 151736 252522 151745
rect 252466 151671 252522 151680
rect 253202 149696 253258 149705
rect 253202 149631 253258 149640
rect 252468 149048 252520 149054
rect 252468 148990 252520 148996
rect 252480 148345 252508 148990
rect 252466 148336 252522 148345
rect 252466 148271 252522 148280
rect 252376 147620 252428 147626
rect 252376 147562 252428 147568
rect 252388 146577 252416 147562
rect 252468 147552 252520 147558
rect 252466 147520 252468 147529
rect 252520 147520 252522 147529
rect 252466 147455 252522 147464
rect 252374 146568 252430 146577
rect 252374 146503 252430 146512
rect 252100 146260 252152 146266
rect 252100 146202 252152 146208
rect 252112 146033 252140 146202
rect 252284 146192 252336 146198
rect 252284 146134 252336 146140
rect 252098 146024 252154 146033
rect 252098 145959 252154 145968
rect 252296 145081 252324 146134
rect 252282 145072 252338 145081
rect 252282 145007 252338 145016
rect 252468 144832 252520 144838
rect 252468 144774 252520 144780
rect 252480 143721 252508 144774
rect 252466 143712 252522 143721
rect 252466 143647 252522 143656
rect 252376 143540 252428 143546
rect 252376 143482 252428 143488
rect 252388 142225 252416 143482
rect 252468 143472 252520 143478
rect 252468 143414 252520 143420
rect 252480 142769 252508 143414
rect 252466 142760 252522 142769
rect 252466 142695 252522 142704
rect 251928 142126 252048 142154
rect 252374 142216 252430 142225
rect 252374 142151 252430 142160
rect 251928 131481 251956 142126
rect 252468 142112 252520 142118
rect 252468 142054 252520 142060
rect 252480 141409 252508 142054
rect 252466 141400 252522 141409
rect 252466 141335 252522 141344
rect 252100 140752 252152 140758
rect 252100 140694 252152 140700
rect 252112 140457 252140 140694
rect 252098 140448 252154 140457
rect 252098 140383 252154 140392
rect 252192 140072 252244 140078
rect 252192 140014 252244 140020
rect 252100 137896 252152 137902
rect 252100 137838 252152 137844
rect 252112 137601 252140 137838
rect 252098 137592 252154 137601
rect 252098 137527 252154 137536
rect 252008 137352 252060 137358
rect 252008 137294 252060 137300
rect 251914 131472 251970 131481
rect 251914 131407 251970 131416
rect 252020 122834 252048 137294
rect 252100 136536 252152 136542
rect 252100 136478 252152 136484
rect 252112 136241 252140 136478
rect 252098 136232 252154 136241
rect 252098 136167 252154 136176
rect 252204 130121 252232 140014
rect 252468 137964 252520 137970
rect 252468 137906 252520 137912
rect 252480 137057 252508 137906
rect 252466 137048 252522 137057
rect 252466 136983 252522 136992
rect 252376 136604 252428 136610
rect 252376 136546 252428 136552
rect 252388 135289 252416 136546
rect 252374 135280 252430 135289
rect 252374 135215 252430 135224
rect 252468 135244 252520 135250
rect 252468 135186 252520 135192
rect 252284 135176 252336 135182
rect 252284 135118 252336 135124
rect 252296 134337 252324 135118
rect 252480 134745 252508 135186
rect 252466 134736 252522 134745
rect 252466 134671 252522 134680
rect 252282 134328 252338 134337
rect 252282 134263 252338 134272
rect 252376 133884 252428 133890
rect 252376 133826 252428 133832
rect 252388 133385 252416 133826
rect 252466 133784 252522 133793
rect 252466 133719 252468 133728
rect 252520 133719 252522 133728
rect 252468 133690 252520 133696
rect 252374 133376 252430 133385
rect 252374 133311 252430 133320
rect 252468 132456 252520 132462
rect 252466 132424 252468 132433
rect 252520 132424 252522 132433
rect 252466 132359 252522 132368
rect 252466 131880 252522 131889
rect 252466 131815 252522 131824
rect 252480 131646 252508 131815
rect 252468 131640 252520 131646
rect 252468 131582 252520 131588
rect 252468 131096 252520 131102
rect 252468 131038 252520 131044
rect 252376 131028 252428 131034
rect 252376 130970 252428 130976
rect 252388 130529 252416 130970
rect 252480 130937 252508 131038
rect 252466 130928 252522 130937
rect 252466 130863 252522 130872
rect 252374 130520 252430 130529
rect 252374 130455 252430 130464
rect 252190 130112 252246 130121
rect 252190 130047 252246 130056
rect 252468 129736 252520 129742
rect 252468 129678 252520 129684
rect 252376 129668 252428 129674
rect 252376 129610 252428 129616
rect 252388 128625 252416 129610
rect 252480 129577 252508 129678
rect 252466 129568 252522 129577
rect 252466 129503 252522 129512
rect 252374 128616 252430 128625
rect 252374 128551 252430 128560
rect 252468 128308 252520 128314
rect 252468 128250 252520 128256
rect 252376 128240 252428 128246
rect 252480 128217 252508 128250
rect 252376 128182 252428 128188
rect 252466 128208 252522 128217
rect 252388 127265 252416 128182
rect 252466 128143 252522 128152
rect 252374 127256 252430 127265
rect 252100 127220 252152 127226
rect 252374 127191 252430 127200
rect 252100 127162 252152 127168
rect 251928 122806 252048 122834
rect 251822 117872 251878 117881
rect 251822 117807 251878 117816
rect 251824 116612 251876 116618
rect 251824 116554 251876 116560
rect 251836 113529 251864 116554
rect 251928 115977 251956 122806
rect 252112 119241 252140 127162
rect 252376 126948 252428 126954
rect 252376 126890 252428 126896
rect 252388 125769 252416 126890
rect 252468 126880 252520 126886
rect 252468 126822 252520 126828
rect 252480 126721 252508 126822
rect 252466 126712 252522 126721
rect 252466 126647 252522 126656
rect 252468 126608 252520 126614
rect 252468 126550 252520 126556
rect 252480 126313 252508 126550
rect 252466 126304 252522 126313
rect 252466 126239 252522 126248
rect 252374 125760 252430 125769
rect 252374 125695 252430 125704
rect 252468 125520 252520 125526
rect 252468 125462 252520 125468
rect 252376 125452 252428 125458
rect 252376 125394 252428 125400
rect 252388 124409 252416 125394
rect 252480 124817 252508 125462
rect 252466 124808 252522 124817
rect 252466 124743 252522 124752
rect 252374 124400 252430 124409
rect 252374 124335 252430 124344
rect 252284 124160 252336 124166
rect 252284 124102 252336 124108
rect 252296 123049 252324 124102
rect 252468 124092 252520 124098
rect 252468 124034 252520 124040
rect 252376 124024 252428 124030
rect 252480 124001 252508 124034
rect 252376 123966 252428 123972
rect 252466 123992 252522 124001
rect 252388 123457 252416 123966
rect 252466 123927 252522 123936
rect 252374 123448 252430 123457
rect 252374 123383 252430 123392
rect 252282 123040 252338 123049
rect 252282 122975 252338 122984
rect 252468 122800 252520 122806
rect 252468 122742 252520 122748
rect 252376 122732 252428 122738
rect 252376 122674 252428 122680
rect 252388 122097 252416 122674
rect 252480 122505 252508 122742
rect 252466 122496 252522 122505
rect 252466 122431 252522 122440
rect 252374 122088 252430 122097
rect 252374 122023 252430 122032
rect 252468 121916 252520 121922
rect 252468 121858 252520 121864
rect 252480 121553 252508 121858
rect 252466 121544 252522 121553
rect 252466 121479 252522 121488
rect 252376 121440 252428 121446
rect 252376 121382 252428 121388
rect 252388 120193 252416 121382
rect 252468 121372 252520 121378
rect 252468 121314 252520 121320
rect 252480 121145 252508 121314
rect 252466 121136 252522 121145
rect 252466 121071 252522 121080
rect 252374 120184 252430 120193
rect 252374 120119 252430 120128
rect 252376 120080 252428 120086
rect 252376 120022 252428 120028
rect 252098 119232 252154 119241
rect 252098 119167 252154 119176
rect 252388 118833 252416 120022
rect 252468 120012 252520 120018
rect 252468 119954 252520 119960
rect 252480 119649 252508 119954
rect 252466 119640 252522 119649
rect 252466 119575 252522 119584
rect 252374 118824 252430 118833
rect 252374 118759 252430 118768
rect 252376 118652 252428 118658
rect 252376 118594 252428 118600
rect 252100 117972 252152 117978
rect 252100 117914 252152 117920
rect 252008 116408 252060 116414
rect 252006 116376 252008 116385
rect 252060 116376 252062 116385
rect 252006 116311 252062 116320
rect 251914 115968 251970 115977
rect 251914 115903 251970 115912
rect 252008 115932 252060 115938
rect 252008 115874 252060 115880
rect 252020 115025 252048 115874
rect 252006 115016 252062 115025
rect 252006 114951 252062 114960
rect 251822 113520 251878 113529
rect 251822 113455 251878 113464
rect 252112 113174 252140 117914
rect 252388 117337 252416 118594
rect 252468 118584 252520 118590
rect 252468 118526 252520 118532
rect 252480 118289 252508 118526
rect 252466 118280 252522 118289
rect 252466 118215 252522 118224
rect 252374 117328 252430 117337
rect 252374 117263 252430 117272
rect 252468 117292 252520 117298
rect 252468 117234 252520 117240
rect 252480 116929 252508 117234
rect 252466 116920 252522 116929
rect 252466 116855 252522 116864
rect 252284 115864 252336 115870
rect 252284 115806 252336 115812
rect 252296 115433 252324 115806
rect 252282 115424 252338 115433
rect 252282 115359 252338 115368
rect 252466 114472 252522 114481
rect 252466 114407 252468 114416
rect 252520 114407 252522 114416
rect 252468 114378 252520 114384
rect 252192 114368 252244 114374
rect 252192 114310 252244 114316
rect 252020 113146 252140 113174
rect 252020 105754 252048 113146
rect 252100 110016 252152 110022
rect 252100 109958 252152 109964
rect 252112 109857 252140 109958
rect 252098 109848 252154 109857
rect 252098 109783 252154 109792
rect 252100 108724 252152 108730
rect 252100 108666 252152 108672
rect 252112 107953 252140 108666
rect 252098 107944 252154 107953
rect 252098 107879 252154 107888
rect 252100 106276 252152 106282
rect 252100 106218 252152 106224
rect 251836 105726 252048 105754
rect 251836 104689 251864 105726
rect 252008 105596 252060 105602
rect 252008 105538 252060 105544
rect 251822 104680 251878 104689
rect 251822 104615 251878 104624
rect 251744 103486 251956 103514
rect 251928 102785 251956 103486
rect 251914 102776 251970 102785
rect 251914 102711 251970 102720
rect 251824 102060 251876 102066
rect 251824 102002 251876 102008
rect 251836 101425 251864 102002
rect 251822 101416 251878 101425
rect 251822 101351 251878 101360
rect 251916 100700 251968 100706
rect 251916 100642 251968 100648
rect 251928 99929 251956 100642
rect 252020 100473 252048 105538
rect 252112 105097 252140 106218
rect 252098 105088 252154 105097
rect 252098 105023 252154 105032
rect 252100 104848 252152 104854
rect 252100 104790 252152 104796
rect 252112 103737 252140 104790
rect 252098 103728 252154 103737
rect 252098 103663 252154 103672
rect 252204 103193 252232 114310
rect 252374 113112 252430 113121
rect 252374 113047 252430 113056
rect 252468 113076 252520 113082
rect 252388 112266 252416 113047
rect 252468 113018 252520 113024
rect 252480 112713 252508 113018
rect 252466 112704 252522 112713
rect 252466 112639 252522 112648
rect 252376 112260 252428 112266
rect 252376 112202 252428 112208
rect 252468 111784 252520 111790
rect 252374 111752 252430 111761
rect 252468 111726 252520 111732
rect 252374 111687 252376 111696
rect 252428 111687 252430 111696
rect 252376 111658 252428 111664
rect 252480 110809 252508 111726
rect 252466 110800 252522 110809
rect 252466 110735 252522 110744
rect 252376 110424 252428 110430
rect 252376 110366 252428 110372
rect 252388 109313 252416 110366
rect 252468 110356 252520 110362
rect 252468 110298 252520 110304
rect 252480 110265 252508 110298
rect 252466 110256 252522 110265
rect 252466 110191 252522 110200
rect 252374 109304 252430 109313
rect 252374 109239 252430 109248
rect 252468 108996 252520 109002
rect 252468 108938 252520 108944
rect 252376 108928 252428 108934
rect 252480 108905 252508 108938
rect 252376 108870 252428 108876
rect 252466 108896 252522 108905
rect 252388 108361 252416 108870
rect 252466 108831 252522 108840
rect 252374 108352 252430 108361
rect 252374 108287 252430 108296
rect 252468 107636 252520 107642
rect 252468 107578 252520 107584
rect 252376 107568 252428 107574
rect 252480 107545 252508 107578
rect 252376 107510 252428 107516
rect 252466 107536 252522 107545
rect 252388 106593 252416 107510
rect 252466 107471 252522 107480
rect 252468 106956 252520 106962
rect 252468 106898 252520 106904
rect 252374 106584 252430 106593
rect 252374 106519 252430 106528
rect 252480 105641 252508 106898
rect 252466 105632 252522 105641
rect 252466 105567 252522 105576
rect 252284 104440 252336 104446
rect 252284 104382 252336 104388
rect 252296 104281 252324 104382
rect 252282 104272 252338 104281
rect 252282 104207 252338 104216
rect 252468 103488 252520 103494
rect 252468 103430 252520 103436
rect 252190 103184 252246 103193
rect 252190 103119 252246 103128
rect 252376 102808 252428 102814
rect 252376 102750 252428 102756
rect 252100 102128 252152 102134
rect 252100 102070 252152 102076
rect 252112 100881 252140 102070
rect 252388 101833 252416 102750
rect 252480 102241 252508 103430
rect 252466 102232 252522 102241
rect 252466 102167 252522 102176
rect 252374 101824 252430 101833
rect 252374 101759 252430 101768
rect 252466 101416 252522 101425
rect 252466 101351 252522 101360
rect 252098 100872 252154 100881
rect 252098 100807 252154 100816
rect 252100 100632 252152 100638
rect 252100 100574 252152 100580
rect 252006 100464 252062 100473
rect 252006 100399 252062 100408
rect 251914 99920 251970 99929
rect 251914 99855 251970 99864
rect 252112 99521 252140 100574
rect 252284 100020 252336 100026
rect 252284 99962 252336 99968
rect 252098 99512 252154 99521
rect 252098 99447 252154 99456
rect 251916 98660 251968 98666
rect 251916 98602 251968 98608
rect 251822 97880 251878 97889
rect 251822 97815 251878 97824
rect 251836 97073 251864 97815
rect 251928 97617 251956 98602
rect 252296 98025 252324 99962
rect 252376 99272 252428 99278
rect 252376 99214 252428 99220
rect 252388 98569 252416 99214
rect 252374 98560 252430 98569
rect 252374 98495 252430 98504
rect 252282 98016 252338 98025
rect 252282 97951 252338 97960
rect 251914 97608 251970 97617
rect 251914 97543 251970 97552
rect 251822 97064 251878 97073
rect 251822 96999 251878 97008
rect 252480 96665 252508 101351
rect 253216 99006 253244 149631
rect 253308 127226 253336 158714
rect 253952 150210 253980 182922
rect 254044 157146 254072 185710
rect 254124 178696 254176 178702
rect 254124 178638 254176 178644
rect 254032 157140 254084 157146
rect 254032 157082 254084 157088
rect 254136 157078 254164 178638
rect 254214 177304 254270 177313
rect 254214 177239 254270 177248
rect 254228 160274 254256 177239
rect 255320 176588 255372 176594
rect 255320 176530 255372 176536
rect 255332 176497 255360 176530
rect 255318 176488 255374 176497
rect 255318 176423 255374 176432
rect 254216 160268 254268 160274
rect 254216 160210 254268 160216
rect 254124 157072 254176 157078
rect 254124 157014 254176 157020
rect 255424 153066 255452 206382
rect 255596 202224 255648 202230
rect 255596 202166 255648 202172
rect 255504 199640 255556 199646
rect 255504 199582 255556 199588
rect 254584 153060 254636 153066
rect 254584 153002 254636 153008
rect 255412 153060 255464 153066
rect 255412 153002 255464 153008
rect 254124 151836 254176 151842
rect 254124 151778 254176 151784
rect 253940 150204 253992 150210
rect 253940 150146 253992 150152
rect 254136 146305 254164 151778
rect 254122 146296 254178 146305
rect 254122 146231 254178 146240
rect 253480 141432 253532 141438
rect 253480 141374 253532 141380
rect 253388 139460 253440 139466
rect 253388 139402 253440 139408
rect 253296 127220 253348 127226
rect 253296 127162 253348 127168
rect 253204 99000 253256 99006
rect 253204 98942 253256 98948
rect 253296 96688 253348 96694
rect 252466 96656 252522 96665
rect 253296 96630 253348 96636
rect 252466 96591 252522 96600
rect 253204 86352 253256 86358
rect 253204 86294 253256 86300
rect 251192 6886 251312 6914
rect 251088 3596 251140 3602
rect 251088 3538 251140 3544
rect 249984 3392 250036 3398
rect 249984 3334 250036 3340
rect 249996 480 250024 3334
rect 251192 480 251220 6886
rect 252376 3596 252428 3602
rect 252376 3538 252428 3544
rect 252388 480 252416 3538
rect 253216 3398 253244 86294
rect 253308 18630 253336 96630
rect 253400 69766 253428 139402
rect 253492 125390 253520 141374
rect 254596 138786 254624 153002
rect 254676 147688 254728 147694
rect 254676 147630 254728 147636
rect 254584 138780 254636 138786
rect 254584 138722 254636 138728
rect 253480 125384 253532 125390
rect 253480 125326 253532 125332
rect 254584 113280 254636 113286
rect 254584 113222 254636 113228
rect 253388 69760 253440 69766
rect 253388 69702 253440 69708
rect 253296 18624 253348 18630
rect 253296 18566 253348 18572
rect 254596 13190 254624 113222
rect 254688 107098 254716 147630
rect 255516 147490 255544 199582
rect 255504 147484 255556 147490
rect 255504 147426 255556 147432
rect 254860 145104 254912 145110
rect 254860 145046 254912 145052
rect 254768 144220 254820 144226
rect 254768 144162 254820 144168
rect 254676 107092 254728 107098
rect 254676 107034 254728 107040
rect 254780 106214 254808 144162
rect 254872 114374 254900 145046
rect 255608 139806 255636 202166
rect 256712 171086 256740 214746
rect 256792 180464 256844 180470
rect 256792 180406 256844 180412
rect 256700 171080 256752 171086
rect 256700 171022 256752 171028
rect 256804 166870 256832 180406
rect 258092 179194 258120 240094
rect 259552 211880 259604 211886
rect 259552 211822 259604 211828
rect 259460 207868 259512 207874
rect 259460 207810 259512 207816
rect 258172 194064 258224 194070
rect 258172 194006 258224 194012
rect 258184 180690 258212 194006
rect 258184 180662 258304 180690
rect 258092 179166 258212 179194
rect 258080 178764 258132 178770
rect 258080 178706 258132 178712
rect 256976 177540 257028 177546
rect 256976 177482 257028 177488
rect 256988 168230 257016 177482
rect 258092 171902 258120 178706
rect 258184 177818 258212 179166
rect 258172 177812 258224 177818
rect 258172 177754 258224 177760
rect 258276 177698 258304 180662
rect 258356 180396 258408 180402
rect 258356 180338 258408 180344
rect 258184 177670 258304 177698
rect 258080 171896 258132 171902
rect 258080 171838 258132 171844
rect 257344 169788 257396 169794
rect 257344 169730 257396 169736
rect 256976 168224 257028 168230
rect 256976 168166 257028 168172
rect 256792 166864 256844 166870
rect 256792 166806 256844 166812
rect 257356 154358 257384 169730
rect 258184 167278 258212 177670
rect 258264 177608 258316 177614
rect 258264 177550 258316 177556
rect 258172 167272 258224 167278
rect 258172 167214 258224 167220
rect 258276 167006 258304 177550
rect 258264 167000 258316 167006
rect 258264 166942 258316 166948
rect 257528 165640 257580 165646
rect 257528 165582 257580 165588
rect 257436 160132 257488 160138
rect 257436 160074 257488 160080
rect 257344 154352 257396 154358
rect 257344 154294 257396 154300
rect 256240 152516 256292 152522
rect 256240 152458 256292 152464
rect 256056 150476 256108 150482
rect 256056 150418 256108 150424
rect 255964 145036 256016 145042
rect 255964 144978 256016 144984
rect 255596 139800 255648 139806
rect 255596 139742 255648 139748
rect 254860 114368 254912 114374
rect 254860 114310 254912 114316
rect 254768 106208 254820 106214
rect 254768 106150 254820 106156
rect 255976 104446 256004 144978
rect 256068 110022 256096 150418
rect 256148 146940 256200 146946
rect 256148 146882 256200 146888
rect 256056 110016 256108 110022
rect 256056 109958 256108 109964
rect 256160 108730 256188 146882
rect 256252 146305 256280 152458
rect 257344 151904 257396 151910
rect 257344 151846 257396 151852
rect 256238 146296 256294 146305
rect 256238 146231 256294 146240
rect 257356 111722 257384 151846
rect 257448 121310 257476 160074
rect 257540 126614 257568 165582
rect 257620 155984 257672 155990
rect 257620 155926 257672 155932
rect 257528 126608 257580 126614
rect 257528 126550 257580 126556
rect 257436 121304 257488 121310
rect 257436 121246 257488 121252
rect 257632 116414 257660 155926
rect 258368 146198 258396 180338
rect 258908 168428 258960 168434
rect 258908 168370 258960 168376
rect 258816 157412 258868 157418
rect 258816 157354 258868 157360
rect 258724 153264 258776 153270
rect 258724 153206 258776 153212
rect 258356 146192 258408 146198
rect 258356 146134 258408 146140
rect 257712 126268 257764 126274
rect 257712 126210 257764 126216
rect 257620 116408 257672 116414
rect 257620 116350 257672 116356
rect 257344 111716 257396 111722
rect 257344 111658 257396 111664
rect 256148 108724 256200 108730
rect 256148 108666 256200 108672
rect 256056 106480 256108 106486
rect 256056 106422 256108 106428
rect 255964 104440 256016 104446
rect 255964 104382 256016 104388
rect 255964 98048 256016 98054
rect 255964 97990 256016 97996
rect 255976 22778 256004 97990
rect 256068 33862 256096 106422
rect 257724 94518 257752 126210
rect 258736 112266 258764 153206
rect 258828 118590 258856 157354
rect 258920 128518 258948 168370
rect 259472 151094 259500 207810
rect 259564 166326 259592 211822
rect 259644 189780 259696 189786
rect 259644 189722 259696 189728
rect 259656 169862 259684 189722
rect 259736 175976 259788 175982
rect 259736 175918 259788 175924
rect 259644 169856 259696 169862
rect 259644 169798 259696 169804
rect 259552 166320 259604 166326
rect 259552 166262 259604 166268
rect 259748 165034 259776 175918
rect 259736 165028 259788 165034
rect 259736 164970 259788 164976
rect 260380 163532 260432 163538
rect 260380 163474 260432 163480
rect 260104 161492 260156 161498
rect 260104 161434 260156 161440
rect 259460 151088 259512 151094
rect 259460 151030 259512 151036
rect 258908 128512 258960 128518
rect 258908 128454 258960 128460
rect 260116 121922 260144 161434
rect 260288 154624 260340 154630
rect 260288 154566 260340 154572
rect 260196 149116 260248 149122
rect 260196 149058 260248 149064
rect 260104 121916 260156 121922
rect 260104 121858 260156 121864
rect 258816 118584 258868 118590
rect 258816 118526 258868 118532
rect 260104 113824 260156 113830
rect 260104 113766 260156 113772
rect 258724 112260 258776 112266
rect 258724 112202 258776 112208
rect 258724 110492 258776 110498
rect 258724 110434 258776 110440
rect 257712 94512 257764 94518
rect 257712 94454 257764 94460
rect 257988 78056 258040 78062
rect 257988 77998 258040 78004
rect 256056 33856 256108 33862
rect 256056 33798 256108 33804
rect 255964 22772 256016 22778
rect 255964 22714 256016 22720
rect 254584 13184 254636 13190
rect 254584 13126 254636 13132
rect 253480 3732 253532 3738
rect 253480 3674 253532 3680
rect 253204 3392 253256 3398
rect 253204 3334 253256 3340
rect 253492 480 253520 3674
rect 254676 3664 254728 3670
rect 254676 3606 254728 3612
rect 254688 480 254716 3606
rect 258000 3602 258028 77998
rect 258736 39438 258764 110434
rect 258816 107908 258868 107914
rect 258816 107850 258868 107856
rect 258828 50454 258856 107850
rect 258816 50448 258868 50454
rect 258816 50390 258868 50396
rect 258816 43648 258868 43654
rect 258816 43590 258868 43596
rect 258724 39432 258776 39438
rect 258724 39374 258776 39380
rect 257988 3596 258040 3602
rect 257988 3538 258040 3544
rect 258828 3534 258856 43590
rect 259458 6352 259514 6361
rect 259458 6287 259514 6296
rect 258816 3528 258868 3534
rect 255870 3496 255926 3505
rect 255870 3431 255926 3440
rect 257066 3496 257122 3505
rect 258816 3470 258868 3476
rect 257066 3431 257122 3440
rect 255884 480 255912 3431
rect 257080 480 257108 3431
rect 258264 3052 258316 3058
rect 258264 2994 258316 3000
rect 258276 480 258304 2994
rect 259472 480 259500 6287
rect 260116 3058 260144 113766
rect 260208 108934 260236 149058
rect 260300 114442 260328 154566
rect 260392 131646 260420 163474
rect 260852 162178 260880 240094
rect 263106 239850 263134 240108
rect 265682 239850 265710 240108
rect 263060 239822 263134 239850
rect 265636 239822 265710 239850
rect 266372 240094 267628 240122
rect 269560 240094 269896 240122
rect 263060 238406 263088 239822
rect 263048 238400 263100 238406
rect 263048 238342 263100 238348
rect 263060 234598 263088 238342
rect 263600 238128 263652 238134
rect 263600 238070 263652 238076
rect 263048 234592 263100 234598
rect 263048 234534 263100 234540
rect 263612 222086 263640 238070
rect 265636 235618 265664 239822
rect 265624 235612 265676 235618
rect 265624 235554 265676 235560
rect 265636 228993 265664 235554
rect 265622 228984 265678 228993
rect 265622 228919 265678 228928
rect 265636 227769 265664 228919
rect 265622 227760 265678 227769
rect 265622 227695 265678 227704
rect 263600 222080 263652 222086
rect 263600 222022 263652 222028
rect 264244 222080 264296 222086
rect 264244 222022 264296 222028
rect 261484 216164 261536 216170
rect 261484 216106 261536 216112
rect 261496 198286 261524 216106
rect 263600 214736 263652 214742
rect 263600 214678 263652 214684
rect 262312 200932 262364 200938
rect 262312 200874 262364 200880
rect 261484 198280 261536 198286
rect 261484 198222 261536 198228
rect 260932 198212 260984 198218
rect 260932 198154 260984 198160
rect 260840 162172 260892 162178
rect 260840 162114 260892 162120
rect 260944 142118 260972 198154
rect 261024 195424 261076 195430
rect 261024 195366 261076 195372
rect 261036 169658 261064 195366
rect 262220 188420 262272 188426
rect 262220 188362 262272 188368
rect 261668 172576 261720 172582
rect 261668 172518 261720 172524
rect 261024 169652 261076 169658
rect 261024 169594 261076 169600
rect 261484 162920 261536 162926
rect 261484 162862 261536 162868
rect 260932 142112 260984 142118
rect 260932 142054 260984 142060
rect 260380 131640 260432 131646
rect 260380 131582 260432 131588
rect 260380 124432 260432 124438
rect 260380 124374 260432 124380
rect 260288 114436 260340 114442
rect 260288 114378 260340 114384
rect 260196 108928 260248 108934
rect 260196 108870 260248 108876
rect 260392 91866 260420 124374
rect 261496 124030 261524 162862
rect 261576 158840 261628 158846
rect 261576 158782 261628 158788
rect 261484 124024 261536 124030
rect 261484 123966 261536 123972
rect 261588 120018 261616 158782
rect 261680 133754 261708 172518
rect 262232 144838 262260 188362
rect 262324 164218 262352 200874
rect 262404 196920 262456 196926
rect 262404 196862 262456 196868
rect 262416 168366 262444 196862
rect 262864 171148 262916 171154
rect 262864 171090 262916 171096
rect 262404 168360 262456 168366
rect 262404 168302 262456 168308
rect 262312 164212 262364 164218
rect 262312 164154 262364 164160
rect 262220 144832 262272 144838
rect 262220 144774 262272 144780
rect 262876 133822 262904 171090
rect 262956 167068 263008 167074
rect 262956 167010 263008 167016
rect 262968 148209 262996 167010
rect 263140 160200 263192 160206
rect 263140 160142 263192 160148
rect 262954 148200 263010 148209
rect 262954 148135 263010 148144
rect 263048 146328 263100 146334
rect 263048 146270 263100 146276
rect 262864 133816 262916 133822
rect 262864 133758 262916 133764
rect 261668 133748 261720 133754
rect 261668 133690 261720 133696
rect 261760 133204 261812 133210
rect 261760 133146 261812 133152
rect 261576 120012 261628 120018
rect 261576 119954 261628 119960
rect 261576 116000 261628 116006
rect 261576 115942 261628 115948
rect 261484 95940 261536 95946
rect 261484 95882 261536 95888
rect 260380 91860 260432 91866
rect 260380 91802 260432 91808
rect 260656 4888 260708 4894
rect 260656 4830 260708 4836
rect 260104 3052 260156 3058
rect 260104 2994 260156 3000
rect 260668 480 260696 4830
rect 261496 3738 261524 95882
rect 261588 51746 261616 115942
rect 261772 100638 261800 133146
rect 262864 131164 262916 131170
rect 262864 131106 262916 131112
rect 261760 100632 261812 100638
rect 261760 100574 261812 100580
rect 261576 51740 261628 51746
rect 261576 51682 261628 51688
rect 262220 29776 262272 29782
rect 262220 29718 262272 29724
rect 262232 16574 262260 29718
rect 262876 24206 262904 131106
rect 262956 120148 263008 120154
rect 262956 120090 263008 120096
rect 262864 24200 262916 24206
rect 262864 24142 262916 24148
rect 262232 16546 262536 16574
rect 261484 3732 261536 3738
rect 261484 3674 261536 3680
rect 261760 3528 261812 3534
rect 261760 3470 261812 3476
rect 261772 480 261800 3470
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16546
rect 262968 15910 262996 120090
rect 263060 106962 263088 146270
rect 263152 121378 263180 160142
rect 263612 155786 263640 214678
rect 263692 180328 263744 180334
rect 263692 180270 263744 180276
rect 263704 162790 263732 180270
rect 264256 177410 264284 222022
rect 265072 206576 265124 206582
rect 265072 206518 265124 206524
rect 264980 202292 265032 202298
rect 264980 202234 265032 202240
rect 264244 177404 264296 177410
rect 264244 177346 264296 177352
rect 264244 173936 264296 173942
rect 264244 173878 264296 173884
rect 263692 162784 263744 162790
rect 263692 162726 263744 162732
rect 263600 155780 263652 155786
rect 263600 155722 263652 155728
rect 264256 136474 264284 173878
rect 264992 165578 265020 202234
rect 264980 165572 265032 165578
rect 264980 165514 265032 165520
rect 264428 164892 264480 164898
rect 264428 164834 264480 164840
rect 264336 153332 264388 153338
rect 264336 153274 264388 153280
rect 264244 136468 264296 136474
rect 264244 136410 264296 136416
rect 263140 121372 263192 121378
rect 263140 121314 263192 121320
rect 264348 116618 264376 153274
rect 264440 129674 264468 164834
rect 264980 155236 265032 155242
rect 264980 155178 265032 155184
rect 264520 137284 264572 137290
rect 264520 137226 264572 137232
rect 264428 129668 264480 129674
rect 264428 129610 264480 129616
rect 264336 116612 264388 116618
rect 264336 116554 264388 116560
rect 264244 107772 264296 107778
rect 264244 107714 264296 107720
rect 263048 106956 263100 106962
rect 263048 106898 263100 106904
rect 264256 68406 264284 107714
rect 264532 103494 264560 137226
rect 264520 103488 264572 103494
rect 264520 103430 264572 103436
rect 264244 68400 264296 68406
rect 264244 68342 264296 68348
rect 262956 15904 263008 15910
rect 262956 15846 263008 15852
rect 264152 3596 264204 3602
rect 264152 3538 264204 3544
rect 264164 480 264192 3538
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 264992 354 265020 155178
rect 265084 147014 265112 206518
rect 265164 178832 265216 178838
rect 265164 178774 265216 178780
rect 265176 162858 265204 178774
rect 265624 169856 265676 169862
rect 265624 169798 265676 169804
rect 265164 162852 265216 162858
rect 265164 162794 265216 162800
rect 265072 147008 265124 147014
rect 265072 146950 265124 146956
rect 265636 131034 265664 169798
rect 265716 157480 265768 157486
rect 265716 157422 265768 157428
rect 265728 142866 265756 157422
rect 265716 142860 265768 142866
rect 265716 142802 265768 142808
rect 265624 131028 265676 131034
rect 265624 130970 265676 130976
rect 265716 129804 265768 129810
rect 265716 129746 265768 129752
rect 265624 128376 265676 128382
rect 265624 128318 265676 128324
rect 265636 4826 265664 128318
rect 265728 75206 265756 129746
rect 266372 86358 266400 240094
rect 269868 237114 269896 240094
rect 270512 240094 271492 240122
rect 269856 237108 269908 237114
rect 269856 237050 269908 237056
rect 269868 230246 269896 237050
rect 269856 230240 269908 230246
rect 269856 230182 269908 230188
rect 269764 227112 269816 227118
rect 269764 227054 269816 227060
rect 268384 225616 268436 225622
rect 268384 225558 268436 225564
rect 267740 207732 267792 207738
rect 267740 207674 267792 207680
rect 266544 184408 266596 184414
rect 266544 184350 266596 184356
rect 266452 181688 266504 181694
rect 266452 181630 266504 181636
rect 266464 151706 266492 181630
rect 266556 155310 266584 184350
rect 267004 156052 267056 156058
rect 267004 155994 267056 156000
rect 266544 155304 266596 155310
rect 266544 155246 266596 155252
rect 266452 151700 266504 151706
rect 266452 151642 266504 151648
rect 267016 137358 267044 155994
rect 267752 155854 267780 207674
rect 267740 155848 267792 155854
rect 267740 155790 267792 155796
rect 267096 142180 267148 142186
rect 267096 142122 267148 142128
rect 267004 137352 267056 137358
rect 267004 137294 267056 137300
rect 267004 121508 267056 121514
rect 267004 121450 267056 121456
rect 266360 86352 266412 86358
rect 266360 86294 266412 86300
rect 265716 75200 265768 75206
rect 265716 75142 265768 75148
rect 267016 38010 267044 121450
rect 267108 102066 267136 142122
rect 267096 102060 267148 102066
rect 267096 102002 267148 102008
rect 267740 84856 267792 84862
rect 267740 84798 267792 84804
rect 267004 38004 267056 38010
rect 267004 37946 267056 37952
rect 265624 4820 265676 4826
rect 265624 4762 265676 4768
rect 266544 3392 266596 3398
rect 266544 3334 266596 3340
rect 266556 480 266584 3334
rect 267752 480 267780 84798
rect 268396 3670 268424 225558
rect 269304 209160 269356 209166
rect 269304 209102 269356 209108
rect 269212 200864 269264 200870
rect 269212 200806 269264 200812
rect 269120 177472 269172 177478
rect 269120 177414 269172 177420
rect 268476 171216 268528 171222
rect 268476 171158 268528 171164
rect 268488 132462 268516 171158
rect 268568 165708 268620 165714
rect 268568 165650 268620 165656
rect 268476 132456 268528 132462
rect 268476 132398 268528 132404
rect 268580 128246 268608 165650
rect 268568 128240 268620 128246
rect 268568 128182 268620 128188
rect 268476 125656 268528 125662
rect 268476 125598 268528 125604
rect 268488 40730 268516 125598
rect 268476 40724 268528 40730
rect 268476 40666 268528 40672
rect 269132 16574 269160 177414
rect 269224 143478 269252 200806
rect 269316 154562 269344 209102
rect 269776 198218 269804 227054
rect 270512 218006 270540 240094
rect 274054 239850 274082 240108
rect 274008 239822 274082 239850
rect 274008 238610 274036 239822
rect 276124 238754 276152 240502
rect 277932 240094 278084 240122
rect 276032 238726 276152 238754
rect 273996 238604 274048 238610
rect 273996 238546 274048 238552
rect 273904 238060 273956 238066
rect 273904 238002 273956 238008
rect 273260 236700 273312 236706
rect 273260 236642 273312 236648
rect 273272 233102 273300 236642
rect 273260 233096 273312 233102
rect 273260 233038 273312 233044
rect 271880 225684 271932 225690
rect 271880 225626 271932 225632
rect 270500 218000 270552 218006
rect 270500 217942 270552 217948
rect 270512 216714 270540 217942
rect 270500 216708 270552 216714
rect 270500 216650 270552 216656
rect 271236 216708 271288 216714
rect 271236 216650 271288 216656
rect 270500 213308 270552 213314
rect 270500 213250 270552 213256
rect 269764 198212 269816 198218
rect 269764 198154 269816 198160
rect 269764 172644 269816 172650
rect 269764 172586 269816 172592
rect 269304 154556 269356 154562
rect 269304 154498 269356 154504
rect 269212 143472 269264 143478
rect 269212 143414 269264 143420
rect 269776 135182 269804 172586
rect 270512 153134 270540 213250
rect 270592 194132 270644 194138
rect 270592 194074 270644 194080
rect 270500 153128 270552 153134
rect 270500 153070 270552 153076
rect 269856 147756 269908 147762
rect 269856 147698 269908 147704
rect 269764 135176 269816 135182
rect 269764 135118 269816 135124
rect 269764 127016 269816 127022
rect 269764 126958 269816 126964
rect 269132 16546 269712 16574
rect 268844 6384 268896 6390
rect 268844 6326 268896 6332
rect 268384 3664 268436 3670
rect 268384 3606 268436 3612
rect 268856 480 268884 6326
rect 269684 1986 269712 16546
rect 269776 2106 269804 126958
rect 269868 107574 269896 147698
rect 270604 144906 270632 194074
rect 271144 183048 271196 183054
rect 271144 182990 271196 182996
rect 270592 144900 270644 144906
rect 270592 144842 270644 144848
rect 269856 107568 269908 107574
rect 269856 107510 269908 107516
rect 269856 102196 269908 102202
rect 269856 102138 269908 102144
rect 269868 21486 269896 102138
rect 269856 21480 269908 21486
rect 269856 21422 269908 21428
rect 271156 3534 271184 182990
rect 271248 181558 271276 216650
rect 271236 181552 271288 181558
rect 271236 181494 271288 181500
rect 271236 167680 271288 167686
rect 271236 167622 271288 167628
rect 271248 129742 271276 167622
rect 271420 138712 271472 138718
rect 271420 138654 271472 138660
rect 271328 133952 271380 133958
rect 271328 133894 271380 133900
rect 271236 129736 271288 129742
rect 271236 129678 271288 129684
rect 271236 100768 271288 100774
rect 271236 100710 271288 100716
rect 271248 11762 271276 100710
rect 271340 57322 271368 133894
rect 271432 114510 271460 138654
rect 271420 114504 271472 114510
rect 271420 114446 271472 114452
rect 271420 106412 271472 106418
rect 271420 106354 271472 106360
rect 271328 57316 271380 57322
rect 271328 57258 271380 57264
rect 271432 42090 271460 106354
rect 271420 42084 271472 42090
rect 271420 42026 271472 42032
rect 271892 16574 271920 225626
rect 273260 211948 273312 211954
rect 273260 211890 273312 211896
rect 271972 192840 272024 192846
rect 271972 192782 272024 192788
rect 271984 137902 272012 192782
rect 272064 180260 272116 180266
rect 272064 180202 272116 180208
rect 272076 153202 272104 180202
rect 272064 153196 272116 153202
rect 272064 153138 272116 153144
rect 273272 151774 273300 211890
rect 273352 196852 273404 196858
rect 273352 196794 273404 196800
rect 273260 151768 273312 151774
rect 273260 151710 273312 151716
rect 272616 147824 272668 147830
rect 272616 147766 272668 147772
rect 271972 137896 272024 137902
rect 271972 137838 272024 137844
rect 272524 113280 272576 113286
rect 272524 113222 272576 113228
rect 272536 35290 272564 113222
rect 272628 107642 272656 147766
rect 273364 140690 273392 196794
rect 273916 191282 273944 238002
rect 274008 235686 274036 238546
rect 273996 235680 274048 235686
rect 273996 235622 274048 235628
rect 273996 234048 274048 234054
rect 273996 233990 274048 233996
rect 274008 213246 274036 233990
rect 275284 232552 275336 232558
rect 275284 232494 275336 232500
rect 274640 218816 274692 218822
rect 274640 218758 274692 218764
rect 273996 213240 274048 213246
rect 273996 213182 274048 213188
rect 273904 191276 273956 191282
rect 273904 191218 273956 191224
rect 273444 189984 273496 189990
rect 273444 189926 273496 189932
rect 273456 158710 273484 189926
rect 274088 174004 274140 174010
rect 274088 173946 274140 173952
rect 273444 158704 273496 158710
rect 273444 158646 273496 158652
rect 273996 151972 274048 151978
rect 273996 151914 274048 151920
rect 273352 140684 273404 140690
rect 273352 140626 273404 140632
rect 273904 135516 273956 135522
rect 273904 135458 273956 135464
rect 272616 107636 272668 107642
rect 272616 107578 272668 107584
rect 272524 35284 272576 35290
rect 272524 35226 272576 35232
rect 273260 20120 273312 20126
rect 273260 20062 273312 20068
rect 271892 16546 272472 16574
rect 271236 11756 271288 11762
rect 271236 11698 271288 11704
rect 271144 3528 271196 3534
rect 271144 3470 271196 3476
rect 271234 3496 271290 3505
rect 271234 3431 271290 3440
rect 269764 2100 269816 2106
rect 269764 2042 269816 2048
rect 269684 1958 270080 1986
rect 270052 480 270080 1958
rect 271248 480 271276 3431
rect 272444 480 272472 16546
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273272 354 273300 20062
rect 273916 7682 273944 135458
rect 274008 111790 274036 151914
rect 274100 136542 274128 173946
rect 274652 146266 274680 218758
rect 274732 188352 274784 188358
rect 274732 188294 274784 188300
rect 274640 146260 274692 146266
rect 274640 146202 274692 146208
rect 274640 144288 274692 144294
rect 274640 144230 274692 144236
rect 274088 136536 274140 136542
rect 274088 136478 274140 136484
rect 273996 111784 274048 111790
rect 273996 111726 274048 111732
rect 274088 110560 274140 110566
rect 274088 110502 274140 110508
rect 273996 109064 274048 109070
rect 273996 109006 274048 109012
rect 274008 66910 274036 109006
rect 274100 72554 274128 110502
rect 274088 72548 274140 72554
rect 274088 72490 274140 72496
rect 273996 66904 274048 66910
rect 273996 66846 274048 66852
rect 274652 16574 274680 144230
rect 274744 143546 274772 188294
rect 275296 177478 275324 232494
rect 276032 224874 276060 238726
rect 278056 238542 278084 240094
rect 279528 240094 279864 240122
rect 281552 240094 282440 240122
rect 279528 238678 279556 240094
rect 279516 238672 279568 238678
rect 279516 238614 279568 238620
rect 278044 238536 278096 238542
rect 278044 238478 278096 238484
rect 278056 231742 278084 238478
rect 279528 231742 279556 238614
rect 278044 231736 278096 231742
rect 278044 231678 278096 231684
rect 279516 231736 279568 231742
rect 279516 231678 279568 231684
rect 280068 231736 280120 231742
rect 280068 231678 280120 231684
rect 276020 224868 276072 224874
rect 276020 224810 276072 224816
rect 276032 224466 276060 224810
rect 276020 224460 276072 224466
rect 276020 224402 276072 224408
rect 276664 224460 276716 224466
rect 276664 224402 276716 224408
rect 276112 198076 276164 198082
rect 276112 198018 276164 198024
rect 275284 177472 275336 177478
rect 275284 177414 275336 177420
rect 275284 164280 275336 164286
rect 275284 164222 275336 164228
rect 274732 143540 274784 143546
rect 274732 143482 274784 143488
rect 275296 125526 275324 164222
rect 276020 153876 276072 153882
rect 276020 153818 276072 153824
rect 275468 141500 275520 141506
rect 275468 141442 275520 141448
rect 275284 125520 275336 125526
rect 275284 125462 275336 125468
rect 275376 124908 275428 124914
rect 275376 124850 275428 124856
rect 275388 113082 275416 124850
rect 275376 113076 275428 113082
rect 275376 113018 275428 113024
rect 275376 100836 275428 100842
rect 275376 100778 275428 100784
rect 275284 96756 275336 96762
rect 275284 96698 275336 96704
rect 275296 24138 275324 96698
rect 275388 28286 275416 100778
rect 275480 78062 275508 141442
rect 275468 78056 275520 78062
rect 275468 77998 275520 78004
rect 275376 28280 275428 28286
rect 275376 28222 275428 28228
rect 275284 24132 275336 24138
rect 275284 24074 275336 24080
rect 274652 16546 274864 16574
rect 273904 7676 273956 7682
rect 273904 7618 273956 7624
rect 274836 480 274864 16546
rect 276032 3602 276060 153818
rect 276124 137970 276152 198018
rect 276112 137964 276164 137970
rect 276112 137906 276164 137912
rect 276112 91792 276164 91798
rect 276112 91734 276164 91740
rect 276020 3596 276072 3602
rect 276020 3538 276072 3544
rect 276124 3482 276152 91734
rect 276676 78674 276704 224402
rect 278136 222896 278188 222902
rect 278136 222838 278188 222844
rect 277400 210588 277452 210594
rect 277400 210530 277452 210536
rect 277412 155922 277440 210530
rect 277492 198144 277544 198150
rect 277492 198086 277544 198092
rect 277400 155916 277452 155922
rect 277400 155858 277452 155864
rect 277504 147558 277532 198086
rect 278148 191826 278176 222838
rect 278780 203720 278832 203726
rect 278780 203662 278832 203668
rect 278136 191820 278188 191826
rect 278136 191762 278188 191768
rect 278044 191412 278096 191418
rect 278044 191354 278096 191360
rect 277492 147552 277544 147558
rect 277492 147494 277544 147500
rect 276664 78668 276716 78674
rect 276664 78610 276716 78616
rect 276756 3596 276808 3602
rect 276756 3538 276808 3544
rect 276032 3454 276152 3482
rect 276032 480 276060 3454
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276768 354 276796 3538
rect 278056 2922 278084 191354
rect 278228 165776 278280 165782
rect 278228 165718 278280 165724
rect 278136 128444 278188 128450
rect 278136 128386 278188 128392
rect 278148 19990 278176 128386
rect 278240 126886 278268 165718
rect 278792 149054 278820 203662
rect 280080 180198 280108 231678
rect 280896 217456 280948 217462
rect 280896 217398 280948 217404
rect 280160 209364 280212 209370
rect 280160 209306 280212 209312
rect 280068 180192 280120 180198
rect 280068 180134 280120 180140
rect 279424 168496 279476 168502
rect 279424 168438 279476 168444
rect 278780 149048 278832 149054
rect 278780 148990 278832 148996
rect 278320 142248 278372 142254
rect 278320 142190 278372 142196
rect 278228 126880 278280 126886
rect 278228 126822 278280 126828
rect 278228 124296 278280 124302
rect 278228 124238 278280 124244
rect 278136 19984 278188 19990
rect 278136 19926 278188 19932
rect 278240 18698 278268 124238
rect 278332 102134 278360 142190
rect 279436 140078 279464 168438
rect 279608 167136 279660 167142
rect 279608 167078 279660 167084
rect 279424 140072 279476 140078
rect 279424 140014 279476 140020
rect 279424 136740 279476 136746
rect 279424 136682 279476 136688
rect 278780 131776 278832 131782
rect 278780 131718 278832 131724
rect 278320 102128 278372 102134
rect 278320 102070 278372 102076
rect 278228 18692 278280 18698
rect 278228 18634 278280 18640
rect 278792 16574 278820 131718
rect 279436 17338 279464 136682
rect 279620 128314 279648 167078
rect 279700 158024 279752 158030
rect 279700 157966 279752 157972
rect 279608 128308 279660 128314
rect 279608 128250 279660 128256
rect 279516 127084 279568 127090
rect 279516 127026 279568 127032
rect 279528 73846 279556 127026
rect 279712 125458 279740 157966
rect 280172 140758 280200 209306
rect 280160 140752 280212 140758
rect 280160 140694 280212 140700
rect 280804 127152 280856 127158
rect 280804 127094 280856 127100
rect 279700 125452 279752 125458
rect 279700 125394 279752 125400
rect 280160 124976 280212 124982
rect 280160 124918 280212 124924
rect 279516 73840 279568 73846
rect 279516 73782 279568 73788
rect 279424 17332 279476 17338
rect 279424 17274 279476 17280
rect 280172 16574 280200 124918
rect 280816 17270 280844 127094
rect 280908 126274 280936 217398
rect 281552 206446 281580 240094
rect 284358 239850 284386 240108
rect 284312 239822 284386 239850
rect 285692 240094 286304 240122
rect 287900 240094 288236 240122
rect 290812 240094 291148 240122
rect 283656 216096 283708 216102
rect 283656 216038 283708 216044
rect 283564 213376 283616 213382
rect 283564 213318 283616 213324
rect 281540 206440 281592 206446
rect 281540 206382 281592 206388
rect 281540 205080 281592 205086
rect 281540 205022 281592 205028
rect 281080 161560 281132 161566
rect 281080 161502 281132 161508
rect 280988 132524 281040 132530
rect 280988 132466 281040 132472
rect 280896 126268 280948 126274
rect 280896 126210 280948 126216
rect 281000 58682 281028 132466
rect 281092 122738 281120 161502
rect 281552 147626 281580 205022
rect 283576 175982 283604 213318
rect 283668 182986 283696 216038
rect 283656 182980 283708 182986
rect 283656 182922 283708 182928
rect 283564 175976 283616 175982
rect 283564 175918 283616 175924
rect 283748 174072 283800 174078
rect 283748 174014 283800 174020
rect 283656 172712 283708 172718
rect 283656 172654 283708 172660
rect 282276 169924 282328 169930
rect 282276 169866 282328 169872
rect 281540 147620 281592 147626
rect 281540 147562 281592 147568
rect 282184 134020 282236 134026
rect 282184 133962 282236 133968
rect 281080 122732 281132 122738
rect 281080 122674 281132 122680
rect 280988 58676 281040 58682
rect 280988 58618 281040 58624
rect 282196 55962 282224 133962
rect 282288 131102 282316 169866
rect 282368 139528 282420 139534
rect 282368 139470 282420 139476
rect 282276 131096 282328 131102
rect 282276 131038 282328 131044
rect 282276 116068 282328 116074
rect 282276 116010 282328 116016
rect 282184 55956 282236 55962
rect 282184 55898 282236 55904
rect 282288 44878 282316 116010
rect 282380 98666 282408 139470
rect 283564 135380 283616 135386
rect 283564 135322 283616 135328
rect 282368 98660 282420 98666
rect 282368 98602 282420 98608
rect 282276 44872 282328 44878
rect 282276 44814 282328 44820
rect 280804 17264 280856 17270
rect 280804 17206 280856 17212
rect 278792 16546 279096 16574
rect 280172 16546 280752 16574
rect 278318 3360 278374 3369
rect 278318 3295 278374 3304
rect 278044 2916 278096 2922
rect 278044 2858 278096 2864
rect 278332 480 278360 3295
rect 277094 354 277206 480
rect 276768 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 280724 480 280752 16546
rect 281540 14544 281592 14550
rect 281540 14486 281592 14492
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281552 354 281580 14486
rect 283576 10334 283604 135322
rect 283668 135250 283696 172654
rect 283760 136610 283788 174014
rect 283840 146396 283892 146402
rect 283840 146338 283892 146344
rect 283748 136604 283800 136610
rect 283748 136546 283800 136552
rect 283656 135244 283708 135250
rect 283656 135186 283708 135192
rect 283748 121576 283800 121582
rect 283748 121518 283800 121524
rect 283656 104916 283708 104922
rect 283656 104858 283708 104864
rect 283564 10328 283616 10334
rect 283564 10270 283616 10276
rect 283668 8974 283696 104858
rect 283760 25634 283788 121518
rect 283852 106282 283880 146338
rect 283930 134464 283986 134473
rect 283930 134399 283986 134408
rect 283944 109002 283972 134399
rect 284312 113830 284340 239822
rect 284944 162172 284996 162178
rect 284944 162114 284996 162120
rect 284300 113824 284352 113830
rect 284300 113766 284352 113772
rect 283932 108996 283984 109002
rect 283932 108938 283984 108944
rect 283840 106276 283892 106282
rect 283840 106218 283892 106224
rect 283748 25628 283800 25634
rect 283748 25570 283800 25576
rect 284300 21548 284352 21554
rect 284300 21490 284352 21496
rect 283656 8968 283708 8974
rect 283656 8910 283708 8916
rect 283104 2916 283156 2922
rect 283104 2858 283156 2864
rect 283116 480 283144 2858
rect 284312 480 284340 21490
rect 284956 3670 284984 162114
rect 285036 135448 285088 135454
rect 285036 135390 285088 135396
rect 285048 9042 285076 135390
rect 285128 103692 285180 103698
rect 285128 103634 285180 103640
rect 285140 57254 285168 103634
rect 285128 57248 285180 57254
rect 285128 57190 285180 57196
rect 285036 9036 285088 9042
rect 285036 8978 285088 8984
rect 285692 6914 285720 240094
rect 287702 238912 287758 238921
rect 287702 238847 287758 238856
rect 287716 215286 287744 238847
rect 287900 238785 287928 240094
rect 289820 239896 289872 239902
rect 289820 239838 289872 239844
rect 287886 238776 287942 238785
rect 287886 238711 287942 238720
rect 287900 238678 287928 238711
rect 287888 238672 287940 238678
rect 287888 238614 287940 238620
rect 289084 217524 289136 217530
rect 289084 217466 289136 217472
rect 287704 215280 287756 215286
rect 287704 215222 287756 215228
rect 289096 178770 289124 217466
rect 289084 178764 289136 178770
rect 289084 178706 289136 178712
rect 289452 171284 289504 171290
rect 289452 171226 289504 171232
rect 289268 162988 289320 162994
rect 289268 162930 289320 162936
rect 287704 161628 287756 161634
rect 287704 161570 287756 161576
rect 286416 131232 286468 131238
rect 286416 131174 286468 131180
rect 286324 129872 286376 129878
rect 286324 129814 286376 129820
rect 286336 37942 286364 129814
rect 286428 64190 286456 131174
rect 287716 122806 287744 161570
rect 289084 158908 289136 158914
rect 289084 158850 289136 158856
rect 287888 155304 287940 155310
rect 287888 155246 287940 155252
rect 287796 122868 287848 122874
rect 287796 122810 287848 122816
rect 287704 122800 287756 122806
rect 287704 122742 287756 122748
rect 287704 118720 287756 118726
rect 287704 118662 287756 118668
rect 286416 64184 286468 64190
rect 286416 64126 286468 64132
rect 286324 37936 286376 37942
rect 286324 37878 286376 37884
rect 287058 27024 287114 27033
rect 287058 26959 287114 26968
rect 285770 26888 285826 26897
rect 285770 26823 285826 26832
rect 285784 16574 285812 26823
rect 287072 16574 287100 26959
rect 285784 16546 286640 16574
rect 287072 16546 287376 16574
rect 285416 6886 285720 6914
rect 284944 3664 284996 3670
rect 284944 3606 284996 3612
rect 285416 480 285444 6886
rect 286612 480 286640 16546
rect 281878 354 281990 480
rect 281552 326 281990 354
rect 281878 -960 281990 326
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287348 354 287376 16546
rect 287716 6186 287744 118662
rect 287808 42158 287836 122810
rect 287900 115870 287928 155246
rect 287978 145616 288034 145625
rect 287978 145551 288034 145560
rect 287992 117298 288020 145551
rect 289096 120086 289124 158850
rect 289176 132592 289228 132598
rect 289176 132534 289228 132540
rect 289084 120080 289136 120086
rect 289084 120022 289136 120028
rect 287980 117292 288032 117298
rect 287980 117234 288032 117240
rect 287888 115864 287940 115870
rect 287888 115806 287940 115812
rect 289084 113348 289136 113354
rect 289084 113290 289136 113296
rect 287888 100904 287940 100910
rect 287888 100846 287940 100852
rect 287796 42152 287848 42158
rect 287796 42094 287848 42100
rect 287900 31074 287928 100846
rect 287888 31068 287940 31074
rect 287888 31010 287940 31016
rect 289096 29646 289124 113290
rect 289188 61470 289216 132534
rect 289280 124098 289308 162930
rect 289360 150544 289412 150550
rect 289360 150486 289412 150492
rect 289268 124092 289320 124098
rect 289268 124034 289320 124040
rect 289268 117360 289320 117366
rect 289268 117302 289320 117308
rect 289280 68338 289308 117302
rect 289372 110362 289400 150486
rect 289464 133890 289492 171226
rect 289452 133884 289504 133890
rect 289452 133826 289504 133832
rect 289360 110356 289412 110362
rect 289360 110298 289412 110304
rect 289268 68332 289320 68338
rect 289268 68274 289320 68280
rect 289176 61464 289228 61470
rect 289176 61406 289228 61412
rect 289084 29640 289136 29646
rect 289084 29582 289136 29588
rect 287704 6180 287756 6186
rect 287704 6122 287756 6128
rect 288992 3596 289044 3602
rect 288992 3538 289044 3544
rect 289004 480 289032 3538
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 289832 354 289860 239838
rect 291120 238785 291148 240094
rect 291106 238776 291162 238785
rect 291106 238711 291162 238720
rect 291844 225616 291896 225622
rect 291844 225558 291896 225564
rect 291200 217388 291252 217394
rect 291200 217330 291252 217336
rect 290648 156664 290700 156670
rect 290648 156606 290700 156612
rect 290556 131300 290608 131306
rect 290556 131242 290608 131248
rect 290464 121644 290516 121650
rect 290464 121586 290516 121592
rect 290476 22846 290504 121586
rect 290568 62898 290596 131242
rect 290660 118658 290688 156606
rect 290648 118652 290700 118658
rect 290648 118594 290700 118600
rect 290556 62892 290608 62898
rect 290556 62834 290608 62840
rect 290464 22840 290516 22846
rect 290464 22782 290516 22788
rect 291212 16574 291240 217330
rect 291856 124982 291884 225558
rect 291948 153882 291976 240586
rect 292592 240094 292744 240122
rect 292028 164348 292080 164354
rect 292028 164290 292080 164296
rect 291936 153876 291988 153882
rect 291936 153818 291988 153824
rect 292040 126954 292068 164290
rect 292028 126948 292080 126954
rect 292028 126890 292080 126896
rect 291936 125724 291988 125730
rect 291936 125666 291988 125672
rect 291844 124976 291896 124982
rect 291844 124918 291896 124924
rect 291844 120216 291896 120222
rect 291844 120158 291896 120164
rect 291856 39370 291884 120158
rect 291948 53106 291976 125666
rect 292028 102264 292080 102270
rect 292028 102206 292080 102212
rect 291936 53100 291988 53106
rect 291936 53042 291988 53048
rect 292040 43450 292068 102206
rect 292592 95946 292620 240094
rect 293052 131782 293080 268087
rect 293144 155242 293172 287671
rect 293236 231674 293264 300834
rect 293958 299296 294014 299305
rect 293958 299231 294014 299240
rect 293314 241496 293370 241505
rect 293314 241431 293370 241440
rect 293328 240650 293356 241431
rect 293316 240644 293368 240650
rect 293316 240586 293368 240592
rect 293224 231668 293276 231674
rect 293224 231610 293276 231616
rect 293132 155236 293184 155242
rect 293132 155178 293184 155184
rect 293408 143608 293460 143614
rect 293408 143550 293460 143556
rect 293040 131776 293092 131782
rect 293040 131718 293092 131724
rect 293224 122936 293276 122942
rect 293224 122878 293276 122884
rect 292672 101448 292724 101454
rect 292672 101390 292724 101396
rect 292580 95940 292632 95946
rect 292580 95882 292632 95888
rect 292028 43444 292080 43450
rect 292028 43386 292080 43392
rect 291844 39364 291896 39370
rect 291844 39306 291896 39312
rect 292684 16574 292712 101390
rect 293236 28354 293264 122878
rect 293316 114640 293368 114646
rect 293316 114582 293368 114588
rect 293328 50386 293356 114582
rect 293420 102814 293448 143550
rect 293408 102808 293460 102814
rect 293408 102750 293460 102756
rect 293972 86290 294000 299231
rect 294050 263936 294106 263945
rect 294050 263871 294106 263880
rect 293960 86284 294012 86290
rect 293960 86226 294012 86232
rect 294064 79422 294092 263871
rect 294156 225690 294184 325751
rect 294234 323096 294290 323105
rect 294234 323031 294290 323040
rect 294248 239902 294276 323031
rect 295338 321056 295394 321065
rect 295338 320991 295394 321000
rect 295352 320210 295380 320991
rect 295340 320204 295392 320210
rect 295340 320146 295392 320152
rect 295338 319016 295394 319025
rect 295338 318951 295394 318960
rect 295352 318850 295380 318951
rect 295340 318844 295392 318850
rect 295340 318786 295392 318792
rect 295340 317416 295392 317422
rect 295340 317358 295392 317364
rect 295352 316985 295380 317358
rect 295338 316976 295394 316985
rect 295338 316911 295394 316920
rect 295338 314256 295394 314265
rect 295338 314191 295394 314200
rect 295352 313954 295380 314191
rect 295340 313948 295392 313954
rect 295340 313890 295392 313896
rect 295338 311944 295394 311953
rect 295338 311879 295340 311888
rect 295392 311879 295394 311888
rect 295340 311850 295392 311856
rect 295340 310480 295392 310486
rect 295340 310422 295392 310428
rect 295352 310185 295380 310422
rect 295338 310176 295394 310185
rect 295338 310111 295394 310120
rect 295338 308136 295394 308145
rect 295338 308071 295394 308080
rect 295352 307834 295380 308071
rect 295340 307828 295392 307834
rect 295340 307770 295392 307776
rect 295338 305416 295394 305425
rect 295338 305351 295394 305360
rect 295352 305046 295380 305351
rect 295340 305040 295392 305046
rect 295340 304982 295392 304988
rect 295340 303612 295392 303618
rect 295340 303554 295392 303560
rect 295352 303385 295380 303554
rect 295338 303376 295394 303385
rect 295338 303311 295394 303320
rect 296076 300144 296128 300150
rect 296076 300086 296128 300092
rect 295338 296576 295394 296585
rect 295338 296511 295394 296520
rect 295352 295390 295380 296511
rect 295340 295384 295392 295390
rect 295340 295326 295392 295332
rect 295338 294536 295394 294545
rect 295338 294471 295394 294480
rect 295352 294030 295380 294471
rect 295340 294024 295392 294030
rect 295340 293966 295392 293972
rect 296088 290465 296116 300086
rect 296626 292496 296682 292505
rect 296732 292482 296760 359042
rect 296824 313954 296852 360334
rect 296916 331906 296944 364346
rect 298284 363044 298336 363050
rect 298284 362986 298336 362992
rect 297364 360596 297416 360602
rect 297364 360538 297416 360544
rect 296904 331900 296956 331906
rect 296904 331842 296956 331848
rect 296812 313948 296864 313954
rect 296812 313890 296864 313896
rect 296682 292454 296760 292482
rect 296626 292431 296682 292440
rect 296074 290456 296130 290465
rect 296074 290391 296130 290400
rect 296732 287706 296760 292454
rect 296720 287700 296772 287706
rect 296720 287642 296772 287648
rect 295340 285728 295392 285734
rect 295338 285696 295340 285705
rect 295392 285696 295394 285705
rect 295338 285631 295394 285640
rect 295338 283656 295394 283665
rect 295338 283591 295394 283600
rect 295352 282946 295380 283591
rect 295340 282940 295392 282946
rect 295340 282882 295392 282888
rect 295352 281738 295380 282882
rect 295352 281710 295472 281738
rect 295338 281616 295394 281625
rect 295338 281551 295340 281560
rect 295392 281551 295394 281560
rect 295340 281522 295392 281528
rect 295338 278896 295394 278905
rect 295338 278831 295340 278840
rect 295392 278831 295394 278840
rect 295340 278802 295392 278808
rect 295338 276856 295394 276865
rect 295338 276791 295394 276800
rect 295352 276078 295380 276791
rect 295340 276072 295392 276078
rect 295340 276014 295392 276020
rect 295338 274816 295394 274825
rect 295338 274751 295394 274760
rect 295352 274718 295380 274751
rect 295340 274712 295392 274718
rect 295340 274654 295392 274660
rect 295338 272776 295394 272785
rect 295338 272711 295394 272720
rect 295352 271930 295380 272711
rect 295340 271924 295392 271930
rect 295340 271866 295392 271872
rect 295338 270056 295394 270065
rect 295338 269991 295394 270000
rect 295352 269142 295380 269991
rect 295340 269136 295392 269142
rect 295340 269078 295392 269084
rect 295338 265976 295394 265985
rect 295338 265911 295394 265920
rect 295352 264246 295380 265911
rect 295340 264240 295392 264246
rect 295340 264182 295392 264188
rect 295338 261216 295394 261225
rect 295338 261151 295340 261160
rect 295392 261151 295394 261160
rect 295340 261122 295392 261128
rect 295338 259176 295394 259185
rect 295338 259111 295394 259120
rect 294236 239896 294288 239902
rect 294236 239838 294288 239844
rect 294144 225684 294196 225690
rect 294144 225626 294196 225632
rect 295352 144294 295380 259111
rect 295444 237182 295472 281710
rect 295524 281580 295576 281586
rect 295524 281522 295576 281528
rect 295536 248414 295564 281522
rect 295984 275392 296036 275398
rect 295984 275334 296036 275340
rect 295996 257145 296024 275334
rect 295982 257136 296038 257145
rect 295982 257071 296038 257080
rect 295614 255096 295670 255105
rect 295614 255031 295670 255040
rect 295628 253978 295656 255031
rect 295616 253972 295668 253978
rect 295616 253914 295668 253920
rect 295536 248386 295656 248414
rect 295522 248296 295578 248305
rect 295522 248231 295578 248240
rect 295536 247110 295564 248231
rect 295524 247104 295576 247110
rect 295524 247046 295576 247052
rect 295524 246356 295576 246362
rect 295524 246298 295576 246304
rect 295536 246265 295564 246298
rect 295522 246256 295578 246265
rect 295522 246191 295578 246200
rect 295628 239426 295656 248386
rect 295800 244248 295852 244254
rect 295800 244190 295852 244196
rect 295812 243545 295840 244190
rect 295798 243536 295854 243545
rect 295798 243471 295854 243480
rect 295616 239420 295668 239426
rect 295616 239362 295668 239368
rect 295996 238754 296024 257071
rect 297180 252272 297232 252278
rect 297180 252214 297232 252220
rect 297192 252113 297220 252214
rect 296534 252104 296590 252113
rect 296534 252039 296590 252048
rect 297178 252104 297234 252113
rect 297178 252039 297234 252048
rect 296548 248441 296576 252039
rect 296626 250336 296682 250345
rect 296682 250294 296760 250322
rect 296626 250271 296682 250280
rect 296534 248432 296590 248441
rect 296534 248367 296590 248376
rect 296732 242214 296760 250294
rect 296720 242208 296772 242214
rect 296720 242150 296772 242156
rect 295628 238726 296024 238754
rect 295432 237176 295484 237182
rect 295432 237118 295484 237124
rect 295628 233170 295656 238726
rect 295616 233164 295668 233170
rect 295616 233106 295668 233112
rect 296260 153400 296312 153406
rect 296260 153342 296312 153348
rect 295984 149728 296036 149734
rect 295984 149670 296036 149676
rect 295340 144288 295392 144294
rect 295340 144230 295392 144236
rect 295996 124166 296024 149670
rect 296076 124364 296128 124370
rect 296076 124306 296128 124312
rect 295984 124160 296036 124166
rect 295984 124102 296036 124108
rect 294604 123004 294656 123010
rect 294604 122946 294656 122952
rect 294052 79416 294104 79422
rect 294052 79358 294104 79364
rect 293316 50380 293368 50386
rect 293316 50322 293368 50328
rect 293960 38072 294012 38078
rect 293960 38014 294012 38020
rect 293224 28348 293276 28354
rect 293224 28290 293276 28296
rect 293972 16574 294000 38014
rect 294616 33794 294644 122946
rect 295984 111852 296036 111858
rect 295984 111794 296036 111800
rect 294604 33788 294656 33794
rect 294604 33730 294656 33736
rect 291212 16546 291424 16574
rect 292684 16546 293264 16574
rect 293972 16546 294920 16574
rect 291396 480 291424 16546
rect 292580 3460 292632 3466
rect 292580 3402 292632 3408
rect 292592 480 292620 3402
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 294892 480 294920 16546
rect 295996 2174 296024 111794
rect 296088 20058 296116 124306
rect 296168 118788 296220 118794
rect 296168 118730 296220 118736
rect 296180 72486 296208 118730
rect 296272 113150 296300 153342
rect 296260 113144 296312 113150
rect 296260 113086 296312 113092
rect 296260 103624 296312 103630
rect 296260 103566 296312 103572
rect 296168 72480 296220 72486
rect 296168 72422 296220 72428
rect 296272 60042 296300 103566
rect 296720 71188 296772 71194
rect 296720 71130 296772 71136
rect 296260 60036 296312 60042
rect 296260 59978 296312 59984
rect 296076 20052 296128 20058
rect 296076 19994 296128 20000
rect 296732 16574 296760 71130
rect 296732 16546 297312 16574
rect 296074 3360 296130 3369
rect 296074 3295 296130 3304
rect 295984 2168 296036 2174
rect 295984 2110 296036 2116
rect 296088 480 296116 3295
rect 297284 480 297312 16546
rect 297376 3398 297404 360538
rect 298100 357672 298152 357678
rect 298100 357614 298152 357620
rect 297548 280356 297600 280362
rect 297548 280298 297600 280304
rect 297456 261180 297508 261186
rect 297456 261122 297508 261128
rect 297468 79354 297496 261122
rect 297560 238406 297588 280298
rect 297548 238400 297600 238406
rect 297548 238342 297600 238348
rect 297548 160268 297600 160274
rect 297548 160210 297600 160216
rect 297560 121446 297588 160210
rect 298112 141506 298140 357614
rect 298192 354952 298244 354958
rect 298192 354894 298244 354900
rect 298204 303618 298232 354894
rect 298296 336734 298324 362986
rect 298284 336728 298336 336734
rect 298284 336670 298336 336676
rect 299388 336728 299440 336734
rect 299388 336670 299440 336676
rect 299400 336054 299428 336670
rect 299388 336048 299440 336054
rect 299388 335990 299440 335996
rect 298192 303612 298244 303618
rect 298192 303554 298244 303560
rect 298928 285728 298980 285734
rect 298928 285670 298980 285676
rect 298836 278860 298888 278866
rect 298836 278802 298888 278808
rect 298744 274712 298796 274718
rect 298744 274654 298796 274660
rect 298192 246356 298244 246362
rect 298192 246298 298244 246304
rect 298204 223446 298232 246298
rect 298756 239970 298784 274654
rect 298848 253230 298876 278802
rect 298940 267102 298968 285670
rect 298928 267096 298980 267102
rect 298928 267038 298980 267044
rect 298928 253972 298980 253978
rect 298928 253914 298980 253920
rect 298836 253224 298888 253230
rect 298836 253166 298888 253172
rect 298940 240786 298968 253914
rect 299492 240825 299520 700266
rect 299572 361752 299624 361758
rect 299572 361694 299624 361700
rect 299584 317422 299612 361694
rect 300860 357808 300912 357814
rect 300860 357750 300912 357756
rect 300124 356448 300176 356454
rect 300124 356390 300176 356396
rect 299572 317416 299624 317422
rect 299572 317358 299624 317364
rect 299572 253224 299624 253230
rect 299572 253166 299624 253172
rect 299478 240816 299534 240825
rect 298928 240780 298980 240786
rect 299478 240751 299534 240760
rect 298928 240722 298980 240728
rect 298744 239964 298796 239970
rect 298744 239906 298796 239912
rect 298192 223440 298244 223446
rect 298192 223382 298244 223388
rect 298744 143676 298796 143682
rect 298744 143618 298796 143624
rect 298100 141500 298152 141506
rect 298100 141442 298152 141448
rect 297730 140040 297786 140049
rect 297730 139975 297786 139984
rect 297548 121440 297600 121446
rect 297548 121382 297600 121388
rect 297640 120284 297692 120290
rect 297640 120226 297692 120232
rect 297548 99408 297600 99414
rect 297548 99350 297600 99356
rect 297456 79348 297508 79354
rect 297456 79290 297508 79296
rect 297560 36582 297588 99350
rect 297652 65618 297680 120226
rect 297744 100706 297772 139975
rect 298756 119406 298784 143618
rect 299112 140820 299164 140826
rect 299112 140762 299164 140768
rect 298928 129940 298980 129946
rect 298928 129882 298980 129888
rect 298744 119400 298796 119406
rect 298744 119342 298796 119348
rect 298744 116136 298796 116142
rect 298744 116078 298796 116084
rect 297732 100700 297784 100706
rect 297732 100642 297784 100648
rect 297640 65612 297692 65618
rect 297640 65554 297692 65560
rect 297548 36576 297600 36582
rect 297548 36518 297600 36524
rect 298756 32434 298784 116078
rect 298836 98116 298888 98122
rect 298836 98058 298888 98064
rect 298744 32428 298796 32434
rect 298744 32370 298796 32376
rect 298848 25566 298876 98058
rect 298940 65550 298968 129882
rect 299020 111920 299072 111926
rect 299020 111862 299072 111868
rect 298928 65544 298980 65550
rect 298928 65486 298980 65492
rect 299032 53174 299060 111862
rect 299124 99278 299152 140762
rect 299112 99272 299164 99278
rect 299112 99214 299164 99220
rect 299020 53168 299072 53174
rect 299020 53110 299072 53116
rect 298928 35352 298980 35358
rect 298928 35294 298980 35300
rect 298836 25560 298888 25566
rect 298836 25502 298888 25508
rect 298468 3664 298520 3670
rect 298468 3606 298520 3612
rect 297364 3392 297416 3398
rect 297364 3334 297416 3340
rect 298480 480 298508 3606
rect 298940 3466 298968 35294
rect 299480 10396 299532 10402
rect 299480 10338 299532 10344
rect 299492 3482 299520 10338
rect 299584 3602 299612 253166
rect 300136 197334 300164 356390
rect 300768 317416 300820 317422
rect 300768 317358 300820 317364
rect 300780 316742 300808 317358
rect 300768 316736 300820 316742
rect 300768 316678 300820 316684
rect 300216 300892 300268 300898
rect 300216 300834 300268 300840
rect 300228 294642 300256 300834
rect 300216 294636 300268 294642
rect 300216 294578 300268 294584
rect 300216 278996 300268 279002
rect 300216 278938 300268 278944
rect 300228 238474 300256 278938
rect 300216 238468 300268 238474
rect 300216 238410 300268 238416
rect 300216 206304 300268 206310
rect 300216 206246 300268 206252
rect 300124 197328 300176 197334
rect 300124 197270 300176 197276
rect 300228 180266 300256 206246
rect 300216 180260 300268 180266
rect 300216 180202 300268 180208
rect 300216 154692 300268 154698
rect 300216 154634 300268 154640
rect 300124 117496 300176 117502
rect 300124 117438 300176 117444
rect 300136 13122 300164 117438
rect 300228 115938 300256 154634
rect 300872 129033 300900 357750
rect 300952 357468 301004 357474
rect 300952 357410 301004 357416
rect 300964 310486 300992 357410
rect 300952 310480 301004 310486
rect 300952 310422 301004 310428
rect 301320 310480 301372 310486
rect 301320 310422 301372 310428
rect 301332 309806 301360 310422
rect 301320 309800 301372 309806
rect 301320 309742 301372 309748
rect 302068 284374 302096 700266
rect 307668 698964 307720 698970
rect 307668 698906 307720 698912
rect 305734 510640 305790 510649
rect 305734 510575 305790 510584
rect 302240 364608 302292 364614
rect 302240 364550 302292 364556
rect 302148 294024 302200 294030
rect 302148 293966 302200 293972
rect 302160 289882 302188 293966
rect 302148 289876 302200 289882
rect 302148 289818 302200 289824
rect 301504 284368 301556 284374
rect 301504 284310 301556 284316
rect 302056 284368 302108 284374
rect 302056 284310 302108 284316
rect 301320 276684 301372 276690
rect 301320 276626 301372 276632
rect 301332 276078 301360 276626
rect 300952 276072 301004 276078
rect 300952 276014 301004 276020
rect 301320 276072 301372 276078
rect 301320 276014 301372 276020
rect 300964 231849 300992 276014
rect 301516 252278 301544 284310
rect 302160 253910 302188 289818
rect 302148 253904 302200 253910
rect 302148 253846 302200 253852
rect 301504 252272 301556 252278
rect 301504 252214 301556 252220
rect 301320 247716 301372 247722
rect 301320 247658 301372 247664
rect 301332 247110 301360 247658
rect 301044 247104 301096 247110
rect 301044 247046 301096 247052
rect 301320 247104 301372 247110
rect 301320 247046 301372 247052
rect 300950 231840 301006 231849
rect 300950 231775 301006 231784
rect 301056 224777 301084 247046
rect 301042 224768 301098 224777
rect 301042 224703 301098 224712
rect 301596 146464 301648 146470
rect 301596 146406 301648 146412
rect 301504 142316 301556 142322
rect 301504 142258 301556 142264
rect 300858 129024 300914 129033
rect 300858 128959 300914 128968
rect 300216 115932 300268 115938
rect 300216 115874 300268 115880
rect 300216 110628 300268 110634
rect 300216 110570 300268 110576
rect 300228 51814 300256 110570
rect 300308 107840 300360 107846
rect 300308 107782 300360 107788
rect 300216 51808 300268 51814
rect 300216 51750 300268 51756
rect 300320 49094 300348 107782
rect 301516 105602 301544 142258
rect 301608 117978 301636 146406
rect 301596 117972 301648 117978
rect 301596 117914 301648 117920
rect 301780 117428 301832 117434
rect 301780 117370 301832 117376
rect 301596 109200 301648 109206
rect 301596 109142 301648 109148
rect 301504 105596 301556 105602
rect 301504 105538 301556 105544
rect 301504 98184 301556 98190
rect 301504 98126 301556 98132
rect 300308 49088 300360 49094
rect 300308 49030 300360 49036
rect 300124 13116 300176 13122
rect 300124 13058 300176 13064
rect 301516 7614 301544 98126
rect 301608 26926 301636 109142
rect 301688 104984 301740 104990
rect 301688 104926 301740 104932
rect 301700 55894 301728 104926
rect 301792 73914 301820 117370
rect 302252 101454 302280 364550
rect 305644 358964 305696 358970
rect 305644 358906 305696 358912
rect 305092 357400 305144 357406
rect 305092 357342 305144 357348
rect 303620 356380 303672 356386
rect 303620 356322 303672 356328
rect 302884 295384 302936 295390
rect 302884 295326 302936 295332
rect 302240 101448 302292 101454
rect 302240 101390 302292 101396
rect 302896 87650 302924 295326
rect 303632 193905 303660 356322
rect 305104 356182 305132 357342
rect 305092 356176 305144 356182
rect 305092 356118 305144 356124
rect 305000 354748 305052 354754
rect 305000 354690 305052 354696
rect 303618 193896 303674 193905
rect 303618 193831 303674 193840
rect 305012 152522 305040 354690
rect 305104 300150 305132 356118
rect 305092 300144 305144 300150
rect 305092 300086 305144 300092
rect 305656 178702 305684 358906
rect 305748 357406 305776 510575
rect 307024 365832 307076 365838
rect 307024 365774 307076 365780
rect 305736 357400 305788 357406
rect 305736 357342 305788 357348
rect 306472 271924 306524 271930
rect 306472 271866 306524 271872
rect 306288 267028 306340 267034
rect 306288 266970 306340 266976
rect 306300 191894 306328 266970
rect 306380 253904 306432 253910
rect 306380 253846 306432 253852
rect 306288 191888 306340 191894
rect 306288 191830 306340 191836
rect 305644 178696 305696 178702
rect 305644 178638 305696 178644
rect 306392 175953 306420 253846
rect 306484 233209 306512 271866
rect 306470 233200 306526 233209
rect 306470 233135 306526 233144
rect 307036 176050 307064 365774
rect 307680 247722 307708 698906
rect 307760 356720 307812 356726
rect 307760 356662 307812 356668
rect 307668 247716 307720 247722
rect 307668 247658 307720 247664
rect 307024 176044 307076 176050
rect 307024 175986 307076 175992
rect 306378 175944 306434 175953
rect 306378 175879 306434 175888
rect 306746 174856 306802 174865
rect 306746 174791 306802 174800
rect 306760 174010 306788 174791
rect 307666 174448 307722 174457
rect 307666 174383 307722 174392
rect 307300 174072 307352 174078
rect 307298 174040 307300 174049
rect 307352 174040 307354 174049
rect 306748 174004 306800 174010
rect 307298 173975 307354 173984
rect 306748 173946 306800 173952
rect 307680 173942 307708 174383
rect 307668 173936 307720 173942
rect 307668 173878 307720 173884
rect 307574 173632 307630 173641
rect 307574 173567 307630 173576
rect 307298 173224 307354 173233
rect 307298 173159 307354 173168
rect 307312 172650 307340 173159
rect 307588 172718 307616 173567
rect 307576 172712 307628 172718
rect 307576 172654 307628 172660
rect 307666 172680 307722 172689
rect 307300 172644 307352 172650
rect 307666 172615 307722 172624
rect 307300 172586 307352 172592
rect 307680 172582 307708 172615
rect 307668 172576 307720 172582
rect 307668 172518 307720 172524
rect 306930 172272 306986 172281
rect 306930 172207 306986 172216
rect 306562 171864 306618 171873
rect 306562 171799 306618 171808
rect 306576 171154 306604 171799
rect 306944 171290 306972 172207
rect 307666 171456 307722 171465
rect 307666 171391 307722 171400
rect 306932 171284 306984 171290
rect 306932 171226 306984 171232
rect 307680 171222 307708 171391
rect 307668 171216 307720 171222
rect 307668 171158 307720 171164
rect 306564 171148 306616 171154
rect 306564 171090 306616 171096
rect 307390 171048 307446 171057
rect 307390 170983 307446 170992
rect 306746 170640 306802 170649
rect 306746 170575 306802 170584
rect 306760 169794 306788 170575
rect 307300 169856 307352 169862
rect 307298 169824 307300 169833
rect 307352 169824 307354 169833
rect 306748 169788 306800 169794
rect 307298 169759 307354 169768
rect 306748 169730 306800 169736
rect 306746 169280 306802 169289
rect 306746 169215 306802 169224
rect 306760 168502 306788 169215
rect 306748 168496 306800 168502
rect 306748 168438 306800 168444
rect 307298 168464 307354 168473
rect 307298 168399 307300 168408
rect 307352 168399 307354 168408
rect 307300 168370 307352 168376
rect 307298 168056 307354 168065
rect 307298 167991 307354 168000
rect 306562 166424 306618 166433
rect 306562 166359 306618 166368
rect 306576 165782 306604 166359
rect 306564 165776 306616 165782
rect 306564 165718 306616 165724
rect 307114 165064 307170 165073
rect 307114 164999 307170 165008
rect 306746 162480 306802 162489
rect 306746 162415 306802 162424
rect 306760 161634 306788 162415
rect 306748 161628 306800 161634
rect 306748 161570 306800 161576
rect 306746 161256 306802 161265
rect 306746 161191 306802 161200
rect 306760 160206 306788 161191
rect 306748 160200 306800 160206
rect 306748 160142 306800 160148
rect 306746 157040 306802 157049
rect 306746 156975 306802 156984
rect 306760 155990 306788 156975
rect 306930 156224 306986 156233
rect 306930 156159 306986 156168
rect 306748 155984 306800 155990
rect 306748 155926 306800 155932
rect 306944 155310 306972 156159
rect 306932 155304 306984 155310
rect 306932 155246 306984 155252
rect 306562 154048 306618 154057
rect 306562 153983 306618 153992
rect 306576 153270 306604 153983
rect 307022 153640 307078 153649
rect 307022 153575 307078 153584
rect 306564 153264 306616 153270
rect 306564 153206 306616 153212
rect 306562 152688 306618 152697
rect 306562 152623 306618 152632
rect 305000 152516 305052 152522
rect 305000 152458 305052 152464
rect 306576 151910 306604 152623
rect 306564 151904 306616 151910
rect 306564 151846 306616 151852
rect 304356 150612 304408 150618
rect 304356 150554 304408 150560
rect 304264 135312 304316 135318
rect 304264 135254 304316 135260
rect 303160 130008 303212 130014
rect 303160 129950 303212 129956
rect 302976 118856 303028 118862
rect 302976 118798 303028 118804
rect 302884 87644 302936 87650
rect 302884 87586 302936 87592
rect 301780 73908 301832 73914
rect 301780 73850 301832 73856
rect 301688 55888 301740 55894
rect 301688 55830 301740 55836
rect 302988 31142 303016 118798
rect 303068 100972 303120 100978
rect 303068 100914 303120 100920
rect 302976 31136 303028 31142
rect 302976 31078 303028 31084
rect 301596 26920 301648 26926
rect 301596 26862 301648 26868
rect 303080 14482 303108 100914
rect 303172 54534 303200 129950
rect 303160 54528 303212 54534
rect 303160 54470 303212 54476
rect 304276 46238 304304 135254
rect 304368 110430 304396 150554
rect 306930 149288 306986 149297
rect 306930 149223 306986 149232
rect 306944 146946 306972 149223
rect 306932 146940 306984 146946
rect 306932 146882 306984 146888
rect 306562 145888 306618 145897
rect 306562 145823 306618 145832
rect 305734 145480 305790 145489
rect 305734 145415 305790 145424
rect 305642 124672 305698 124681
rect 305642 124607 305698 124616
rect 304356 110424 304408 110430
rect 304356 110366 304408 110372
rect 304540 109132 304592 109138
rect 304540 109074 304592 109080
rect 304448 107704 304500 107710
rect 304448 107646 304500 107652
rect 304356 102332 304408 102338
rect 304356 102274 304408 102280
rect 304368 62830 304396 102274
rect 304460 69698 304488 107646
rect 304552 71126 304580 109074
rect 304540 71120 304592 71126
rect 304540 71062 304592 71068
rect 304448 69692 304500 69698
rect 304448 69634 304500 69640
rect 304356 62824 304408 62830
rect 304356 62766 304408 62772
rect 304264 46232 304316 46238
rect 304264 46174 304316 46180
rect 303068 14476 303120 14482
rect 303068 14418 303120 14424
rect 305656 11830 305684 124607
rect 305748 104854 305776 145415
rect 306576 145042 306604 145823
rect 306932 145104 306984 145110
rect 306930 145072 306932 145081
rect 306984 145072 306986 145081
rect 306564 145036 306616 145042
rect 306930 145007 306986 145016
rect 306564 144978 306616 144984
rect 306930 144664 306986 144673
rect 306930 144599 306986 144608
rect 306562 144256 306618 144265
rect 306562 144191 306618 144200
rect 306010 140856 306066 140865
rect 306010 140791 306066 140800
rect 305826 106312 305882 106321
rect 305826 106247 305882 106256
rect 305736 104848 305788 104854
rect 305736 104790 305788 104796
rect 305734 99512 305790 99521
rect 305734 99447 305790 99456
rect 305748 35222 305776 99447
rect 305840 44946 305868 106247
rect 305918 103864 305974 103873
rect 305918 103799 305974 103808
rect 305932 61402 305960 103799
rect 306024 100026 306052 140791
rect 306576 137290 306604 144191
rect 306944 143682 306972 144599
rect 306932 143676 306984 143682
rect 306932 143618 306984 143624
rect 306746 142488 306802 142497
rect 306746 142423 306802 142432
rect 306760 142322 306788 142423
rect 306748 142316 306800 142322
rect 306748 142258 306800 142264
rect 306930 139088 306986 139097
rect 306930 139023 306986 139032
rect 306944 138038 306972 139023
rect 306932 138032 306984 138038
rect 306932 137974 306984 137980
rect 306930 137864 306986 137873
rect 306930 137799 306986 137808
rect 306564 137284 306616 137290
rect 306564 137226 306616 137232
rect 306944 136746 306972 137799
rect 306932 136740 306984 136746
rect 306932 136682 306984 136688
rect 306930 136640 306986 136649
rect 306930 136575 306986 136584
rect 306944 135522 306972 136575
rect 306932 135516 306984 135522
rect 306932 135458 306984 135464
rect 306746 134872 306802 134881
rect 306746 134807 306802 134816
rect 306760 134026 306788 134807
rect 306748 134020 306800 134026
rect 306748 133962 306800 133968
rect 306930 133648 306986 133657
rect 306930 133583 306986 133592
rect 306944 132530 306972 133583
rect 306932 132524 306984 132530
rect 306932 132466 306984 132472
rect 306746 131064 306802 131073
rect 306746 130999 306802 131008
rect 306760 130014 306788 130999
rect 306748 130008 306800 130014
rect 306748 129950 306800 129956
rect 306746 125488 306802 125497
rect 306746 125423 306802 125432
rect 306760 124438 306788 125423
rect 307036 124914 307064 153575
rect 307128 141438 307156 164999
rect 307312 164898 307340 167991
rect 307300 164892 307352 164898
rect 307300 164834 307352 164840
rect 307298 164248 307354 164257
rect 307298 164183 307354 164192
rect 307206 163024 307262 163033
rect 307206 162959 307262 162968
rect 307220 149734 307248 162959
rect 307312 158030 307340 164183
rect 307404 163538 307432 170983
rect 307666 170232 307722 170241
rect 307666 170167 307722 170176
rect 307680 169930 307708 170167
rect 307668 169924 307720 169930
rect 307668 169866 307720 169872
rect 307574 168872 307630 168881
rect 307574 168807 307630 168816
rect 307588 167686 307616 168807
rect 307576 167680 307628 167686
rect 307576 167622 307628 167628
rect 307666 167648 307722 167657
rect 307666 167583 307722 167592
rect 307482 167240 307538 167249
rect 307482 167175 307538 167184
rect 307496 167074 307524 167175
rect 307680 167142 307708 167583
rect 307668 167136 307720 167142
rect 307668 167078 307720 167084
rect 307484 167068 307536 167074
rect 307484 167010 307536 167016
rect 307666 166832 307722 166841
rect 307666 166767 307722 166776
rect 307482 165880 307538 165889
rect 307482 165815 307538 165824
rect 307496 165646 307524 165815
rect 307680 165714 307708 166767
rect 307668 165708 307720 165714
rect 307668 165650 307720 165656
rect 307484 165640 307536 165646
rect 307484 165582 307536 165588
rect 307574 165472 307630 165481
rect 307574 165407 307630 165416
rect 307588 164354 307616 165407
rect 307666 164656 307722 164665
rect 307666 164591 307722 164600
rect 307576 164348 307628 164354
rect 307576 164290 307628 164296
rect 307680 164286 307708 164591
rect 307668 164280 307720 164286
rect 307668 164222 307720 164228
rect 307482 163840 307538 163849
rect 307482 163775 307538 163784
rect 307392 163532 307444 163538
rect 307392 163474 307444 163480
rect 307496 162994 307524 163775
rect 307666 163432 307722 163441
rect 307666 163367 307722 163376
rect 307484 162988 307536 162994
rect 307484 162930 307536 162936
rect 307680 162926 307708 163367
rect 307668 162920 307720 162926
rect 307668 162862 307720 162868
rect 307666 162072 307722 162081
rect 307666 162007 307722 162016
rect 307482 161664 307538 161673
rect 307482 161599 307538 161608
rect 307496 161498 307524 161599
rect 307680 161566 307708 162007
rect 307668 161560 307720 161566
rect 307668 161502 307720 161508
rect 307484 161492 307536 161498
rect 307484 161434 307536 161440
rect 307574 160848 307630 160857
rect 307574 160783 307630 160792
rect 307588 160138 307616 160783
rect 307666 160440 307722 160449
rect 307666 160375 307722 160384
rect 307680 160274 307708 160375
rect 307668 160268 307720 160274
rect 307668 160210 307720 160216
rect 307576 160132 307628 160138
rect 307576 160074 307628 160080
rect 307574 160032 307630 160041
rect 307574 159967 307630 159976
rect 307482 159624 307538 159633
rect 307482 159559 307538 159568
rect 307496 158778 307524 159559
rect 307588 158846 307616 159967
rect 307666 159080 307722 159089
rect 307666 159015 307722 159024
rect 307680 158914 307708 159015
rect 307668 158908 307720 158914
rect 307668 158850 307720 158856
rect 307576 158840 307628 158846
rect 307576 158782 307628 158788
rect 307484 158772 307536 158778
rect 307484 158714 307536 158720
rect 307666 158672 307722 158681
rect 307666 158607 307722 158616
rect 307482 158264 307538 158273
rect 307482 158199 307538 158208
rect 307300 158024 307352 158030
rect 307300 157966 307352 157972
rect 307496 157486 307524 158199
rect 307574 157856 307630 157865
rect 307574 157791 307630 157800
rect 307484 157480 307536 157486
rect 307484 157422 307536 157428
rect 307588 156670 307616 157791
rect 307680 157418 307708 158607
rect 307668 157412 307720 157418
rect 307668 157354 307720 157360
rect 307576 156664 307628 156670
rect 307576 156606 307628 156612
rect 307666 156632 307722 156641
rect 307666 156567 307722 156576
rect 307680 156058 307708 156567
rect 307668 156052 307720 156058
rect 307668 155994 307720 156000
rect 307666 155680 307722 155689
rect 307666 155615 307722 155624
rect 307482 155272 307538 155281
rect 307482 155207 307538 155216
rect 307298 154864 307354 154873
rect 307298 154799 307354 154808
rect 307208 149728 307260 149734
rect 307208 149670 307260 149676
rect 307116 141432 307168 141438
rect 307116 141374 307168 141380
rect 307312 138718 307340 154799
rect 307496 154630 307524 155207
rect 307680 154698 307708 155615
rect 307668 154692 307720 154698
rect 307668 154634 307720 154640
rect 307484 154624 307536 154630
rect 307484 154566 307536 154572
rect 307574 154456 307630 154465
rect 307574 154391 307630 154400
rect 307588 153338 307616 154391
rect 307668 153400 307720 153406
rect 307668 153342 307720 153348
rect 307576 153332 307628 153338
rect 307576 153274 307628 153280
rect 307680 153241 307708 153342
rect 307666 153232 307722 153241
rect 307666 153167 307722 153176
rect 307574 152280 307630 152289
rect 307574 152215 307630 152224
rect 307588 151842 307616 152215
rect 307668 151972 307720 151978
rect 307668 151914 307720 151920
rect 307680 151881 307708 151914
rect 307666 151872 307722 151881
rect 307576 151836 307628 151842
rect 307666 151807 307722 151816
rect 307576 151778 307628 151784
rect 307482 151464 307538 151473
rect 307482 151399 307538 151408
rect 307496 150550 307524 151399
rect 307574 151056 307630 151065
rect 307574 150991 307630 151000
rect 307484 150544 307536 150550
rect 307484 150486 307536 150492
rect 307588 150482 307616 150991
rect 307666 150648 307722 150657
rect 307666 150583 307668 150592
rect 307720 150583 307722 150592
rect 307668 150554 307720 150560
rect 307576 150476 307628 150482
rect 307576 150418 307628 150424
rect 307482 149832 307538 149841
rect 307482 149767 307538 149776
rect 307496 149122 307524 149767
rect 307484 149116 307536 149122
rect 307484 149058 307536 149064
rect 307574 148880 307630 148889
rect 307574 148815 307630 148824
rect 307482 148472 307538 148481
rect 307482 148407 307538 148416
rect 307496 147694 307524 148407
rect 307588 147830 307616 148815
rect 307666 148064 307722 148073
rect 307666 147999 307722 148008
rect 307576 147824 307628 147830
rect 307576 147766 307628 147772
rect 307680 147762 307708 147999
rect 307668 147756 307720 147762
rect 307668 147698 307720 147704
rect 307484 147688 307536 147694
rect 307390 147656 307446 147665
rect 307484 147630 307536 147636
rect 307390 147591 307446 147600
rect 307404 144226 307432 147591
rect 307482 147248 307538 147257
rect 307482 147183 307538 147192
rect 307496 146334 307524 147183
rect 307574 146840 307630 146849
rect 307574 146775 307630 146784
rect 307588 146402 307616 146775
rect 307668 146464 307720 146470
rect 307666 146432 307668 146441
rect 307720 146432 307722 146441
rect 307576 146396 307628 146402
rect 307666 146367 307722 146376
rect 307576 146338 307628 146344
rect 307484 146328 307536 146334
rect 307484 146270 307536 146276
rect 307392 144220 307444 144226
rect 307392 144162 307444 144168
rect 307666 143848 307722 143857
rect 307666 143783 307722 143792
rect 307680 143614 307708 143783
rect 307668 143608 307720 143614
rect 307668 143550 307720 143556
rect 307666 143440 307722 143449
rect 307666 143375 307722 143384
rect 307482 143032 307538 143041
rect 307482 142967 307538 142976
rect 307496 142254 307524 142967
rect 307484 142248 307536 142254
rect 307484 142190 307536 142196
rect 307680 142186 307708 143375
rect 307668 142180 307720 142186
rect 307668 142122 307720 142128
rect 307390 141672 307446 141681
rect 307390 141607 307446 141616
rect 307300 138712 307352 138718
rect 307300 138654 307352 138660
rect 307206 138272 307262 138281
rect 307206 138207 307262 138216
rect 307116 129872 307168 129878
rect 307114 129840 307116 129849
rect 307168 129840 307170 129849
rect 307114 129775 307170 129784
rect 307024 124908 307076 124914
rect 307024 124850 307076 124856
rect 306748 124432 306800 124438
rect 306748 124374 306800 124380
rect 307114 123040 307170 123049
rect 307114 122975 307116 122984
rect 307168 122975 307170 122984
rect 307116 122946 307168 122952
rect 306746 121272 306802 121281
rect 306746 121207 306802 121216
rect 306760 120154 306788 121207
rect 306748 120148 306800 120154
rect 306748 120090 306800 120096
rect 306562 119640 306618 119649
rect 306562 119575 306618 119584
rect 306576 118726 306604 119575
rect 307114 119096 307170 119105
rect 307114 119031 307170 119040
rect 307128 118794 307156 119031
rect 307116 118788 307168 118794
rect 307116 118730 307168 118736
rect 306564 118720 306616 118726
rect 306564 118662 306616 118668
rect 306930 118688 306986 118697
rect 306930 118623 306986 118632
rect 306562 118280 306618 118289
rect 306562 118215 306618 118224
rect 306576 117502 306604 118215
rect 306564 117496 306616 117502
rect 306564 117438 306616 117444
rect 306944 117366 306972 118623
rect 306932 117360 306984 117366
rect 306932 117302 306984 117308
rect 307022 115696 307078 115705
rect 307022 115631 307078 115640
rect 306562 114064 306618 114073
rect 306562 113999 306618 114008
rect 306576 113218 306604 113999
rect 306564 113212 306616 113218
rect 306564 113154 306616 113160
rect 307036 113174 307064 115631
rect 307114 114880 307170 114889
rect 307114 114815 307170 114824
rect 307128 114578 307156 114815
rect 307116 114572 307168 114578
rect 307116 114514 307168 114520
rect 307036 113146 307156 113174
rect 306930 110256 306986 110265
rect 306930 110191 306986 110200
rect 306944 109138 306972 110191
rect 306932 109132 306984 109138
rect 306932 109074 306984 109080
rect 306746 103456 306802 103465
rect 306746 103391 306802 103400
rect 306760 102338 306788 103391
rect 306748 102332 306800 102338
rect 306748 102274 306800 102280
rect 306746 102096 306802 102105
rect 306746 102031 306802 102040
rect 306760 100978 306788 102031
rect 306748 100972 306800 100978
rect 306748 100914 306800 100920
rect 306012 100020 306064 100026
rect 306012 99962 306064 99968
rect 306562 99104 306618 99113
rect 306562 99039 306618 99048
rect 306576 98190 306604 99039
rect 306564 98184 306616 98190
rect 306564 98126 306616 98132
rect 307022 97880 307078 97889
rect 307022 97815 307078 97824
rect 305920 61396 305972 61402
rect 305920 61338 305972 61344
rect 306380 47592 306432 47598
rect 306380 47534 306432 47540
rect 305828 44940 305880 44946
rect 305828 44882 305880 44888
rect 305736 35216 305788 35222
rect 305736 35158 305788 35164
rect 305644 11824 305696 11830
rect 305644 11766 305696 11772
rect 301504 7608 301556 7614
rect 301504 7550 301556 7556
rect 305552 6316 305604 6322
rect 305552 6258 305604 6264
rect 304354 6216 304410 6225
rect 303160 6180 303212 6186
rect 304354 6151 304410 6160
rect 303160 6122 303212 6128
rect 299572 3596 299624 3602
rect 299572 3538 299624 3544
rect 300768 3596 300820 3602
rect 300768 3538 300820 3544
rect 298928 3460 298980 3466
rect 299492 3454 299704 3482
rect 298928 3402 298980 3408
rect 299676 480 299704 3454
rect 300780 480 300808 3538
rect 301964 3460 302016 3466
rect 301964 3402 302016 3408
rect 301976 480 302004 3402
rect 303172 480 303200 6122
rect 304368 480 304396 6151
rect 305564 480 305592 6258
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306392 354 306420 47534
rect 307036 21418 307064 97815
rect 307128 49026 307156 113146
rect 307220 80714 307248 138207
rect 307298 137048 307354 137057
rect 307298 136983 307354 136992
rect 307312 89010 307340 136983
rect 307404 133210 307432 141607
rect 307666 141264 307722 141273
rect 307666 141199 307722 141208
rect 307680 140826 307708 141199
rect 307668 140820 307720 140826
rect 307668 140762 307720 140768
rect 307574 140448 307630 140457
rect 307574 140383 307630 140392
rect 307588 139534 307616 140383
rect 307666 139632 307722 139641
rect 307666 139567 307722 139576
rect 307576 139528 307628 139534
rect 307576 139470 307628 139476
rect 307680 139466 307708 139567
rect 307668 139460 307720 139466
rect 307668 139402 307720 139408
rect 307666 137456 307722 137465
rect 307666 137391 307722 137400
rect 307680 136678 307708 137391
rect 307668 136672 307720 136678
rect 307668 136614 307720 136620
rect 307482 136232 307538 136241
rect 307482 136167 307538 136176
rect 307496 135454 307524 136167
rect 307574 135688 307630 135697
rect 307574 135623 307630 135632
rect 307484 135448 307536 135454
rect 307484 135390 307536 135396
rect 307588 135386 307616 135623
rect 307576 135380 307628 135386
rect 307576 135322 307628 135328
rect 307668 135312 307720 135318
rect 307666 135280 307668 135289
rect 307720 135280 307722 135289
rect 307666 135215 307722 135224
rect 307666 134464 307722 134473
rect 307666 134399 307722 134408
rect 307680 133958 307708 134399
rect 307668 133952 307720 133958
rect 307668 133894 307720 133900
rect 307482 133240 307538 133249
rect 307392 133204 307444 133210
rect 307482 133175 307538 133184
rect 307392 133146 307444 133152
rect 307496 132598 307524 133175
rect 307484 132592 307536 132598
rect 307484 132534 307536 132540
rect 307482 132288 307538 132297
rect 307482 132223 307538 132232
rect 307496 131306 307524 132223
rect 307574 131880 307630 131889
rect 307574 131815 307630 131824
rect 307484 131300 307536 131306
rect 307484 131242 307536 131248
rect 307588 131238 307616 131815
rect 307666 131472 307722 131481
rect 307666 131407 307722 131416
rect 307576 131232 307628 131238
rect 307576 131174 307628 131180
rect 307680 131170 307708 131407
rect 307668 131164 307720 131170
rect 307668 131106 307720 131112
rect 307574 130656 307630 130665
rect 307574 130591 307630 130600
rect 307588 129810 307616 130591
rect 307666 130248 307722 130257
rect 307666 130183 307722 130192
rect 307680 129946 307708 130183
rect 307668 129940 307720 129946
rect 307668 129882 307720 129888
rect 307576 129804 307628 129810
rect 307576 129746 307628 129752
rect 307482 129296 307538 129305
rect 307482 129231 307538 129240
rect 307496 128450 307524 129231
rect 307666 128888 307722 128897
rect 307666 128823 307722 128832
rect 307484 128444 307536 128450
rect 307484 128386 307536 128392
rect 307680 128382 307708 128823
rect 307668 128376 307720 128382
rect 307668 128318 307720 128324
rect 307482 128072 307538 128081
rect 307482 128007 307538 128016
rect 307496 127090 307524 128007
rect 307666 127664 307722 127673
rect 307666 127599 307722 127608
rect 307574 127256 307630 127265
rect 307574 127191 307630 127200
rect 307484 127084 307536 127090
rect 307484 127026 307536 127032
rect 307588 127022 307616 127191
rect 307680 127158 307708 127599
rect 307668 127152 307720 127158
rect 307668 127094 307720 127100
rect 307576 127016 307628 127022
rect 307576 126958 307628 126964
rect 307574 126440 307630 126449
rect 307574 126375 307630 126384
rect 307588 125730 307616 126375
rect 307666 125896 307722 125905
rect 307666 125831 307722 125840
rect 307576 125724 307628 125730
rect 307576 125666 307628 125672
rect 307680 125662 307708 125831
rect 307668 125656 307720 125662
rect 307668 125598 307720 125604
rect 307482 125080 307538 125089
rect 307482 125015 307538 125024
rect 307496 124370 307524 125015
rect 307484 124364 307536 124370
rect 307484 124306 307536 124312
rect 307668 124296 307720 124302
rect 307666 124264 307668 124273
rect 307720 124264 307722 124273
rect 307666 124199 307722 124208
rect 307482 123856 307538 123865
rect 307482 123791 307538 123800
rect 307496 122874 307524 123791
rect 307666 123448 307722 123457
rect 307666 123383 307722 123392
rect 307680 122942 307708 123383
rect 307668 122936 307720 122942
rect 307668 122878 307720 122884
rect 307484 122868 307536 122874
rect 307484 122810 307536 122816
rect 307482 122496 307538 122505
rect 307482 122431 307538 122440
rect 307496 121514 307524 122431
rect 307574 122088 307630 122097
rect 307574 122023 307630 122032
rect 307588 121582 307616 122023
rect 307666 121680 307722 121689
rect 307666 121615 307668 121624
rect 307720 121615 307722 121624
rect 307668 121586 307720 121592
rect 307576 121576 307628 121582
rect 307576 121518 307628 121524
rect 307484 121508 307536 121514
rect 307484 121450 307536 121456
rect 307574 120864 307630 120873
rect 307574 120799 307630 120808
rect 307588 120290 307616 120799
rect 307666 120456 307722 120465
rect 307666 120391 307722 120400
rect 307576 120284 307628 120290
rect 307576 120226 307628 120232
rect 307680 120222 307708 120391
rect 307668 120216 307720 120222
rect 307668 120158 307720 120164
rect 307666 120048 307722 120057
rect 307666 119983 307722 119992
rect 307680 118862 307708 119983
rect 307668 118856 307720 118862
rect 307668 118798 307720 118804
rect 307666 117464 307722 117473
rect 307666 117399 307668 117408
rect 307720 117399 307722 117408
rect 307668 117370 307720 117376
rect 307574 117056 307630 117065
rect 307574 116991 307630 117000
rect 307482 116648 307538 116657
rect 307482 116583 307538 116592
rect 307496 116006 307524 116583
rect 307588 116142 307616 116991
rect 307666 116240 307722 116249
rect 307666 116175 307722 116184
rect 307576 116136 307628 116142
rect 307576 116078 307628 116084
rect 307680 116074 307708 116175
rect 307668 116068 307720 116074
rect 307668 116010 307720 116016
rect 307484 116000 307536 116006
rect 307484 115942 307536 115948
rect 307482 115288 307538 115297
rect 307482 115223 307538 115232
rect 307496 114646 307524 115223
rect 307484 114640 307536 114646
rect 307484 114582 307536 114588
rect 307574 114472 307630 114481
rect 307574 114407 307630 114416
rect 307588 113286 307616 114407
rect 307668 113348 307720 113354
rect 307668 113290 307720 113296
rect 307576 113280 307628 113286
rect 307680 113257 307708 113290
rect 307576 113222 307628 113228
rect 307666 113248 307722 113257
rect 307666 113183 307722 113192
rect 307574 112296 307630 112305
rect 307574 112231 307630 112240
rect 307588 111926 307616 112231
rect 307576 111920 307628 111926
rect 307576 111862 307628 111868
rect 307666 111888 307722 111897
rect 307666 111823 307668 111832
rect 307720 111823 307722 111832
rect 307668 111794 307720 111800
rect 307482 111480 307538 111489
rect 307482 111415 307538 111424
rect 307496 110566 307524 111415
rect 307666 111072 307722 111081
rect 307666 111007 307722 111016
rect 307574 110664 307630 110673
rect 307680 110634 307708 111007
rect 307574 110599 307630 110608
rect 307668 110628 307720 110634
rect 307484 110560 307536 110566
rect 307484 110502 307536 110508
rect 307588 110498 307616 110599
rect 307668 110570 307720 110576
rect 307576 110492 307628 110498
rect 307576 110434 307628 110440
rect 307666 109848 307722 109857
rect 307666 109783 307722 109792
rect 307574 109304 307630 109313
rect 307574 109239 307630 109248
rect 307588 109070 307616 109239
rect 307680 109206 307708 109783
rect 307668 109200 307720 109206
rect 307668 109142 307720 109148
rect 307576 109064 307628 109070
rect 307576 109006 307628 109012
rect 307390 108896 307446 108905
rect 307390 108831 307446 108840
rect 307404 107778 307432 108831
rect 307482 108488 307538 108497
rect 307482 108423 307538 108432
rect 307392 107772 307444 107778
rect 307392 107714 307444 107720
rect 307496 107710 307524 108423
rect 307666 108080 307722 108089
rect 307666 108015 307722 108024
rect 307680 107914 307708 108015
rect 307668 107908 307720 107914
rect 307668 107850 307720 107856
rect 307576 107840 307628 107846
rect 307576 107782 307628 107788
rect 307484 107704 307536 107710
rect 307588 107681 307616 107782
rect 307484 107646 307536 107652
rect 307574 107672 307630 107681
rect 307574 107607 307630 107616
rect 307482 107264 307538 107273
rect 307482 107199 307538 107208
rect 307496 106321 307524 107199
rect 307574 106856 307630 106865
rect 307574 106791 307630 106800
rect 307588 106418 307616 106791
rect 307668 106480 307720 106486
rect 307666 106448 307668 106457
rect 307720 106448 307722 106457
rect 307576 106412 307628 106418
rect 307666 106383 307722 106392
rect 307576 106354 307628 106360
rect 307482 106312 307538 106321
rect 307482 106247 307538 106256
rect 307574 105496 307630 105505
rect 307574 105431 307630 105440
rect 307588 104990 307616 105431
rect 307666 105088 307722 105097
rect 307666 105023 307722 105032
rect 307576 104984 307628 104990
rect 307576 104926 307628 104932
rect 307680 104922 307708 105023
rect 307668 104916 307720 104922
rect 307668 104858 307720 104864
rect 307482 104680 307538 104689
rect 307482 104615 307538 104624
rect 307496 103698 307524 104615
rect 307666 104272 307722 104281
rect 307666 104207 307722 104216
rect 307484 103692 307536 103698
rect 307484 103634 307536 103640
rect 307680 103630 307708 104207
rect 307668 103624 307720 103630
rect 307668 103566 307720 103572
rect 307482 103048 307538 103057
rect 307482 102983 307538 102992
rect 307496 102270 307524 102983
rect 307666 102504 307722 102513
rect 307666 102439 307722 102448
rect 307484 102264 307536 102270
rect 307484 102206 307536 102212
rect 307680 102202 307708 102439
rect 307668 102196 307720 102202
rect 307668 102138 307720 102144
rect 307482 101688 307538 101697
rect 307482 101623 307538 101632
rect 307496 100910 307524 101623
rect 307574 101280 307630 101289
rect 307574 101215 307630 101224
rect 307484 100904 307536 100910
rect 307484 100846 307536 100852
rect 307588 100774 307616 101215
rect 307666 100872 307722 100881
rect 307666 100807 307668 100816
rect 307720 100807 307722 100816
rect 307668 100778 307720 100784
rect 307576 100768 307628 100774
rect 307576 100710 307628 100716
rect 307666 100464 307722 100473
rect 307666 100399 307722 100408
rect 307482 100056 307538 100065
rect 307482 99991 307538 100000
rect 307496 99414 307524 99991
rect 307680 99521 307708 100399
rect 307666 99512 307722 99521
rect 307666 99447 307722 99456
rect 307484 99408 307536 99414
rect 307484 99350 307536 99356
rect 307574 98696 307630 98705
rect 307574 98631 307630 98640
rect 307588 98122 307616 98631
rect 307666 98288 307722 98297
rect 307666 98223 307722 98232
rect 307576 98116 307628 98122
rect 307576 98058 307628 98064
rect 307680 98054 307708 98223
rect 307668 98048 307720 98054
rect 307668 97990 307720 97996
rect 307482 97472 307538 97481
rect 307482 97407 307538 97416
rect 307496 96694 307524 97407
rect 307668 96756 307720 96762
rect 307668 96698 307720 96704
rect 307484 96688 307536 96694
rect 307680 96665 307708 96698
rect 307484 96630 307536 96636
rect 307666 96656 307722 96665
rect 307666 96591 307722 96600
rect 307666 96248 307722 96257
rect 307666 96183 307722 96192
rect 307680 95266 307708 96183
rect 307668 95260 307720 95266
rect 307668 95202 307720 95208
rect 307300 89004 307352 89010
rect 307300 88946 307352 88952
rect 307208 80708 307260 80714
rect 307208 80650 307260 80656
rect 307116 49020 307168 49026
rect 307116 48962 307168 48968
rect 307024 21412 307076 21418
rect 307024 21354 307076 21360
rect 307772 16574 307800 356662
rect 308404 339516 308456 339522
rect 308404 339458 308456 339464
rect 308416 90370 308444 339458
rect 309152 231742 309180 700334
rect 309784 354884 309836 354890
rect 309784 354826 309836 354832
rect 309140 231736 309192 231742
rect 309140 231678 309192 231684
rect 308496 205148 308548 205154
rect 308496 205090 308548 205096
rect 308404 90364 308456 90370
rect 308404 90306 308456 90312
rect 307772 16546 307984 16574
rect 307956 480 307984 16546
rect 308508 2990 308536 205090
rect 309048 6316 309100 6322
rect 309048 6258 309100 6264
rect 308496 2984 308548 2990
rect 308496 2926 308548 2932
rect 309060 480 309088 6258
rect 309796 3398 309824 354826
rect 310532 235618 310560 700402
rect 331232 374678 331260 702986
rect 348804 696250 348832 703520
rect 364996 700398 365024 703520
rect 354588 700392 354640 700398
rect 354588 700334 354640 700340
rect 364984 700392 365036 700398
rect 364984 700334 365036 700340
rect 383568 700392 383620 700398
rect 383568 700334 383620 700340
rect 348792 696244 348844 696250
rect 348792 696186 348844 696192
rect 331220 374672 331272 374678
rect 331220 374614 331272 374620
rect 313924 371340 313976 371346
rect 313924 371282 313976 371288
rect 311900 354816 311952 354822
rect 311900 354758 311952 354764
rect 310612 305040 310664 305046
rect 310612 304982 310664 304988
rect 310520 235612 310572 235618
rect 310520 235554 310572 235560
rect 310428 222080 310480 222086
rect 310428 222022 310480 222028
rect 310440 221474 310468 222022
rect 310428 221468 310480 221474
rect 310428 221410 310480 221416
rect 309876 202360 309928 202366
rect 309876 202302 309928 202308
rect 309784 3392 309836 3398
rect 309784 3334 309836 3340
rect 309888 3330 309916 202302
rect 310440 180033 310468 221410
rect 310624 216617 310652 304982
rect 311164 233912 311216 233918
rect 311164 233854 311216 233860
rect 310610 216608 310666 216617
rect 310610 216543 310666 216552
rect 310624 215393 310652 216543
rect 310610 215384 310666 215393
rect 310610 215319 310666 215328
rect 311176 181694 311204 233854
rect 311912 217462 311940 354758
rect 313280 307828 313332 307834
rect 313280 307770 313332 307776
rect 313292 239873 313320 307770
rect 313278 239864 313334 239873
rect 313278 239799 313334 239808
rect 311900 217456 311952 217462
rect 311900 217398 311952 217404
rect 311254 215384 311310 215393
rect 311254 215319 311310 215328
rect 311164 181688 311216 181694
rect 311164 181630 311216 181636
rect 310426 180024 310482 180033
rect 310426 179959 310482 179968
rect 311268 177546 311296 215319
rect 312544 211812 312596 211818
rect 312544 211754 312596 211760
rect 311256 177540 311308 177546
rect 311256 177482 311308 177488
rect 312556 176118 312584 211754
rect 313936 177313 313964 371282
rect 340880 367328 340932 367334
rect 340880 367270 340932 367276
rect 331220 364540 331272 364546
rect 331220 364482 331272 364488
rect 318064 363180 318116 363186
rect 318064 363122 318116 363128
rect 315304 361888 315356 361894
rect 315304 361830 315356 361836
rect 314016 278044 314068 278050
rect 314016 277986 314068 277992
rect 314028 222086 314056 277986
rect 314016 222080 314068 222086
rect 314016 222022 314068 222028
rect 314016 215960 314068 215966
rect 314016 215902 314068 215908
rect 314028 177614 314056 215902
rect 315316 203726 315344 361830
rect 316038 352608 316094 352617
rect 316038 352543 316094 352552
rect 315396 231124 315448 231130
rect 315396 231066 315448 231072
rect 315304 203720 315356 203726
rect 315304 203662 315356 203668
rect 315408 180334 315436 231066
rect 316052 225622 316080 352543
rect 316040 225616 316092 225622
rect 316040 225558 316092 225564
rect 315488 206372 315540 206378
rect 315488 206314 315540 206320
rect 315396 180328 315448 180334
rect 315396 180270 315448 180276
rect 314016 177608 314068 177614
rect 314016 177550 314068 177556
rect 313922 177304 313978 177313
rect 313922 177239 313978 177248
rect 312544 176112 312596 176118
rect 312544 176054 312596 176060
rect 315500 175953 315528 206314
rect 318076 199646 318104 363122
rect 319444 361820 319496 361826
rect 319444 361762 319496 361768
rect 318156 289944 318208 289950
rect 318156 289886 318208 289892
rect 318168 227662 318196 289886
rect 318156 227656 318208 227662
rect 318156 227598 318208 227604
rect 318064 199640 318116 199646
rect 318064 199582 318116 199588
rect 318156 199572 318208 199578
rect 318156 199514 318208 199520
rect 318064 184204 318116 184210
rect 318064 184146 318116 184152
rect 317328 178832 317380 178838
rect 317328 178774 317380 178780
rect 317340 178129 317368 178774
rect 318076 178566 318104 184146
rect 318064 178560 318116 178566
rect 318064 178502 318116 178508
rect 316038 178120 316094 178129
rect 316038 178055 316094 178064
rect 317326 178120 317382 178129
rect 317326 178055 317382 178064
rect 315486 175944 315542 175953
rect 316052 175930 316080 178055
rect 318168 176089 318196 199514
rect 319456 195265 319484 361762
rect 329196 360528 329248 360534
rect 329196 360470 329248 360476
rect 324962 357776 325018 357785
rect 324962 357711 325018 357720
rect 323584 320204 323636 320210
rect 323584 320146 323636 320152
rect 319536 292596 319588 292602
rect 319536 292538 319588 292544
rect 319548 237114 319576 292538
rect 319536 237108 319588 237114
rect 319536 237050 319588 237056
rect 323596 211818 323624 320146
rect 323676 291236 323728 291242
rect 323676 291178 323728 291184
rect 323688 235822 323716 291178
rect 323676 235816 323728 235822
rect 323676 235758 323728 235764
rect 323584 211812 323636 211818
rect 323584 211754 323636 211760
rect 322940 200796 322992 200802
rect 322940 200738 322992 200744
rect 319536 196784 319588 196790
rect 319536 196726 319588 196732
rect 319442 195256 319498 195265
rect 319442 195191 319498 195200
rect 319548 176186 319576 196726
rect 320824 196648 320876 196654
rect 320824 196590 320876 196596
rect 320836 190454 320864 196590
rect 321652 193860 321704 193866
rect 321652 193802 321704 193808
rect 321560 191140 321612 191146
rect 321560 191082 321612 191088
rect 320836 190426 321324 190454
rect 320180 186992 320232 186998
rect 320180 186934 320232 186940
rect 320192 176769 320220 186934
rect 320178 176760 320234 176769
rect 320178 176695 320234 176704
rect 319536 176180 319588 176186
rect 319536 176122 319588 176128
rect 318154 176080 318210 176089
rect 318154 176015 318210 176024
rect 316020 175902 316080 175930
rect 315486 175879 315542 175888
rect 321296 165753 321324 190426
rect 321282 165744 321338 165753
rect 321282 165679 321338 165688
rect 321572 106865 321600 191082
rect 321664 122806 321692 193802
rect 321836 184272 321888 184278
rect 321836 184214 321888 184220
rect 321744 180124 321796 180130
rect 321744 180066 321796 180072
rect 321756 139097 321784 180066
rect 321848 148345 321876 184214
rect 321834 148336 321890 148345
rect 321834 148271 321890 148280
rect 322846 147792 322902 147801
rect 322846 147727 322902 147736
rect 322860 147694 322888 147727
rect 322848 147688 322900 147694
rect 322848 147630 322900 147636
rect 321742 139088 321798 139097
rect 321742 139023 321798 139032
rect 322846 138544 322902 138553
rect 322846 138479 322902 138488
rect 322860 138038 322888 138479
rect 322848 138032 322900 138038
rect 322848 137974 322900 137980
rect 321652 122800 321704 122806
rect 321652 122742 321704 122748
rect 321664 122233 321692 122742
rect 321650 122224 321706 122233
rect 321650 122159 321706 122168
rect 321558 106856 321614 106865
rect 321558 106791 321614 106800
rect 321742 106856 321798 106865
rect 321742 106791 321798 106800
rect 321572 106350 321600 106791
rect 321560 106344 321612 106350
rect 321560 106286 321612 106292
rect 321650 101144 321706 101153
rect 321650 101079 321706 101088
rect 321558 96656 321614 96665
rect 321558 96591 321614 96600
rect 321572 95169 321600 96591
rect 321558 95160 321614 95169
rect 321558 95095 321614 95104
rect 317420 90364 317472 90370
rect 317420 90306 317472 90312
rect 311900 77988 311952 77994
rect 311900 77930 311952 77936
rect 311912 16574 311940 77930
rect 316132 68468 316184 68474
rect 316132 68410 316184 68416
rect 313278 50280 313334 50289
rect 313278 50215 313334 50224
rect 313292 16574 313320 50215
rect 316144 16574 316172 68410
rect 317432 16574 317460 90306
rect 321664 84194 321692 101079
rect 321756 96626 321784 106791
rect 322952 104009 322980 200738
rect 323124 185700 323176 185706
rect 323124 185642 323176 185648
rect 323032 178560 323084 178566
rect 323032 178502 323084 178508
rect 323044 129441 323072 178502
rect 323136 164801 323164 185642
rect 323688 185065 323716 235758
rect 324320 203584 324372 203590
rect 324320 203526 324372 203532
rect 324332 186314 324360 203526
rect 324412 191344 324464 191350
rect 324412 191286 324464 191292
rect 324424 190466 324452 191286
rect 324976 191146 325004 357711
rect 325056 318844 325108 318850
rect 325056 318786 325108 318792
rect 325068 271182 325096 318786
rect 327724 296744 327776 296750
rect 327724 296686 327776 296692
rect 326344 280220 326396 280226
rect 326344 280162 326396 280168
rect 325056 271176 325108 271182
rect 325056 271118 325108 271124
rect 325056 269136 325108 269142
rect 325056 269078 325108 269084
rect 325068 214742 325096 269078
rect 326356 233170 326384 280162
rect 325700 233164 325752 233170
rect 325700 233106 325752 233112
rect 326344 233164 326396 233170
rect 326344 233106 326396 233112
rect 325056 214736 325108 214742
rect 325056 214678 325108 214684
rect 324964 191140 325016 191146
rect 324964 191082 325016 191088
rect 324412 190460 324464 190466
rect 324412 190402 324464 190408
rect 324424 189145 324452 190402
rect 324504 189848 324556 189854
rect 324504 189790 324556 189796
rect 324410 189136 324466 189145
rect 324410 189071 324466 189080
rect 324516 189038 324544 189790
rect 324504 189032 324556 189038
rect 324504 188974 324556 188980
rect 325056 189032 325108 189038
rect 325056 188974 325108 188980
rect 324332 186286 324728 186314
rect 324504 185632 324556 185638
rect 324504 185574 324556 185580
rect 323674 185056 323730 185065
rect 323674 184991 323730 185000
rect 324320 176656 324372 176662
rect 324320 176598 324372 176604
rect 324332 175545 324360 176598
rect 324318 175536 324374 175545
rect 324318 175471 324374 175480
rect 324320 175228 324372 175234
rect 324320 175170 324372 175176
rect 324332 174049 324360 175170
rect 324318 174040 324374 174049
rect 324318 173975 324374 173984
rect 324320 172508 324372 172514
rect 324320 172450 324372 172456
rect 324332 171737 324360 172450
rect 324318 171728 324374 171737
rect 324318 171663 324374 171672
rect 324320 171080 324372 171086
rect 324320 171022 324372 171028
rect 324332 170921 324360 171022
rect 324318 170912 324374 170921
rect 324318 170847 324374 170856
rect 324318 170096 324374 170105
rect 324318 170031 324374 170040
rect 324332 169794 324360 170031
rect 324320 169788 324372 169794
rect 324320 169730 324372 169736
rect 324516 169726 324544 185574
rect 324504 169720 324556 169726
rect 324504 169662 324556 169668
rect 324318 169416 324374 169425
rect 324318 169351 324374 169360
rect 324332 169046 324360 169351
rect 324320 169040 324372 169046
rect 324320 168982 324372 168988
rect 324516 168609 324544 169662
rect 324502 168600 324558 168609
rect 324502 168535 324558 168544
rect 324320 168360 324372 168366
rect 324320 168302 324372 168308
rect 324332 167113 324360 168302
rect 324700 168298 324728 186286
rect 324964 185836 325016 185842
rect 324964 185778 325016 185784
rect 324870 172136 324926 172145
rect 324870 172071 324926 172080
rect 324884 171154 324912 172071
rect 324872 171148 324924 171154
rect 324872 171090 324924 171096
rect 324412 168292 324464 168298
rect 324412 168234 324464 168240
rect 324688 168292 324740 168298
rect 324688 168234 324740 168240
rect 324424 167793 324452 168234
rect 324410 167784 324466 167793
rect 324410 167719 324466 167728
rect 324318 167104 324374 167113
rect 324318 167039 324374 167048
rect 324320 167000 324372 167006
rect 324320 166942 324372 166948
rect 324332 166297 324360 166942
rect 324318 166288 324374 166297
rect 324318 166223 324374 166232
rect 324318 165472 324374 165481
rect 324318 165407 324374 165416
rect 323122 164792 323178 164801
rect 323122 164727 323178 164736
rect 323398 164792 323454 164801
rect 323398 164727 323454 164736
rect 323412 164286 323440 164727
rect 324332 164354 324360 165407
rect 324320 164348 324372 164354
rect 324320 164290 324372 164296
rect 323400 164280 323452 164286
rect 323400 164222 323452 164228
rect 324320 164212 324372 164218
rect 324320 164154 324372 164160
rect 324332 163985 324360 164154
rect 324412 164144 324464 164150
rect 324412 164086 324464 164092
rect 324318 163976 324374 163985
rect 324318 163911 324374 163920
rect 324424 163169 324452 164086
rect 324410 163160 324466 163169
rect 324410 163095 324466 163104
rect 324318 160848 324374 160857
rect 324318 160783 324374 160792
rect 324332 160750 324360 160783
rect 324320 160744 324372 160750
rect 324320 160686 324372 160692
rect 324320 159384 324372 159390
rect 324318 159352 324320 159361
rect 324372 159352 324374 159361
rect 324318 159287 324374 159296
rect 324412 158704 324464 158710
rect 324412 158646 324464 158652
rect 324320 158636 324372 158642
rect 324320 158578 324372 158584
rect 324332 158545 324360 158578
rect 324318 158536 324374 158545
rect 324318 158471 324374 158480
rect 324424 157865 324452 158646
rect 324410 157856 324466 157865
rect 324410 157791 324466 157800
rect 324320 157344 324372 157350
rect 324320 157286 324372 157292
rect 324332 157049 324360 157286
rect 324412 157276 324464 157282
rect 324412 157218 324464 157224
rect 324318 157040 324374 157049
rect 324318 156975 324374 156984
rect 324424 156369 324452 157218
rect 324410 156360 324466 156369
rect 324410 156295 324466 156304
rect 324320 155916 324372 155922
rect 324320 155858 324372 155864
rect 324332 154737 324360 155858
rect 324318 154728 324374 154737
rect 324318 154663 324374 154672
rect 324320 154556 324372 154562
rect 324320 154498 324372 154504
rect 324332 154057 324360 154498
rect 324412 154488 324464 154494
rect 324412 154430 324464 154436
rect 324318 154048 324374 154057
rect 324318 153983 324374 153992
rect 324424 153241 324452 154430
rect 324976 153270 325004 185778
rect 325068 174729 325096 188974
rect 325054 174720 325110 174729
rect 325054 174655 325110 174664
rect 325606 160168 325662 160177
rect 325712 160154 325740 233106
rect 327736 230382 327764 296686
rect 328460 267096 328512 267102
rect 328460 267038 328512 267044
rect 327816 252612 327868 252618
rect 327816 252554 327868 252560
rect 327724 230376 327776 230382
rect 327724 230318 327776 230324
rect 327828 223582 327856 252554
rect 327172 223576 327224 223582
rect 327172 223518 327224 223524
rect 327816 223576 327868 223582
rect 327816 223518 327868 223524
rect 327080 209228 327132 209234
rect 327080 209170 327132 209176
rect 325792 178764 325844 178770
rect 325792 178706 325844 178712
rect 325662 160126 325740 160154
rect 325606 160103 325662 160112
rect 324964 153264 325016 153270
rect 324410 153232 324466 153241
rect 324964 153206 325016 153212
rect 324410 153167 324466 153176
rect 324976 152425 325004 153206
rect 324962 152416 325018 152425
rect 324962 152351 325018 152360
rect 324320 151768 324372 151774
rect 324320 151710 324372 151716
rect 324410 151736 324466 151745
rect 324332 150929 324360 151710
rect 324410 151671 324466 151680
rect 324318 150920 324374 150929
rect 324318 150855 324374 150864
rect 324424 150482 324452 151671
rect 324412 150476 324464 150482
rect 324412 150418 324464 150424
rect 324320 150408 324372 150414
rect 324320 150350 324372 150356
rect 324332 150113 324360 150350
rect 324412 150340 324464 150346
rect 324412 150282 324464 150288
rect 324318 150104 324374 150113
rect 324318 150039 324374 150048
rect 324424 149433 324452 150282
rect 324410 149424 324466 149433
rect 324410 149359 324466 149368
rect 324320 147620 324372 147626
rect 324320 147562 324372 147568
rect 324332 147121 324360 147562
rect 324318 147112 324374 147121
rect 324318 147047 324374 147056
rect 324320 145580 324372 145586
rect 324320 145522 324372 145528
rect 324332 145489 324360 145522
rect 324318 145480 324374 145489
rect 324318 145415 324374 145424
rect 324412 144900 324464 144906
rect 324412 144842 324464 144848
rect 324320 144832 324372 144838
rect 324318 144800 324320 144809
rect 324372 144800 324374 144809
rect 324318 144735 324374 144744
rect 324424 143993 324452 144842
rect 324410 143984 324466 143993
rect 324410 143919 324466 143928
rect 324412 143540 324464 143546
rect 324412 143482 324464 143488
rect 324320 143404 324372 143410
rect 324320 143346 324372 143352
rect 324332 143177 324360 143346
rect 324318 143168 324374 143177
rect 324318 143103 324374 143112
rect 324424 142497 324452 143482
rect 324410 142488 324466 142497
rect 324410 142423 324466 142432
rect 324412 142112 324464 142118
rect 324412 142054 324464 142060
rect 324320 142044 324372 142050
rect 324320 141986 324372 141992
rect 324332 141681 324360 141986
rect 324318 141672 324374 141681
rect 324318 141607 324374 141616
rect 324424 140865 324452 142054
rect 324410 140856 324466 140865
rect 324410 140791 324466 140800
rect 324320 140752 324372 140758
rect 324320 140694 324372 140700
rect 324332 140185 324360 140694
rect 324318 140176 324374 140185
rect 324318 140111 324374 140120
rect 324320 137964 324372 137970
rect 324320 137906 324372 137912
rect 324332 137873 324360 137906
rect 324412 137896 324464 137902
rect 324318 137864 324374 137873
rect 324412 137838 324464 137844
rect 324318 137799 324374 137808
rect 324424 137057 324452 137838
rect 324410 137048 324466 137057
rect 324410 136983 324466 136992
rect 324320 136604 324372 136610
rect 324320 136546 324372 136552
rect 324332 136377 324360 136546
rect 324412 136536 324464 136542
rect 324412 136478 324464 136484
rect 324318 136368 324374 136377
rect 324318 136303 324374 136312
rect 324424 135561 324452 136478
rect 324410 135552 324466 135561
rect 324410 135487 324466 135496
rect 324320 135244 324372 135250
rect 324320 135186 324372 135192
rect 324332 134745 324360 135186
rect 324412 135176 324464 135182
rect 324412 135118 324464 135124
rect 324318 134736 324374 134745
rect 324318 134671 324374 134680
rect 324424 134065 324452 135118
rect 325516 134564 325568 134570
rect 325516 134506 325568 134512
rect 324410 134056 324466 134065
rect 324410 133991 324466 134000
rect 324320 133884 324372 133890
rect 324320 133826 324372 133832
rect 324332 133249 324360 133826
rect 324318 133240 324374 133249
rect 324318 133175 324374 133184
rect 324320 132456 324372 132462
rect 324318 132424 324320 132433
rect 324372 132424 324374 132433
rect 324318 132359 324374 132368
rect 324412 132388 324464 132394
rect 324412 132330 324464 132336
rect 324424 131753 324452 132330
rect 324410 131744 324466 131753
rect 324410 131679 324466 131688
rect 324412 131096 324464 131102
rect 324412 131038 324464 131044
rect 324320 131028 324372 131034
rect 324320 130970 324372 130976
rect 324332 130937 324360 130970
rect 324318 130928 324374 130937
rect 324318 130863 324374 130872
rect 324424 130121 324452 131038
rect 324410 130112 324466 130121
rect 324410 130047 324466 130056
rect 323030 129432 323086 129441
rect 323030 129367 323086 129376
rect 325054 129432 325110 129441
rect 325054 129367 325110 129376
rect 324320 129056 324372 129062
rect 324320 128998 324372 129004
rect 324332 128625 324360 128998
rect 324318 128616 324374 128625
rect 324318 128551 324374 128560
rect 324320 128308 324372 128314
rect 324320 128250 324372 128256
rect 324332 127809 324360 128250
rect 324318 127800 324374 127809
rect 324318 127735 324374 127744
rect 324502 127120 324558 127129
rect 324502 127055 324558 127064
rect 324320 126948 324372 126954
rect 324320 126890 324372 126896
rect 324332 126313 324360 126890
rect 324318 126304 324374 126313
rect 324318 126239 324374 126248
rect 324320 125588 324372 125594
rect 324320 125530 324372 125536
rect 324332 125497 324360 125530
rect 324412 125520 324464 125526
rect 324318 125488 324374 125497
rect 324412 125462 324464 125468
rect 324318 125423 324374 125432
rect 324424 124817 324452 125462
rect 324410 124808 324466 124817
rect 324410 124743 324466 124752
rect 324516 124166 324544 127055
rect 324504 124160 324556 124166
rect 324504 124102 324556 124108
rect 324320 124092 324372 124098
rect 324320 124034 324372 124040
rect 324332 124001 324360 124034
rect 324412 124024 324464 124030
rect 324318 123992 324374 124001
rect 324412 123966 324464 123972
rect 324318 123927 324374 123936
rect 324424 123185 324452 123966
rect 324410 123176 324466 123185
rect 324410 123111 324466 123120
rect 324320 122528 324372 122534
rect 324318 122496 324320 122505
rect 324372 122496 324374 122505
rect 324318 122431 324374 122440
rect 324320 121440 324372 121446
rect 324320 121382 324372 121388
rect 324332 120873 324360 121382
rect 324412 121372 324464 121378
rect 324412 121314 324464 121320
rect 324318 120864 324374 120873
rect 324318 120799 324374 120808
rect 324424 120193 324452 121314
rect 324410 120184 324466 120193
rect 324410 120119 324466 120128
rect 324320 120080 324372 120086
rect 324320 120022 324372 120028
rect 324332 119377 324360 120022
rect 324318 119368 324374 119377
rect 324318 119303 324374 119312
rect 324412 118652 324464 118658
rect 324412 118594 324464 118600
rect 324320 118584 324372 118590
rect 324318 118552 324320 118561
rect 324372 118552 324374 118561
rect 324318 118487 324374 118496
rect 324424 117881 324452 118594
rect 324504 117972 324556 117978
rect 324504 117914 324556 117920
rect 324410 117872 324466 117881
rect 324410 117807 324466 117816
rect 324320 117292 324372 117298
rect 324320 117234 324372 117240
rect 324332 117065 324360 117234
rect 324318 117056 324374 117065
rect 324318 116991 324374 117000
rect 324516 116385 324544 117914
rect 324502 116376 324558 116385
rect 324502 116311 324558 116320
rect 324412 115932 324464 115938
rect 324412 115874 324464 115880
rect 324318 115560 324374 115569
rect 324318 115495 324374 115504
rect 324332 115122 324360 115495
rect 324320 115116 324372 115122
rect 324320 115058 324372 115064
rect 324424 114753 324452 115874
rect 324780 115252 324832 115258
rect 324780 115194 324832 115200
rect 324410 114744 324466 114753
rect 324410 114679 324466 114688
rect 324412 114504 324464 114510
rect 324412 114446 324464 114452
rect 324320 114436 324372 114442
rect 324320 114378 324372 114384
rect 324332 114073 324360 114378
rect 324318 114064 324374 114073
rect 324318 113999 324374 114008
rect 324424 113257 324452 114446
rect 324410 113248 324466 113257
rect 324410 113183 324466 113192
rect 324320 113144 324372 113150
rect 324320 113086 324372 113092
rect 324332 112441 324360 113086
rect 324318 112432 324374 112441
rect 324318 112367 324374 112376
rect 324320 111784 324372 111790
rect 324320 111726 324372 111732
rect 324410 111752 324466 111761
rect 324332 110945 324360 111726
rect 324410 111687 324466 111696
rect 324318 110936 324374 110945
rect 324318 110871 324374 110880
rect 324424 110770 324452 111687
rect 324412 110764 324464 110770
rect 324412 110706 324464 110712
rect 324320 110424 324372 110430
rect 324320 110366 324372 110372
rect 324332 109449 324360 110366
rect 324792 110129 324820 115194
rect 325068 112470 325096 129367
rect 325056 112464 325108 112470
rect 325056 112406 325108 112412
rect 324778 110120 324834 110129
rect 324778 110055 324834 110064
rect 324318 109440 324374 109449
rect 324318 109375 324374 109384
rect 324410 108624 324466 108633
rect 324410 108559 324466 108568
rect 324320 108384 324372 108390
rect 324320 108326 324372 108332
rect 324332 107817 324360 108326
rect 324424 108322 324452 108559
rect 324412 108316 324464 108322
rect 324412 108258 324464 108264
rect 324318 107808 324374 107817
rect 324318 107743 324374 107752
rect 324320 106276 324372 106282
rect 324320 106218 324372 106224
rect 324332 105505 324360 106218
rect 324318 105496 324374 105505
rect 324318 105431 324374 105440
rect 324424 105346 324452 108258
rect 325528 107137 325556 134506
rect 325804 108390 325832 178706
rect 326434 178664 326490 178673
rect 326434 178599 326490 178608
rect 326448 178022 326476 178599
rect 326436 178016 326488 178022
rect 326436 177958 326488 177964
rect 325884 177336 325936 177342
rect 325884 177278 325936 177284
rect 325896 162178 325924 177278
rect 325884 162172 325936 162178
rect 325884 162114 325936 162120
rect 325896 161673 325924 162114
rect 325882 161664 325938 161673
rect 325882 161599 325938 161608
rect 326448 161474 326476 177958
rect 326356 161446 326476 161474
rect 326356 143410 326384 161446
rect 326344 143404 326396 143410
rect 326344 143346 326396 143352
rect 327092 122534 327120 209170
rect 327184 144838 327212 223518
rect 327908 209228 327960 209234
rect 327908 209170 327960 209176
rect 327920 208418 327948 209170
rect 327908 208412 327960 208418
rect 327908 208354 327960 208360
rect 327264 187060 327316 187066
rect 327264 187002 327316 187008
rect 327276 169046 327304 187002
rect 327356 176112 327408 176118
rect 327356 176054 327408 176060
rect 327264 169040 327316 169046
rect 327264 168982 327316 168988
rect 327368 159390 327396 176054
rect 327356 159384 327408 159390
rect 327356 159326 327408 159332
rect 327172 144832 327224 144838
rect 327172 144774 327224 144780
rect 328368 144220 328420 144226
rect 328368 144162 328420 144168
rect 328380 131170 328408 144162
rect 328368 131164 328420 131170
rect 328368 131106 328420 131112
rect 328380 131034 328408 131106
rect 328368 131028 328420 131034
rect 328368 130970 328420 130976
rect 327080 122528 327132 122534
rect 327080 122470 327132 122476
rect 327538 121408 327594 121417
rect 327538 121343 327540 121352
rect 327592 121343 327594 121352
rect 327540 121314 327592 121320
rect 327724 115116 327776 115122
rect 327724 115058 327776 115064
rect 327080 110764 327132 110770
rect 327080 110706 327132 110712
rect 325792 108384 325844 108390
rect 325792 108326 325844 108332
rect 325514 107128 325570 107137
rect 325514 107063 325570 107072
rect 324332 105318 324452 105346
rect 322938 104000 322994 104009
rect 322938 103935 322994 103944
rect 322952 103562 322980 103935
rect 322940 103556 322992 103562
rect 322940 103498 322992 103504
rect 324332 101538 324360 105318
rect 324412 103488 324464 103494
rect 324412 103430 324464 103436
rect 324424 102513 324452 103430
rect 325606 103184 325662 103193
rect 325662 103142 325740 103170
rect 325606 103119 325662 103128
rect 324410 102504 324466 102513
rect 324410 102439 324466 102448
rect 324332 101510 324728 101538
rect 324596 101448 324648 101454
rect 324596 101390 324648 101396
rect 324608 100881 324636 101390
rect 324594 100872 324650 100881
rect 324594 100807 324650 100816
rect 322938 100192 322994 100201
rect 322938 100127 322994 100136
rect 321744 96620 321796 96626
rect 321744 96562 321796 96568
rect 322952 94926 322980 100127
rect 324318 99376 324374 99385
rect 324318 99311 324320 99320
rect 324372 99311 324374 99320
rect 324320 99282 324372 99288
rect 324412 99272 324464 99278
rect 324412 99214 324464 99220
rect 324424 98569 324452 99214
rect 324410 98560 324466 98569
rect 324410 98495 324466 98504
rect 324608 98410 324636 100807
rect 324424 98382 324636 98410
rect 324320 96620 324372 96626
rect 324320 96562 324372 96568
rect 324332 96393 324360 96562
rect 324318 96384 324374 96393
rect 324318 96319 324374 96328
rect 322940 94920 322992 94926
rect 322940 94862 322992 94868
rect 322952 93906 322980 94862
rect 322940 93900 322992 93906
rect 322940 93842 322992 93848
rect 324318 93256 324374 93265
rect 324318 93191 324374 93200
rect 324332 93158 324360 93191
rect 324320 93152 324372 93158
rect 324320 93094 324372 93100
rect 324332 91050 324360 93094
rect 324320 91044 324372 91050
rect 324320 90986 324372 90992
rect 321572 84166 321692 84194
rect 321572 81394 321600 84166
rect 324424 82822 324452 98382
rect 324594 97880 324650 97889
rect 324594 97815 324650 97824
rect 324502 93800 324558 93809
rect 324608 93786 324636 97815
rect 324700 95198 324728 101510
rect 324688 95192 324740 95198
rect 324688 95134 324740 95140
rect 325712 95130 325740 103142
rect 325700 95124 325752 95130
rect 325700 95066 325752 95072
rect 325712 93906 325740 95066
rect 325700 93900 325752 93906
rect 325700 93842 325752 93848
rect 324558 93758 324636 93786
rect 324502 93735 324558 93744
rect 324504 87644 324556 87650
rect 324504 87586 324556 87592
rect 324412 82816 324464 82822
rect 324412 82758 324464 82764
rect 321560 81388 321612 81394
rect 321560 81330 321612 81336
rect 320180 79348 320232 79354
rect 320180 79290 320232 79296
rect 320192 16574 320220 79290
rect 323584 32564 323636 32570
rect 323584 32506 323636 32512
rect 311912 16546 312216 16574
rect 313292 16546 313872 16574
rect 316144 16546 316264 16574
rect 317432 16546 318104 16574
rect 320192 16546 320496 16574
rect 311440 15972 311492 15978
rect 311440 15914 311492 15920
rect 309876 3324 309928 3330
rect 309876 3266 309928 3272
rect 310244 2984 310296 2990
rect 310244 2926 310296 2932
rect 310256 480 310284 2926
rect 311452 480 311480 15914
rect 306718 354 306830 480
rect 306392 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 354 312216 16546
rect 313844 480 313872 16546
rect 315028 3324 315080 3330
rect 315028 3266 315080 3272
rect 315040 480 315068 3266
rect 316236 480 316264 16546
rect 317328 3392 317380 3398
rect 317328 3334 317380 3340
rect 317340 480 317368 3334
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 319720 3596 319772 3602
rect 319720 3538 319772 3544
rect 319732 480 319760 3538
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 322112 3460 322164 3466
rect 322112 3402 322164 3408
rect 323308 3460 323360 3466
rect 323308 3402 323360 3408
rect 322124 480 322152 3402
rect 323320 480 323348 3402
rect 323596 3398 323624 32506
rect 324516 6914 324544 87586
rect 324608 84194 324636 93758
rect 327092 89690 327120 110706
rect 327736 93854 327764 115058
rect 327736 93826 327948 93854
rect 327080 89684 327132 89690
rect 327080 89626 327132 89632
rect 327920 86970 327948 93826
rect 328368 89684 328420 89690
rect 328368 89626 328420 89632
rect 328380 88194 328408 89626
rect 328368 88188 328420 88194
rect 328368 88130 328420 88136
rect 327908 86964 327960 86970
rect 327908 86906 327960 86912
rect 327920 85513 327948 86906
rect 327906 85504 327962 85513
rect 327906 85439 327962 85448
rect 324608 84166 325004 84194
rect 324976 80034 325004 84166
rect 327080 83496 327132 83502
rect 327080 83438 327132 83444
rect 324964 80028 325016 80034
rect 324964 79970 325016 79976
rect 327092 16574 327120 83438
rect 328472 16574 328500 267038
rect 329104 191140 329156 191146
rect 329104 191082 329156 191088
rect 328552 177472 328604 177478
rect 328552 177414 328604 177420
rect 328564 137970 328592 177414
rect 328552 137964 328604 137970
rect 328552 137906 328604 137912
rect 327092 16546 328040 16574
rect 328472 16546 328776 16574
rect 324424 6886 324544 6914
rect 323584 3392 323636 3398
rect 323584 3334 323636 3340
rect 324424 480 324452 6886
rect 326804 3528 326856 3534
rect 326804 3470 326856 3476
rect 325608 3392 325660 3398
rect 325608 3334 325660 3340
rect 325620 480 325648 3334
rect 326816 480 326844 3470
rect 328012 480 328040 16546
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 328748 354 328776 16546
rect 329116 3534 329144 191082
rect 329208 187678 329236 360470
rect 330484 214600 330536 214606
rect 330484 214542 330536 214548
rect 329840 210452 329892 210458
rect 329840 210394 329892 210400
rect 329196 187672 329248 187678
rect 329196 187614 329248 187620
rect 329196 185632 329248 185638
rect 329196 185574 329248 185580
rect 329208 169726 329236 185574
rect 329196 169720 329248 169726
rect 329196 169662 329248 169668
rect 329196 149116 329248 149122
rect 329196 149058 329248 149064
rect 329208 124030 329236 149058
rect 329852 137902 329880 210394
rect 330496 193866 330524 214542
rect 330484 193860 330536 193866
rect 330484 193802 330536 193808
rect 330496 190454 330524 193802
rect 330496 190426 330616 190454
rect 330484 188624 330536 188630
rect 330484 188566 330536 188572
rect 330496 187610 330524 188566
rect 330484 187604 330536 187610
rect 330484 187546 330536 187552
rect 329932 175976 329984 175982
rect 329932 175918 329984 175924
rect 329840 137896 329892 137902
rect 329840 137838 329892 137844
rect 329196 124024 329248 124030
rect 329196 123966 329248 123972
rect 329944 110430 329972 175918
rect 330496 144906 330524 187546
rect 330588 164150 330616 190426
rect 330576 164144 330628 164150
rect 330576 164086 330628 164092
rect 330576 145648 330628 145654
rect 330576 145590 330628 145596
rect 330484 144900 330536 144906
rect 330484 144842 330536 144848
rect 330300 137896 330352 137902
rect 330300 137838 330352 137844
rect 330312 137290 330340 137838
rect 330300 137284 330352 137290
rect 330300 137226 330352 137232
rect 330588 118590 330616 145590
rect 330576 118584 330628 118590
rect 330576 118526 330628 118532
rect 329932 110424 329984 110430
rect 329932 110366 329984 110372
rect 329944 109721 329972 110366
rect 329930 109712 329986 109721
rect 329930 109647 329986 109656
rect 329196 108384 329248 108390
rect 329196 108326 329248 108332
rect 329208 85542 329236 108326
rect 329196 85536 329248 85542
rect 329196 85478 329248 85484
rect 331232 3602 331260 364482
rect 332600 360460 332652 360466
rect 332600 360402 332652 360408
rect 331864 264240 331916 264246
rect 331864 264182 331916 264188
rect 331312 213920 331364 213926
rect 331312 213862 331364 213868
rect 331324 150414 331352 213862
rect 331494 161256 331550 161265
rect 331494 161191 331550 161200
rect 331508 160750 331536 161191
rect 331496 160744 331548 160750
rect 331496 160686 331548 160692
rect 331312 150408 331364 150414
rect 331312 150350 331364 150356
rect 331312 75268 331364 75274
rect 331312 75210 331364 75216
rect 331220 3596 331272 3602
rect 331220 3538 331272 3544
rect 329104 3528 329156 3534
rect 329104 3470 329156 3476
rect 330392 3528 330444 3534
rect 330392 3470 330444 3476
rect 330404 480 330432 3470
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331324 354 331352 75210
rect 331876 3602 331904 264182
rect 331956 262268 332008 262274
rect 331956 262210 332008 262216
rect 331968 213926 331996 262210
rect 331956 213920 332008 213926
rect 331956 213862 332008 213868
rect 332048 189916 332100 189922
rect 332048 189858 332100 189864
rect 332060 169726 332088 189858
rect 332048 169720 332100 169726
rect 332048 169662 332100 169668
rect 331956 169040 332008 169046
rect 331956 168982 332008 168988
rect 331968 95062 331996 168982
rect 331956 95056 332008 95062
rect 331956 94998 332008 95004
rect 332612 6186 332640 360402
rect 337476 316736 337528 316742
rect 337476 316678 337528 316684
rect 337384 287156 337436 287162
rect 337384 287098 337436 287104
rect 333242 274816 333298 274825
rect 333242 274751 333298 274760
rect 333256 228954 333284 274751
rect 333980 242208 334032 242214
rect 333980 242150 334032 242156
rect 333244 228948 333296 228954
rect 333244 228890 333296 228896
rect 333256 228342 333284 228890
rect 332692 228336 332744 228342
rect 332692 228278 332744 228284
rect 333244 228336 333296 228342
rect 333244 228278 333296 228284
rect 332704 143546 332732 228278
rect 333244 199504 333296 199510
rect 333244 199446 333296 199452
rect 333256 190398 333284 199446
rect 333244 190392 333296 190398
rect 333244 190334 333296 190340
rect 332784 177608 332836 177614
rect 332784 177550 332836 177556
rect 332692 143540 332744 143546
rect 332692 143482 332744 143488
rect 332796 131102 332824 177550
rect 333256 164218 333284 190334
rect 333244 164212 333296 164218
rect 333244 164154 333296 164160
rect 333888 150476 333940 150482
rect 333888 150418 333940 150424
rect 332784 131096 332836 131102
rect 332784 131038 332836 131044
rect 332796 130422 332824 131038
rect 332784 130416 332836 130422
rect 332784 130358 332836 130364
rect 333900 81326 333928 150418
rect 333888 81320 333940 81326
rect 333888 81262 333940 81268
rect 333244 43580 333296 43586
rect 333244 43522 333296 43528
rect 332692 33924 332744 33930
rect 332692 33866 332744 33872
rect 332600 6180 332652 6186
rect 332600 6122 332652 6128
rect 331864 3596 331916 3602
rect 331864 3538 331916 3544
rect 332704 480 332732 33866
rect 333256 3534 333284 43522
rect 333992 16574 334020 242150
rect 335360 240780 335412 240786
rect 335360 240722 335412 240728
rect 334164 198280 334216 198286
rect 334164 198222 334216 198228
rect 334072 191888 334124 191894
rect 334072 191830 334124 191836
rect 334084 124098 334112 191830
rect 334176 150414 334204 198222
rect 334256 176180 334308 176186
rect 334256 176122 334308 176128
rect 334268 154494 334296 176122
rect 334256 154488 334308 154494
rect 334256 154430 334308 154436
rect 334624 154488 334676 154494
rect 334624 154430 334676 154436
rect 334636 153882 334664 154430
rect 334624 153876 334676 153882
rect 334624 153818 334676 153824
rect 334164 150408 334216 150414
rect 334164 150350 334216 150356
rect 334176 149122 334204 150350
rect 334164 149116 334216 149122
rect 334164 149058 334216 149064
rect 334072 124092 334124 124098
rect 334072 124034 334124 124040
rect 333992 16546 334664 16574
rect 333888 3596 333940 3602
rect 333888 3538 333940 3544
rect 333244 3528 333296 3534
rect 333244 3470 333296 3476
rect 333900 480 333928 3538
rect 331558 354 331670 480
rect 331324 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 16546
rect 335372 3482 335400 240722
rect 336740 214668 336792 214674
rect 336740 214610 336792 214616
rect 335544 209092 335596 209098
rect 335544 209034 335596 209040
rect 335452 199640 335504 199646
rect 335452 199582 335504 199588
rect 335464 6322 335492 199582
rect 335556 150482 335584 209034
rect 335636 181620 335688 181626
rect 335636 181562 335688 181568
rect 335544 150476 335596 150482
rect 335544 150418 335596 150424
rect 335648 147626 335676 181562
rect 335636 147620 335688 147626
rect 335636 147562 335688 147568
rect 336752 114442 336780 214610
rect 336832 207664 336884 207670
rect 336832 207606 336884 207612
rect 336844 145586 336872 207606
rect 337396 178838 337424 287098
rect 337488 242214 337516 316678
rect 340142 273864 340198 273873
rect 340142 273799 340198 273808
rect 337476 242208 337528 242214
rect 337476 242150 337528 242156
rect 338212 218748 338264 218754
rect 338212 218690 338264 218696
rect 338118 211848 338174 211857
rect 338118 211783 338174 211792
rect 337476 184340 337528 184346
rect 337476 184282 337528 184288
rect 337384 178832 337436 178838
rect 337384 178774 337436 178780
rect 337488 166326 337516 184282
rect 337476 166320 337528 166326
rect 337476 166262 337528 166268
rect 337384 164348 337436 164354
rect 337384 164290 337436 164296
rect 336832 145580 336884 145586
rect 336832 145522 336884 145528
rect 336740 114436 336792 114442
rect 336740 114378 336792 114384
rect 337396 105602 337424 164290
rect 337488 151774 337516 166262
rect 337476 151768 337528 151774
rect 337476 151710 337528 151716
rect 337476 145580 337528 145586
rect 337476 145522 337528 145528
rect 337488 133210 337516 145522
rect 337476 133204 337528 133210
rect 337476 133146 337528 133152
rect 337476 122120 337528 122126
rect 337476 122062 337528 122068
rect 337384 105596 337436 105602
rect 337384 105538 337436 105544
rect 337488 101454 337516 122062
rect 338028 114436 338080 114442
rect 338028 114378 338080 114384
rect 338040 113830 338068 114378
rect 338028 113824 338080 113830
rect 338028 113766 338080 113772
rect 338132 113150 338160 211783
rect 338224 150346 338252 218690
rect 340156 210662 340184 273799
rect 340144 210656 340196 210662
rect 340144 210598 340196 210604
rect 340144 204944 340196 204950
rect 340144 204886 340196 204892
rect 340156 202230 340184 204886
rect 340144 202224 340196 202230
rect 340144 202166 340196 202172
rect 338856 195288 338908 195294
rect 338856 195230 338908 195236
rect 338764 177540 338816 177546
rect 338764 177482 338816 177488
rect 338212 150340 338264 150346
rect 338212 150282 338264 150288
rect 338224 149734 338252 150282
rect 338212 149728 338264 149734
rect 338212 149670 338264 149676
rect 338120 113144 338172 113150
rect 338120 113086 338172 113092
rect 338132 112538 338160 113086
rect 338120 112532 338172 112538
rect 338120 112474 338172 112480
rect 337476 101448 337528 101454
rect 337476 101390 337528 101396
rect 338776 85474 338804 177482
rect 338868 143546 338896 195230
rect 339500 182912 339552 182918
rect 339500 182854 339552 182860
rect 339512 144226 339540 182854
rect 339500 144220 339552 144226
rect 339500 144162 339552 144168
rect 338856 143540 338908 143546
rect 338856 143482 338908 143488
rect 338868 136542 338896 143482
rect 338856 136536 338908 136542
rect 338856 136478 338908 136484
rect 340156 115258 340184 202166
rect 340236 199436 340288 199442
rect 340236 199378 340288 199384
rect 340248 120018 340276 199378
rect 340788 129056 340840 129062
rect 340786 129024 340788 129033
rect 340840 129024 340842 129033
rect 340786 128959 340842 128968
rect 340236 120012 340288 120018
rect 340236 119954 340288 119960
rect 340248 118658 340276 119954
rect 340236 118652 340288 118658
rect 340236 118594 340288 118600
rect 340144 115252 340196 115258
rect 340144 115194 340196 115200
rect 338764 85468 338816 85474
rect 338764 85410 338816 85416
rect 339498 51776 339554 51785
rect 339498 51711 339554 51720
rect 336738 42120 336794 42129
rect 336738 42055 336794 42064
rect 336752 16574 336780 42055
rect 336752 16546 337056 16574
rect 335452 6316 335504 6322
rect 335452 6258 335504 6264
rect 335372 3454 336320 3482
rect 336292 480 336320 3454
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337028 354 337056 16546
rect 338670 3496 338726 3505
rect 338670 3431 338726 3440
rect 338684 480 338712 3431
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339512 354 339540 51711
rect 340892 3466 340920 367270
rect 347044 356244 347096 356250
rect 347044 356186 347096 356192
rect 345664 291304 345716 291310
rect 345664 291246 345716 291252
rect 342904 287088 342956 287094
rect 342904 287030 342956 287036
rect 341524 283008 341576 283014
rect 341524 282950 341576 282956
rect 341536 233238 341564 282950
rect 341524 233232 341576 233238
rect 341524 233174 341576 233180
rect 342916 226166 342944 287030
rect 342996 244928 343048 244934
rect 342996 244870 343048 244876
rect 342904 226160 342956 226166
rect 342904 226102 342956 226108
rect 343008 222154 343036 244870
rect 345676 237250 345704 291246
rect 345756 273284 345808 273290
rect 345756 273226 345808 273232
rect 345664 237244 345716 237250
rect 345664 237186 345716 237192
rect 345768 227730 345796 273226
rect 345020 227724 345072 227730
rect 345020 227666 345072 227672
rect 345756 227724 345808 227730
rect 345756 227666 345808 227672
rect 342352 222148 342404 222154
rect 342352 222090 342404 222096
rect 342996 222148 343048 222154
rect 342996 222090 343048 222096
rect 340972 211812 341024 211818
rect 340972 211754 341024 211760
rect 340880 3460 340932 3466
rect 340880 3402 340932 3408
rect 340984 480 341012 211754
rect 342260 206440 342312 206446
rect 342260 206382 342312 206388
rect 341524 182232 341576 182238
rect 341524 182174 341576 182180
rect 341064 181688 341116 181694
rect 341064 181630 341116 181636
rect 341076 133890 341104 181630
rect 341064 133884 341116 133890
rect 341064 133826 341116 133832
rect 341248 133884 341300 133890
rect 341248 133826 341300 133832
rect 341260 133278 341288 133826
rect 341248 133272 341300 133278
rect 341248 133214 341300 133220
rect 341536 122806 341564 182174
rect 341524 122800 341576 122806
rect 341524 122742 341576 122748
rect 342272 16574 342300 206382
rect 342364 96626 342392 222090
rect 344284 211812 344336 211818
rect 344284 211754 344336 211760
rect 342442 207632 342498 207641
rect 342442 207567 342498 207576
rect 342456 155922 342484 207567
rect 343732 196716 343784 196722
rect 343732 196658 343784 196664
rect 342536 182980 342588 182986
rect 342536 182922 342588 182928
rect 342444 155916 342496 155922
rect 342444 155858 342496 155864
rect 342456 155242 342484 155858
rect 342444 155236 342496 155242
rect 342444 155178 342496 155184
rect 342548 151814 342576 182922
rect 343640 176044 343692 176050
rect 343640 175986 343692 175992
rect 342456 151786 342576 151814
rect 342456 146266 342484 151786
rect 342444 146260 342496 146266
rect 342444 146202 342496 146208
rect 342456 145654 342484 146202
rect 342444 145648 342496 145654
rect 342444 145590 342496 145596
rect 342352 96620 342404 96626
rect 342352 96562 342404 96568
rect 342272 16546 342944 16574
rect 342168 3460 342220 3466
rect 342168 3402 342220 3408
rect 342180 480 342208 3402
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 16546
rect 343652 3466 343680 175986
rect 343744 121446 343772 196658
rect 343824 192500 343876 192506
rect 343824 192442 343876 192448
rect 343836 136610 343864 192442
rect 344296 167006 344324 211754
rect 344284 167000 344336 167006
rect 344284 166942 344336 166948
rect 343824 136604 343876 136610
rect 343824 136546 343876 136552
rect 344468 136604 344520 136610
rect 344468 136546 344520 136552
rect 344480 135930 344508 136546
rect 344468 135924 344520 135930
rect 344468 135866 344520 135872
rect 343732 121440 343784 121446
rect 343732 121382 343784 121388
rect 343744 120766 343772 121382
rect 343732 120760 343784 120766
rect 343732 120702 343784 120708
rect 345032 99278 345060 227666
rect 346400 213240 346452 213246
rect 346400 213182 346452 213188
rect 345296 198008 345348 198014
rect 345296 197950 345348 197956
rect 345204 192568 345256 192574
rect 345204 192510 345256 192516
rect 345112 180260 345164 180266
rect 345112 180202 345164 180208
rect 345124 115938 345152 180202
rect 345216 142118 345244 192510
rect 345308 157282 345336 197950
rect 345296 157276 345348 157282
rect 345296 157218 345348 157224
rect 346308 157276 346360 157282
rect 346308 157218 346360 157224
rect 346320 156670 346348 157218
rect 346308 156664 346360 156670
rect 346308 156606 346360 156612
rect 345204 142112 345256 142118
rect 345204 142054 345256 142060
rect 345112 115932 345164 115938
rect 345112 115874 345164 115880
rect 346308 115932 346360 115938
rect 346308 115874 346360 115880
rect 346320 115161 346348 115874
rect 346306 115152 346362 115161
rect 346306 115087 346362 115096
rect 346412 103494 346440 213182
rect 346492 180328 346544 180334
rect 346492 180270 346544 180276
rect 346504 154562 346532 180270
rect 346492 154556 346544 154562
rect 346492 154498 346544 154504
rect 346400 103488 346452 103494
rect 346400 103430 346452 103436
rect 345020 99272 345072 99278
rect 345020 99214 345072 99220
rect 347056 77178 347084 356186
rect 351184 346452 351236 346458
rect 351184 346394 351236 346400
rect 349804 342916 349856 342922
rect 349804 342858 349856 342864
rect 347686 285696 347742 285705
rect 347686 285631 347742 285640
rect 347700 227633 347728 285631
rect 347686 227624 347742 227633
rect 347686 227559 347742 227568
rect 347700 226386 347728 227559
rect 347700 226358 347820 226386
rect 347792 224874 347820 226358
rect 347136 224868 347188 224874
rect 347136 224810 347188 224816
rect 347780 224868 347832 224874
rect 347780 224810 347832 224816
rect 347148 132394 347176 224810
rect 349160 214736 349212 214742
rect 349160 214678 349212 214684
rect 347688 213240 347740 213246
rect 347688 213182 347740 213188
rect 347700 212566 347728 213182
rect 347688 212560 347740 212566
rect 347688 212502 347740 212508
rect 347872 203652 347924 203658
rect 347872 203594 347924 203600
rect 347780 198212 347832 198218
rect 347780 198154 347832 198160
rect 347688 154556 347740 154562
rect 347688 154498 347740 154504
rect 347700 153950 347728 154498
rect 347688 153944 347740 153950
rect 347688 153886 347740 153892
rect 347136 132388 347188 132394
rect 347136 132330 347188 132336
rect 347792 111790 347820 198154
rect 347884 125526 347912 203594
rect 347964 202156 348016 202162
rect 347964 202098 348016 202104
rect 347976 135250 348004 202098
rect 347964 135244 348016 135250
rect 347964 135186 348016 135192
rect 347872 125520 347924 125526
rect 347872 125462 347924 125468
rect 347780 111784 347832 111790
rect 347780 111726 347832 111732
rect 347792 111110 347820 111726
rect 347780 111104 347832 111110
rect 347780 111046 347832 111052
rect 347044 77172 347096 77178
rect 347044 77114 347096 77120
rect 345018 24168 345074 24177
rect 345018 24103 345074 24112
rect 345032 16574 345060 24103
rect 345032 16546 345336 16574
rect 344560 3528 344612 3534
rect 344560 3470 344612 3476
rect 343640 3460 343692 3466
rect 343640 3402 343692 3408
rect 344572 480 344600 3470
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345308 354 345336 16546
rect 348056 6248 348108 6254
rect 348056 6190 348108 6196
rect 346952 2984 347004 2990
rect 346952 2926 347004 2932
rect 346964 480 346992 2926
rect 348068 480 348096 6190
rect 349172 3534 349200 214678
rect 349250 200696 349306 200705
rect 349250 200631 349306 200640
rect 349264 125594 349292 200631
rect 349344 192908 349396 192914
rect 349344 192850 349396 192856
rect 349252 125588 349304 125594
rect 349252 125530 349304 125536
rect 349356 120086 349384 192850
rect 349816 153202 349844 342858
rect 350540 271176 350592 271182
rect 350540 271118 350592 271124
rect 349804 153196 349856 153202
rect 349804 153138 349856 153144
rect 349620 125588 349672 125594
rect 349620 125530 349672 125536
rect 349632 124914 349660 125530
rect 349620 124908 349672 124914
rect 349620 124850 349672 124856
rect 349344 120080 349396 120086
rect 349344 120022 349396 120028
rect 349356 119406 349384 120022
rect 349344 119400 349396 119406
rect 349344 119342 349396 119348
rect 350552 16574 350580 271118
rect 350632 182844 350684 182850
rect 350632 182786 350684 182792
rect 350644 124166 350672 182786
rect 350632 124160 350684 124166
rect 350632 124102 350684 124108
rect 350644 123486 350672 124102
rect 350632 123480 350684 123486
rect 350632 123422 350684 123428
rect 351196 92206 351224 346394
rect 352564 278112 352616 278118
rect 352564 278054 352616 278060
rect 352576 228886 352604 278054
rect 354600 276078 354628 700334
rect 374644 359032 374696 359038
rect 374644 358974 374696 358980
rect 363604 357604 363656 357610
rect 363604 357546 363656 357552
rect 355322 357504 355378 357513
rect 355322 357439 355378 357448
rect 353944 276072 353996 276078
rect 353944 276014 353996 276020
rect 354588 276072 354640 276078
rect 354588 276014 354640 276020
rect 353300 246424 353352 246430
rect 353300 246366 353352 246372
rect 353312 244254 353340 246366
rect 353300 244248 353352 244254
rect 353300 244190 353352 244196
rect 353956 230314 353984 276014
rect 354680 237380 354732 237386
rect 354680 237322 354732 237328
rect 353944 230308 353996 230314
rect 353944 230250 353996 230256
rect 352564 228880 352616 228886
rect 352564 228822 352616 228828
rect 353944 227180 353996 227186
rect 353944 227122 353996 227128
rect 353298 222864 353354 222873
rect 353298 222799 353354 222808
rect 352564 210520 352616 210526
rect 352564 210462 352616 210468
rect 351276 205692 351328 205698
rect 351276 205634 351328 205640
rect 351288 108322 351316 205634
rect 351920 193996 351972 194002
rect 351920 193938 351972 193944
rect 351276 108316 351328 108322
rect 351276 108258 351328 108264
rect 351184 92200 351236 92206
rect 351184 92142 351236 92148
rect 350552 16546 351224 16574
rect 349252 13252 349304 13258
rect 349252 13194 349304 13200
rect 349160 3528 349212 3534
rect 349160 3470 349212 3476
rect 349264 480 349292 13194
rect 350448 3528 350500 3534
rect 350448 3470 350500 3476
rect 350460 480 350488 3470
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 351932 2990 351960 193938
rect 352576 114578 352604 210462
rect 353312 135182 353340 222799
rect 353300 135176 353352 135182
rect 353300 135118 353352 135124
rect 352564 114572 352616 114578
rect 352564 114514 352616 114520
rect 353956 109002 353984 227122
rect 354036 192636 354088 192642
rect 354036 192578 354088 192584
rect 354048 173874 354076 192578
rect 354036 173868 354088 173874
rect 354036 173810 354088 173816
rect 354036 171148 354088 171154
rect 354036 171090 354088 171096
rect 353944 108996 353996 109002
rect 353944 108938 353996 108944
rect 354048 89486 354076 171090
rect 354692 117978 354720 237322
rect 354770 184376 354826 184385
rect 354770 184311 354826 184320
rect 354784 128314 354812 184311
rect 354772 128308 354824 128314
rect 354772 128250 354824 128256
rect 354680 117972 354732 117978
rect 354680 117914 354732 117920
rect 354680 114572 354732 114578
rect 354680 114514 354732 114520
rect 354692 106282 354720 114514
rect 354680 106276 354732 106282
rect 354680 106218 354732 106224
rect 355336 95266 355364 357439
rect 359464 349852 359516 349858
rect 359464 349794 359516 349800
rect 356796 288448 356848 288454
rect 356796 288390 356848 288396
rect 356704 281580 356756 281586
rect 356704 281522 356756 281528
rect 355416 255332 355468 255338
rect 355416 255274 355468 255280
rect 355428 237386 355456 255274
rect 355416 237380 355468 237386
rect 355416 237322 355468 237328
rect 356060 220108 356112 220114
rect 356060 220050 356112 220056
rect 355968 128308 356020 128314
rect 355968 128250 356020 128256
rect 355980 127634 356008 128250
rect 355968 127628 356020 127634
rect 355968 127570 356020 127576
rect 356072 117298 356100 220050
rect 356716 129062 356744 281522
rect 356808 228857 356836 288390
rect 358082 272504 358138 272513
rect 358082 272439 358138 272448
rect 358096 246362 358124 272439
rect 358084 246356 358136 246362
rect 358084 246298 358136 246304
rect 356794 228848 356850 228857
rect 356794 228783 356850 228792
rect 357992 217320 358044 217326
rect 357992 217262 358044 217268
rect 358004 216578 358032 217262
rect 357992 216572 358044 216578
rect 357992 216514 358044 216520
rect 358176 216572 358228 216578
rect 358176 216514 358228 216520
rect 358084 191276 358136 191282
rect 358084 191218 358136 191224
rect 356888 181484 356940 181490
rect 356888 181426 356940 181432
rect 356900 170338 356928 181426
rect 356888 170332 356940 170338
rect 356888 170274 356940 170280
rect 356796 169788 356848 169794
rect 356796 169730 356848 169736
rect 356704 129056 356756 129062
rect 356704 128998 356756 129004
rect 356060 117292 356112 117298
rect 356060 117234 356112 117240
rect 355324 95260 355376 95266
rect 355324 95202 355376 95208
rect 356808 93634 356836 169730
rect 357348 117292 357400 117298
rect 357348 117234 357400 117240
rect 357360 116521 357388 117234
rect 357346 116512 357402 116521
rect 357346 116447 357402 116456
rect 356796 93628 356848 93634
rect 356796 93570 356848 93576
rect 354036 89480 354088 89486
rect 354036 89422 354088 89428
rect 358096 82822 358124 191218
rect 358188 140758 358216 216514
rect 358820 191208 358872 191214
rect 358820 191150 358872 191156
rect 358176 140752 358228 140758
rect 358176 140694 358228 140700
rect 358832 132462 358860 191150
rect 358820 132456 358872 132462
rect 358820 132398 358872 132404
rect 359476 89418 359504 349794
rect 360844 338156 360896 338162
rect 360844 338098 360896 338104
rect 359648 283212 359700 283218
rect 359648 283154 359700 283160
rect 359554 280256 359610 280265
rect 359554 280191 359610 280200
rect 359568 234569 359596 280191
rect 359660 240038 359688 283154
rect 360856 260846 360884 338098
rect 362224 290012 362276 290018
rect 362224 289954 362276 289960
rect 360934 281616 360990 281625
rect 360934 281551 360990 281560
rect 360844 260840 360896 260846
rect 360844 260782 360896 260788
rect 360844 256760 360896 256766
rect 360844 256702 360896 256708
rect 359648 240032 359700 240038
rect 359648 239974 359700 239980
rect 359554 234560 359610 234569
rect 359554 234495 359610 234504
rect 360292 225480 360344 225486
rect 360292 225422 360344 225428
rect 360200 224936 360252 224942
rect 360200 224878 360252 224884
rect 360212 224534 360240 224878
rect 360200 224528 360252 224534
rect 360200 224470 360252 224476
rect 359554 178800 359610 178809
rect 359554 178735 359610 178744
rect 359568 142050 359596 178735
rect 359648 170332 359700 170338
rect 359648 170274 359700 170280
rect 359660 158778 359688 170274
rect 359648 158772 359700 158778
rect 359648 158714 359700 158720
rect 359660 158642 359688 158714
rect 360212 158710 360240 224470
rect 360304 175234 360332 225422
rect 360856 224534 360884 256702
rect 360844 224528 360896 224534
rect 360844 224470 360896 224476
rect 360948 219366 360976 281551
rect 361028 233912 361080 233918
rect 361028 233854 361080 233860
rect 361040 226302 361068 233854
rect 361028 226296 361080 226302
rect 361028 226238 361080 226244
rect 361040 225486 361068 226238
rect 361028 225480 361080 225486
rect 361028 225422 361080 225428
rect 360936 219360 360988 219366
rect 360936 219302 360988 219308
rect 360844 203720 360896 203726
rect 360844 203662 360896 203668
rect 360292 175228 360344 175234
rect 360292 175170 360344 175176
rect 360200 158704 360252 158710
rect 360200 158646 360252 158652
rect 359648 158636 359700 158642
rect 359648 158578 359700 158584
rect 360108 142180 360160 142186
rect 360108 142122 360160 142128
rect 360120 142050 360148 142122
rect 359556 142044 359608 142050
rect 359556 141986 359608 141992
rect 360108 142044 360160 142050
rect 360108 141986 360160 141992
rect 359556 133272 359608 133278
rect 359556 133214 359608 133220
rect 359464 89412 359516 89418
rect 359464 89354 359516 89360
rect 359568 84182 359596 133214
rect 360856 92274 360884 203662
rect 360936 153944 360988 153950
rect 360936 153886 360988 153892
rect 360844 92268 360896 92274
rect 360844 92210 360896 92216
rect 360948 85338 360976 153886
rect 362236 96393 362264 289954
rect 362316 281580 362368 281586
rect 362316 281522 362368 281528
rect 362328 240106 362356 281522
rect 363616 276010 363644 357546
rect 367744 331900 367796 331906
rect 367744 331842 367796 331848
rect 363788 285864 363840 285870
rect 363788 285806 363840 285812
rect 363694 284880 363750 284889
rect 363694 284815 363750 284824
rect 363604 276004 363656 276010
rect 363604 275946 363656 275952
rect 363604 240168 363656 240174
rect 363604 240110 363656 240116
rect 362316 240100 362368 240106
rect 362316 240042 362368 240048
rect 363616 120018 363644 240110
rect 363708 231606 363736 284815
rect 363800 256766 363828 285806
rect 366364 284572 366416 284578
rect 366364 284514 366416 284520
rect 365076 284504 365128 284510
rect 365076 284446 365128 284452
rect 364984 277704 365036 277710
rect 364984 277646 365036 277652
rect 364248 276004 364300 276010
rect 364248 275946 364300 275952
rect 363788 256760 363840 256766
rect 363788 256702 363840 256708
rect 364260 243574 364288 275946
rect 363788 243568 363840 243574
rect 363788 243510 363840 243516
rect 364248 243568 364300 243574
rect 364248 243510 364300 243516
rect 363696 231600 363748 231606
rect 363696 231542 363748 231548
rect 363800 219434 363828 243510
rect 363788 219428 363840 219434
rect 363788 219370 363840 219376
rect 363696 178696 363748 178702
rect 363696 178638 363748 178644
rect 363604 120012 363656 120018
rect 363604 119954 363656 119960
rect 362222 96384 362278 96393
rect 362222 96319 362278 96328
rect 363708 89622 363736 178638
rect 364996 135182 365024 277646
rect 365088 238542 365116 284446
rect 365166 279032 365222 279041
rect 365166 278967 365222 278976
rect 365076 238536 365128 238542
rect 365076 238478 365128 238484
rect 365180 237318 365208 278967
rect 365168 237312 365220 237318
rect 365168 237254 365220 237260
rect 365076 177404 365128 177410
rect 365076 177346 365128 177352
rect 364984 135176 365036 135182
rect 364984 135118 365036 135124
rect 363696 89616 363748 89622
rect 363696 89558 363748 89564
rect 360936 85332 360988 85338
rect 360936 85274 360988 85280
rect 359556 84176 359608 84182
rect 359556 84118 359608 84124
rect 358084 82816 358136 82822
rect 358084 82758 358136 82764
rect 365088 79966 365116 177346
rect 366376 134570 366404 284514
rect 366456 269816 366508 269822
rect 366456 269758 366508 269764
rect 366468 235754 366496 269758
rect 366456 235748 366508 235754
rect 366456 235690 366508 235696
rect 366364 134564 366416 134570
rect 366364 134506 366416 134512
rect 367756 82754 367784 331842
rect 369124 329860 369176 329866
rect 369124 329802 369176 329808
rect 367928 280492 367980 280498
rect 367928 280434 367980 280440
rect 367836 276208 367888 276214
rect 367836 276150 367888 276156
rect 367848 125526 367876 276150
rect 367940 231810 367968 280434
rect 368478 241496 368534 241505
rect 368478 241431 368534 241440
rect 368492 241233 368520 241431
rect 368478 241224 368534 241233
rect 368478 241159 368534 241168
rect 367928 231804 367980 231810
rect 367928 231746 367980 231752
rect 367928 159384 367980 159390
rect 367928 159326 367980 159332
rect 367836 125520 367888 125526
rect 367836 125462 367888 125468
rect 367940 95470 367968 159326
rect 368492 99346 368520 241159
rect 369136 135998 369164 329802
rect 369308 288584 369360 288590
rect 369308 288526 369360 288532
rect 369216 281784 369268 281790
rect 369216 281726 369268 281732
rect 369228 234530 369256 281726
rect 369320 241505 369348 288526
rect 370596 285796 370648 285802
rect 370596 285738 370648 285744
rect 370504 275324 370556 275330
rect 370504 275266 370556 275272
rect 369306 241496 369362 241505
rect 369306 241431 369362 241440
rect 369216 234524 369268 234530
rect 369216 234466 369268 234472
rect 370516 187610 370544 275266
rect 370608 237153 370636 285738
rect 371884 284436 371936 284442
rect 371884 284378 371936 284384
rect 370594 237144 370650 237153
rect 370594 237079 370650 237088
rect 371896 230450 371924 284378
rect 371976 283144 372028 283150
rect 371976 283086 372028 283092
rect 371988 238649 372016 283086
rect 373356 283076 373408 283082
rect 373356 283018 373408 283024
rect 373264 278928 373316 278934
rect 373264 278870 373316 278876
rect 371974 238640 372030 238649
rect 371974 238575 372030 238584
rect 371884 230444 371936 230450
rect 371884 230386 371936 230392
rect 373276 216578 373304 278870
rect 373368 235890 373396 283018
rect 373356 235884 373408 235890
rect 373356 235826 373408 235832
rect 373998 224904 374054 224913
rect 373998 224839 374054 224848
rect 373264 216572 373316 216578
rect 373264 216514 373316 216520
rect 373354 200832 373410 200841
rect 373354 200767 373410 200776
rect 370596 195356 370648 195362
rect 370596 195298 370648 195304
rect 370504 187604 370556 187610
rect 370504 187546 370556 187552
rect 369216 162172 369268 162178
rect 369216 162114 369268 162120
rect 369124 135992 369176 135998
rect 369124 135934 369176 135940
rect 368480 99340 368532 99346
rect 368480 99282 368532 99288
rect 367928 95464 367980 95470
rect 367928 95406 367980 95412
rect 369228 88262 369256 162114
rect 370608 120086 370636 195298
rect 373264 144968 373316 144974
rect 373264 144910 373316 144916
rect 373276 137970 373304 144910
rect 373264 137964 373316 137970
rect 373264 137906 373316 137912
rect 373264 131776 373316 131782
rect 373264 131718 373316 131724
rect 370596 120080 370648 120086
rect 370596 120022 370648 120028
rect 369216 88256 369268 88262
rect 369216 88198 369268 88204
rect 367744 82748 367796 82754
rect 367744 82690 367796 82696
rect 365076 79960 365128 79966
rect 365076 79902 365128 79908
rect 373276 59362 373304 131718
rect 373368 129742 373396 200767
rect 373448 140072 373500 140078
rect 373448 140014 373500 140020
rect 373460 132462 373488 140014
rect 373448 132456 373500 132462
rect 373448 132398 373500 132404
rect 373356 129736 373408 129742
rect 373356 129678 373408 129684
rect 373446 129024 373502 129033
rect 373446 128959 373502 128968
rect 373460 81258 373488 128959
rect 374012 114510 374040 224839
rect 374000 114504 374052 114510
rect 374000 114446 374052 114452
rect 374656 92449 374684 358974
rect 377402 341456 377458 341465
rect 377402 341391 377458 341400
rect 374828 281920 374880 281926
rect 374828 281862 374880 281868
rect 374736 281852 374788 281858
rect 374736 281794 374788 281800
rect 374748 224913 374776 281794
rect 374840 238746 374868 281862
rect 376024 280424 376076 280430
rect 376024 280366 376076 280372
rect 374828 238740 374880 238746
rect 374828 238682 374880 238688
rect 374734 224904 374790 224913
rect 374734 224839 374790 224848
rect 376036 168298 376064 280366
rect 376024 168292 376076 168298
rect 376024 168234 376076 168240
rect 376024 153264 376076 153270
rect 376024 153206 376076 153212
rect 374736 127628 374788 127634
rect 374736 127570 374788 127576
rect 374642 92440 374698 92449
rect 374642 92375 374698 92384
rect 374748 84114 374776 127570
rect 376036 93430 376064 153206
rect 377416 122806 377444 341391
rect 381544 285728 381596 285734
rect 381544 285670 381596 285676
rect 377496 281716 377548 281722
rect 377496 281658 377548 281664
rect 377508 238610 377536 281658
rect 377680 280560 377732 280566
rect 377680 280502 377732 280508
rect 377586 280392 377642 280401
rect 377586 280327 377642 280336
rect 377600 238678 377628 280327
rect 377692 241466 377720 280502
rect 378876 279132 378928 279138
rect 378876 279074 378928 279080
rect 378784 247716 378836 247722
rect 378784 247658 378836 247664
rect 377680 241460 377732 241466
rect 377680 241402 377732 241408
rect 377588 238672 377640 238678
rect 377588 238614 377640 238620
rect 377496 238604 377548 238610
rect 377496 238546 377548 238552
rect 378140 225208 378192 225214
rect 378140 225150 378192 225156
rect 377496 156664 377548 156670
rect 377496 156606 377548 156612
rect 377404 122800 377456 122806
rect 377404 122742 377456 122748
rect 376116 112532 376168 112538
rect 376116 112474 376168 112480
rect 376128 95169 376156 112474
rect 376114 95160 376170 95169
rect 376114 95095 376170 95104
rect 376024 93424 376076 93430
rect 376024 93366 376076 93372
rect 374736 84108 374788 84114
rect 374736 84050 374788 84056
rect 377508 82686 377536 156606
rect 378152 126954 378180 225150
rect 378140 126948 378192 126954
rect 378140 126890 378192 126896
rect 378796 90914 378824 247658
rect 378888 226234 378916 279074
rect 380346 278896 380402 278905
rect 380346 278831 380402 278840
rect 379428 278792 379480 278798
rect 379428 278734 379480 278740
rect 379440 247042 379468 278734
rect 380164 277568 380216 277574
rect 380164 277510 380216 277516
rect 379428 247036 379480 247042
rect 379428 246978 379480 246984
rect 379440 246430 379468 246978
rect 379428 246424 379480 246430
rect 379428 246366 379480 246372
rect 378876 226228 378928 226234
rect 378876 226170 378928 226176
rect 378888 225214 378916 226170
rect 378876 225208 378928 225214
rect 378876 225150 378928 225156
rect 380176 147626 380204 277510
rect 380254 274952 380310 274961
rect 380254 274887 380310 274896
rect 380268 190466 380296 274887
rect 380360 237289 380388 278831
rect 381556 276690 381584 285670
rect 381636 279064 381688 279070
rect 381636 279006 381688 279012
rect 381544 276684 381596 276690
rect 381544 276626 381596 276632
rect 381544 271924 381596 271930
rect 381544 271866 381596 271872
rect 380346 237280 380402 237289
rect 380346 237215 380402 237224
rect 380900 234864 380952 234870
rect 380900 234806 380952 234812
rect 380348 229764 380400 229770
rect 380348 229706 380400 229712
rect 380256 190460 380308 190466
rect 380256 190402 380308 190408
rect 380360 176662 380388 229706
rect 380440 180192 380492 180198
rect 380440 180134 380492 180140
rect 380348 176656 380400 176662
rect 380348 176598 380400 176604
rect 380256 164280 380308 164286
rect 380256 164222 380308 164228
rect 380164 147620 380216 147626
rect 380164 147562 380216 147568
rect 380164 142180 380216 142186
rect 380164 142122 380216 142128
rect 378876 131164 378928 131170
rect 378876 131106 378928 131112
rect 378888 96626 378916 131106
rect 378968 119400 379020 119406
rect 378968 119342 379020 119348
rect 378876 96620 378928 96626
rect 378876 96562 378928 96568
rect 378784 90908 378836 90914
rect 378784 90850 378836 90856
rect 378980 89690 379008 119342
rect 380176 95033 380204 142122
rect 380268 95334 380296 164222
rect 380452 162858 380480 180134
rect 380912 168366 380940 234806
rect 380900 168360 380952 168366
rect 380900 168302 380952 168308
rect 380440 162852 380492 162858
rect 380440 162794 380492 162800
rect 380348 158772 380400 158778
rect 380348 158714 380400 158720
rect 380256 95328 380308 95334
rect 380256 95270 380308 95276
rect 380162 95024 380218 95033
rect 380162 94959 380218 94968
rect 380360 92478 380388 158714
rect 380348 92472 380400 92478
rect 380348 92414 380400 92420
rect 381556 92138 381584 271866
rect 381648 235958 381676 279006
rect 382188 276684 382240 276690
rect 382188 276626 382240 276632
rect 381636 235952 381688 235958
rect 381636 235894 381688 235900
rect 381648 234870 381676 235894
rect 381636 234864 381688 234870
rect 381636 234806 381688 234812
rect 382200 197334 382228 276626
rect 382924 276276 382976 276282
rect 382924 276218 382976 276224
rect 382278 234696 382334 234705
rect 382278 234631 382334 234640
rect 382188 197328 382240 197334
rect 382188 197270 382240 197276
rect 381636 181552 381688 181558
rect 381636 181494 381688 181500
rect 381648 99346 381676 181494
rect 382292 171086 382320 234631
rect 382936 173913 382964 276218
rect 383016 276140 383068 276146
rect 383016 276082 383068 276088
rect 383028 189038 383056 276082
rect 383106 274680 383162 274689
rect 383106 274615 383162 274624
rect 383120 235929 383148 274615
rect 383106 235920 383162 235929
rect 383106 235855 383162 235864
rect 383120 234705 383148 235855
rect 383106 234696 383162 234705
rect 383106 234631 383162 234640
rect 383016 189032 383068 189038
rect 383016 188974 383068 188980
rect 383014 179480 383070 179489
rect 383014 179415 383070 179424
rect 382922 173904 382978 173913
rect 382922 173839 382978 173848
rect 382280 171080 382332 171086
rect 382280 171022 382332 171028
rect 382924 147688 382976 147694
rect 382924 147630 382976 147636
rect 381728 130416 381780 130422
rect 381728 130358 381780 130364
rect 381636 99340 381688 99346
rect 381636 99282 381688 99288
rect 381544 92132 381596 92138
rect 381544 92074 381596 92080
rect 378968 89684 379020 89690
rect 378968 89626 379020 89632
rect 381740 86834 381768 130358
rect 382936 94994 382964 147630
rect 383028 96558 383056 179415
rect 383108 120760 383160 120766
rect 383108 120702 383160 120708
rect 383016 96552 383068 96558
rect 383016 96494 383068 96500
rect 382924 94988 382976 94994
rect 382924 94930 382976 94936
rect 383120 88126 383148 120702
rect 383580 91089 383608 700334
rect 397472 698970 397500 703520
rect 397460 698964 397512 698970
rect 397460 698906 397512 698912
rect 391204 576904 391256 576910
rect 391204 576846 391256 576852
rect 388444 404388 388496 404394
rect 388444 404330 388496 404336
rect 387708 358080 387760 358086
rect 387708 358022 387760 358028
rect 385868 288516 385920 288522
rect 385868 288458 385920 288464
rect 384212 281648 384264 281654
rect 384212 281590 384264 281596
rect 384224 278118 384252 281590
rect 385038 279168 385094 279177
rect 385038 279103 385094 279112
rect 384212 278112 384264 278118
rect 384212 278054 384264 278060
rect 384302 277672 384358 277681
rect 384302 277607 384358 277616
rect 384316 142118 384344 277607
rect 384486 277536 384542 277545
rect 384486 277471 384542 277480
rect 384500 161401 384528 277471
rect 385052 274650 385080 279103
rect 385880 278050 385908 288458
rect 387616 284640 387668 284646
rect 387616 284582 387668 284588
rect 385868 278044 385920 278050
rect 385868 277986 385920 277992
rect 385684 277636 385736 277642
rect 385684 277578 385736 277584
rect 385040 274644 385092 274650
rect 385040 274586 385092 274592
rect 385132 223576 385184 223582
rect 385132 223518 385184 223524
rect 385040 220720 385092 220726
rect 385040 220662 385092 220668
rect 384486 161392 384542 161401
rect 384486 161327 384542 161336
rect 385052 157350 385080 220662
rect 385144 172514 385172 223518
rect 385132 172508 385184 172514
rect 385132 172450 385184 172456
rect 385040 157344 385092 157350
rect 385040 157286 385092 157292
rect 384396 155236 384448 155242
rect 384396 155178 384448 155184
rect 384304 142112 384356 142118
rect 384304 142054 384356 142060
rect 384304 138032 384356 138038
rect 384304 137974 384356 137980
rect 384316 93702 384344 137974
rect 384304 93696 384356 93702
rect 384304 93638 384356 93644
rect 383566 91080 383622 91089
rect 383566 91015 383622 91024
rect 383108 88120 383160 88126
rect 383108 88062 383160 88068
rect 384408 86902 384436 155178
rect 385696 143546 385724 277578
rect 385776 277500 385828 277506
rect 385776 277442 385828 277448
rect 385788 220726 385816 277442
rect 385868 276344 385920 276350
rect 385868 276286 385920 276292
rect 385880 223582 385908 276286
rect 386878 273456 386934 273465
rect 386878 273391 386934 273400
rect 386892 273290 386920 273391
rect 386880 273284 386932 273290
rect 386880 273226 386932 273232
rect 387154 270056 387210 270065
rect 387154 269991 387210 270000
rect 387168 269822 387196 269991
rect 387156 269816 387208 269822
rect 387156 269758 387208 269764
rect 387062 266656 387118 266665
rect 387062 266591 387118 266600
rect 386878 263256 386934 263265
rect 386878 263191 386934 263200
rect 386892 262274 386920 263191
rect 386880 262268 386932 262274
rect 386880 262210 386932 262216
rect 386880 260840 386932 260846
rect 386880 260782 386932 260788
rect 386892 260001 386920 260782
rect 386878 259992 386934 260001
rect 386878 259927 386934 259936
rect 386878 256456 386934 256465
rect 386878 256391 386934 256400
rect 386892 255338 386920 256391
rect 386880 255332 386932 255338
rect 386880 255274 386932 255280
rect 386878 253056 386934 253065
rect 386878 252991 386934 253000
rect 386892 252618 386920 252991
rect 386880 252612 386932 252618
rect 386880 252554 386932 252560
rect 386880 247036 386932 247042
rect 386880 246978 386932 246984
rect 386892 246401 386920 246978
rect 386878 246392 386934 246401
rect 386878 246327 386934 246336
rect 386604 243568 386656 243574
rect 386602 243536 386604 243545
rect 386656 243536 386658 243545
rect 386602 243471 386658 243480
rect 386878 240272 386934 240281
rect 386878 240207 386934 240216
rect 386892 240174 386920 240207
rect 386880 240168 386932 240174
rect 386880 240110 386932 240116
rect 387076 238814 387104 266591
rect 387522 249656 387578 249665
rect 387522 249591 387578 249600
rect 387536 244934 387564 249591
rect 387524 244928 387576 244934
rect 387524 244870 387576 244876
rect 387156 242208 387208 242214
rect 387156 242150 387208 242156
rect 387064 238808 387116 238814
rect 387064 238750 387116 238756
rect 386786 236736 386842 236745
rect 386786 236671 386842 236680
rect 386512 233980 386564 233986
rect 386512 233922 386564 233928
rect 386524 233481 386552 233922
rect 386800 233918 386828 236671
rect 386788 233912 386840 233918
rect 386788 233854 386840 233860
rect 386510 233472 386566 233481
rect 386510 233407 386566 233416
rect 386420 229764 386472 229770
rect 386420 229706 386472 229712
rect 386432 226681 386460 229706
rect 386972 227044 387024 227050
rect 386972 226986 387024 226992
rect 386418 226672 386474 226681
rect 386418 226607 386474 226616
rect 385868 223576 385920 223582
rect 385868 223518 385920 223524
rect 386984 223281 387012 226986
rect 386970 223272 387026 223281
rect 386970 223207 387026 223216
rect 387076 222193 387104 238750
rect 387168 230081 387196 242150
rect 387154 230072 387210 230081
rect 387154 230007 387210 230016
rect 387168 228750 387196 230007
rect 387156 228744 387208 228750
rect 387156 228686 387208 228692
rect 387154 223272 387210 223281
rect 387154 223207 387210 223216
rect 387062 222184 387118 222193
rect 387062 222119 387118 222128
rect 386880 220788 386932 220794
rect 386880 220730 386932 220736
rect 385776 220720 385828 220726
rect 385776 220662 385828 220668
rect 386892 219881 386920 220730
rect 386878 219872 386934 219881
rect 386878 219807 386934 219816
rect 386878 212936 386934 212945
rect 386878 212871 386934 212880
rect 386892 212566 386920 212871
rect 386880 212560 386932 212566
rect 386880 212502 386932 212508
rect 387168 211818 387196 223207
rect 387524 216640 387576 216646
rect 387524 216582 387576 216588
rect 387536 216481 387564 216582
rect 387522 216472 387578 216481
rect 387522 216407 387578 216416
rect 387156 211812 387208 211818
rect 387156 211754 387208 211760
rect 386878 209536 386934 209545
rect 386878 209471 386934 209480
rect 386892 208418 386920 209471
rect 386880 208412 386932 208418
rect 386880 208354 386932 208360
rect 386878 206136 386934 206145
rect 386878 206071 386934 206080
rect 386892 205698 386920 206071
rect 386880 205692 386932 205698
rect 386880 205634 386932 205640
rect 386878 202736 386934 202745
rect 386878 202671 386934 202680
rect 386892 202230 386920 202671
rect 386880 202224 386932 202230
rect 386880 202166 386932 202172
rect 387062 199336 387118 199345
rect 387062 199271 387118 199280
rect 386880 197328 386932 197334
rect 386880 197270 386932 197276
rect 386892 196081 386920 197270
rect 386878 196072 386934 196081
rect 386878 196007 386934 196016
rect 386420 193860 386472 193866
rect 386420 193802 386472 193808
rect 386432 193361 386460 193802
rect 386418 193352 386474 193361
rect 386418 193287 386474 193296
rect 387076 190398 387104 199271
rect 387064 190392 387116 190398
rect 387064 190334 387116 190340
rect 386878 189816 386934 189825
rect 386878 189751 386934 189760
rect 386788 187672 386840 187678
rect 386788 187614 386840 187620
rect 386800 186561 386828 187614
rect 386786 186552 386842 186561
rect 386786 186487 386842 186496
rect 386892 185638 386920 189751
rect 386880 185632 386932 185638
rect 386880 185574 386932 185580
rect 386418 183016 386474 183025
rect 386418 182951 386474 182960
rect 386432 182238 386460 182951
rect 386420 182232 386472 182238
rect 386420 182174 386472 182180
rect 386878 179616 386934 179625
rect 386878 179551 386934 179560
rect 386892 178022 386920 179551
rect 386880 178016 386932 178022
rect 386880 177958 386932 177964
rect 387628 173874 387656 284582
rect 387720 270065 387748 358022
rect 387706 270056 387762 270065
rect 387706 269991 387762 270000
rect 387800 229084 387852 229090
rect 387800 229026 387852 229032
rect 387708 228744 387760 228750
rect 387708 228686 387760 228692
rect 387156 173868 387208 173874
rect 387156 173810 387208 173816
rect 387616 173868 387668 173874
rect 387616 173810 387668 173816
rect 387168 172961 387196 173810
rect 387154 172952 387210 172961
rect 387154 172887 387210 172896
rect 386880 169720 386932 169726
rect 386880 169662 386932 169668
rect 386892 169561 386920 169662
rect 386878 169552 386934 169561
rect 386878 169487 386934 169496
rect 386880 166320 386932 166326
rect 386880 166262 386932 166268
rect 386892 166161 386920 166262
rect 386878 166152 386934 166161
rect 386878 166087 386934 166096
rect 386880 162852 386932 162858
rect 386880 162794 386932 162800
rect 386892 162761 386920 162794
rect 386878 162752 386934 162761
rect 386878 162687 386934 162696
rect 387062 159216 387118 159225
rect 387062 159151 387118 159160
rect 385776 153876 385828 153882
rect 385776 153818 385828 153824
rect 385684 143540 385736 143546
rect 385684 143482 385736 143488
rect 385684 135924 385736 135930
rect 385684 135866 385736 135872
rect 385696 95130 385724 135866
rect 385788 95402 385816 153818
rect 386880 153196 386932 153202
rect 386880 153138 386932 153144
rect 386892 152561 386920 153138
rect 386878 152552 386934 152561
rect 386878 152487 386934 152496
rect 386604 150408 386656 150414
rect 386604 150350 386656 150356
rect 386616 149161 386644 150350
rect 386602 149152 386658 149161
rect 386602 149087 386658 149096
rect 387076 146266 387104 159151
rect 387064 146260 387116 146266
rect 387064 146202 387116 146208
rect 386602 145616 386658 145625
rect 386602 145551 386658 145560
rect 386616 144974 386644 145551
rect 386604 144968 386656 144974
rect 386604 144910 386656 144916
rect 387614 142896 387670 142905
rect 387614 142831 387670 142840
rect 387628 140078 387656 142831
rect 387616 140072 387668 140078
rect 387616 140014 387668 140020
rect 387154 139496 387210 139505
rect 387154 139431 387210 139440
rect 386694 136096 386750 136105
rect 386694 136031 386750 136040
rect 386708 135998 386736 136031
rect 386420 135992 386472 135998
rect 386420 135934 386472 135940
rect 386696 135992 386748 135998
rect 386696 135934 386748 135940
rect 386432 131782 386460 135934
rect 386420 131776 386472 131782
rect 386420 131718 386472 131724
rect 386604 129736 386656 129742
rect 386604 129678 386656 129684
rect 386616 129441 386644 129678
rect 386602 129432 386658 129441
rect 386602 129367 386658 129376
rect 387064 129056 387116 129062
rect 387064 128998 387116 129004
rect 385868 123480 385920 123486
rect 385868 123422 385920 123428
rect 385776 95396 385828 95402
rect 385776 95338 385828 95344
rect 385684 95124 385736 95130
rect 385684 95066 385736 95072
rect 385880 93498 385908 123422
rect 386788 122800 386840 122806
rect 386788 122742 386840 122748
rect 386800 122641 386828 122742
rect 386786 122632 386842 122641
rect 386786 122567 386842 122576
rect 386880 120080 386932 120086
rect 386880 120022 386932 120028
rect 386892 119241 386920 120022
rect 386878 119232 386934 119241
rect 386878 119167 386934 119176
rect 386878 115696 386934 115705
rect 386878 115631 386934 115640
rect 386892 114578 386920 115631
rect 386880 114572 386932 114578
rect 386880 114514 386932 114520
rect 386602 109032 386658 109041
rect 386602 108967 386604 108976
rect 386656 108967 386658 108976
rect 386604 108938 386656 108944
rect 387076 106185 387104 128998
rect 387168 122126 387196 139431
rect 387616 133204 387668 133210
rect 387616 133146 387668 133152
rect 387628 126041 387656 133146
rect 387614 126032 387670 126041
rect 387614 125967 387670 125976
rect 387156 122120 387208 122126
rect 387156 122062 387208 122068
rect 387156 112464 387208 112470
rect 387156 112406 387208 112412
rect 387062 106176 387118 106185
rect 387062 106111 387118 106120
rect 385960 103556 386012 103562
rect 385960 103498 386012 103504
rect 385868 93492 385920 93498
rect 385868 93434 385920 93440
rect 384396 86896 384448 86902
rect 384396 86838 384448 86844
rect 381728 86828 381780 86834
rect 381728 86770 381780 86776
rect 385972 85406 386000 103498
rect 386880 99340 386932 99346
rect 386880 99282 386932 99288
rect 386892 98841 386920 99282
rect 386878 98832 386934 98841
rect 386878 98767 386934 98776
rect 387168 93566 387196 112406
rect 387248 106344 387300 106350
rect 387248 106286 387300 106292
rect 387156 93560 387208 93566
rect 387156 93502 387208 93508
rect 387260 90846 387288 106286
rect 387614 106176 387670 106185
rect 387614 106111 387670 106120
rect 387628 105641 387656 106111
rect 387614 105632 387670 105641
rect 387614 105567 387670 105576
rect 387248 90840 387300 90846
rect 387248 90782 387300 90788
rect 385960 85400 386012 85406
rect 385960 85342 386012 85348
rect 377496 82680 377548 82686
rect 377496 82622 377548 82628
rect 373448 81252 373500 81258
rect 373448 81194 373500 81200
rect 387628 60722 387656 105567
rect 387720 92342 387748 228686
rect 387812 228478 387840 229026
rect 388456 228478 388484 404330
rect 389088 349852 389140 349858
rect 389088 349794 389140 349800
rect 388996 304292 389048 304298
rect 388996 304234 389048 304240
rect 388534 277808 388590 277817
rect 388534 277743 388590 277752
rect 387800 228472 387852 228478
rect 387800 228414 387852 228420
rect 388444 228472 388496 228478
rect 388444 228414 388496 228420
rect 387812 175953 387840 228414
rect 388442 213888 388498 213897
rect 388442 213823 388498 213832
rect 387798 175944 387854 175953
rect 387798 175879 387854 175888
rect 388456 155961 388484 213823
rect 388442 155952 388498 155961
rect 388442 155887 388498 155896
rect 388444 149728 388496 149734
rect 388444 149670 388496 149676
rect 388456 92410 388484 149670
rect 388548 135250 388576 277743
rect 389008 216481 389036 304234
rect 388994 216472 389050 216481
rect 388994 216407 389050 216416
rect 388628 137284 388680 137290
rect 388628 137226 388680 137232
rect 388536 135244 388588 135250
rect 388536 135186 388588 135192
rect 388536 113824 388588 113830
rect 388536 113766 388588 113772
rect 388444 92404 388496 92410
rect 388444 92346 388496 92352
rect 387708 92336 387760 92342
rect 387708 92278 387760 92284
rect 388548 90778 388576 113766
rect 388640 94858 388668 137226
rect 389100 132841 389128 349794
rect 391216 301481 391244 576846
rect 392584 430636 392636 430642
rect 392584 430578 392636 430584
rect 391202 301472 391258 301481
rect 391202 301407 391258 301416
rect 392596 284646 392624 430578
rect 412652 303618 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 429856 700330 429884 703520
rect 429844 700324 429896 700330
rect 429844 700266 429896 700272
rect 421564 358828 421616 358834
rect 421564 358770 421616 358776
rect 415768 352572 415820 352578
rect 415768 352514 415820 352520
rect 412640 303612 412692 303618
rect 412640 303554 412692 303560
rect 413284 303612 413336 303618
rect 413284 303554 413336 303560
rect 413296 287706 413324 303554
rect 406108 287700 406160 287706
rect 406108 287642 406160 287648
rect 413284 287700 413336 287706
rect 413284 287642 413336 287648
rect 392584 284640 392636 284646
rect 392584 284582 392636 284588
rect 389916 283280 389968 283286
rect 389916 283222 389968 283228
rect 389640 280288 389692 280294
rect 389640 280230 389692 280236
rect 389652 275330 389680 280230
rect 389824 277772 389876 277778
rect 389824 277714 389876 277720
rect 389640 275324 389692 275330
rect 389640 275266 389692 275272
rect 389732 275256 389784 275262
rect 389732 275198 389784 275204
rect 389744 267034 389772 275198
rect 389732 267028 389784 267034
rect 389732 266970 389784 266976
rect 389836 162489 389864 277714
rect 389928 275262 389956 283222
rect 397092 280560 397144 280566
rect 397092 280502 397144 280508
rect 393872 279132 393924 279138
rect 393872 279074 393924 279080
rect 391940 278860 391992 278866
rect 391940 278802 391992 278808
rect 391952 276690 391980 278802
rect 391940 276684 391992 276690
rect 391940 276626 391992 276632
rect 393884 275876 393912 279074
rect 397104 275876 397132 280502
rect 403532 279064 403584 279070
rect 403532 279006 403584 279012
rect 400312 278928 400364 278934
rect 400312 278870 400364 278876
rect 400324 275876 400352 278870
rect 403544 275876 403572 279006
rect 406120 275876 406148 287642
rect 409236 280492 409288 280498
rect 409236 280434 409288 280440
rect 390466 275632 390522 275641
rect 409248 275618 409276 280434
rect 410340 276412 410392 276418
rect 410340 276354 410392 276360
rect 410352 276010 410380 276354
rect 412548 276208 412600 276214
rect 412548 276150 412600 276156
rect 410340 276004 410392 276010
rect 410340 275946 410392 275952
rect 412560 275876 412588 276150
rect 415780 275876 415808 352514
rect 418988 288584 419040 288590
rect 418988 288526 419040 288532
rect 419000 275876 419028 288526
rect 421576 278934 421604 358770
rect 435088 357536 435140 357542
rect 435088 357478 435140 357484
rect 428648 284572 428700 284578
rect 428648 284514 428700 284520
rect 425428 280356 425480 280362
rect 425428 280298 425480 280304
rect 421564 278928 421616 278934
rect 421564 278870 421616 278876
rect 421840 278928 421892 278934
rect 421840 278870 421892 278876
rect 421852 275890 421880 278870
rect 421852 275862 422234 275890
rect 425440 275876 425468 280298
rect 428660 275876 428688 284514
rect 431868 277704 431920 277710
rect 431868 277646 431920 277652
rect 431880 275876 431908 277646
rect 435100 275876 435128 357478
rect 462332 311137 462360 703520
rect 478524 700398 478552 703520
rect 494808 702545 494836 703520
rect 494794 702536 494850 702545
rect 494794 702471 494850 702480
rect 478512 700392 478564 700398
rect 478512 700334 478564 700340
rect 527192 700330 527220 703520
rect 543476 702434 543504 703520
rect 559668 702506 559696 703520
rect 559656 702500 559708 702506
rect 559656 702442 559708 702448
rect 542372 702406 543504 702434
rect 527180 700324 527232 700330
rect 527180 700266 527232 700272
rect 502984 630692 503036 630698
rect 502984 630634 503036 630640
rect 463424 361684 463476 361690
rect 463424 361626 463476 361632
rect 462318 311128 462374 311137
rect 462318 311063 462374 311072
rect 449900 289876 449952 289882
rect 449900 289818 449952 289824
rect 449912 287054 449940 289818
rect 456984 287700 457036 287706
rect 456984 287642 457036 287648
rect 449912 287026 450768 287054
rect 441528 283280 441580 283286
rect 441528 283222 441580 283228
rect 438308 281920 438360 281926
rect 438308 281862 438360 281868
rect 438320 275876 438348 281862
rect 441540 275876 441568 283222
rect 447968 278996 448020 279002
rect 447968 278938 448020 278944
rect 444746 276312 444802 276321
rect 444746 276247 444802 276256
rect 444760 275876 444788 276247
rect 447980 275876 448008 278938
rect 450740 275890 450768 287026
rect 452660 277704 452712 277710
rect 452660 277646 452712 277652
rect 450740 275862 451214 275890
rect 390522 275590 390678 275618
rect 409248 275602 409736 275618
rect 452672 275602 452700 277646
rect 453764 277636 453816 277642
rect 453764 277578 453816 277584
rect 453776 275876 453804 277578
rect 456996 275876 457024 287642
rect 460202 277808 460258 277817
rect 460202 277743 460258 277752
rect 460216 275876 460244 277743
rect 463436 275876 463464 361626
rect 498844 337408 498896 337414
rect 498844 337350 498896 337356
rect 471244 311908 471296 311914
rect 471244 311850 471296 311856
rect 468484 309800 468536 309806
rect 468484 309742 468536 309748
rect 468496 287706 468524 309742
rect 468484 287700 468536 287706
rect 468484 287642 468536 287648
rect 471256 284986 471284 311850
rect 492404 294636 492456 294642
rect 492404 294578 492456 294584
rect 486424 287700 486476 287706
rect 486424 287642 486476 287648
rect 471244 284980 471296 284986
rect 471244 284922 471296 284928
rect 473084 284504 473136 284510
rect 473084 284446 473136 284452
rect 469864 280424 469916 280430
rect 469864 280366 469916 280372
rect 466644 276344 466696 276350
rect 466644 276286 466696 276292
rect 466656 275876 466684 276286
rect 469876 275876 469904 280366
rect 473096 275876 473124 284446
rect 482744 281852 482796 281858
rect 482744 281794 482796 281800
rect 476302 279168 476358 279177
rect 476302 279103 476358 279112
rect 476316 275876 476344 279103
rect 479522 277672 479578 277681
rect 479522 277607 479578 277616
rect 479536 275876 479564 277607
rect 482756 275876 482784 281794
rect 486436 277642 486464 287642
rect 489184 277704 489236 277710
rect 489184 277646 489236 277652
rect 486424 277636 486476 277642
rect 486424 277578 486476 277584
rect 486436 277394 486464 277578
rect 486344 277366 486464 277394
rect 486344 275890 486372 277366
rect 485990 275862 486372 275890
rect 489196 275876 489224 277646
rect 492416 275876 492444 294578
rect 495624 277568 495676 277574
rect 495624 277510 495676 277516
rect 495636 275876 495664 277510
rect 498856 275876 498884 337350
rect 502996 298110 503024 630634
rect 530584 590708 530636 590714
rect 530584 590650 530636 590656
rect 520924 341556 520976 341562
rect 520924 341498 520976 341504
rect 502340 298104 502392 298110
rect 502340 298046 502392 298052
rect 502984 298104 503036 298110
rect 502984 298046 503036 298052
rect 502352 296750 502380 298046
rect 502340 296744 502392 296750
rect 520936 296714 520964 341498
rect 502340 296686 502392 296692
rect 520752 296686 520964 296714
rect 502352 278730 502380 296686
rect 520752 292602 520780 296686
rect 520740 292596 520792 292602
rect 520740 292538 520792 292544
rect 514300 285864 514352 285870
rect 514300 285806 514352 285812
rect 507860 283212 507912 283218
rect 507860 283154 507912 283160
rect 501420 278724 501472 278730
rect 501420 278666 501472 278672
rect 502340 278724 502392 278730
rect 502340 278666 502392 278672
rect 501432 275876 501460 278666
rect 507872 275876 507900 283154
rect 510802 276040 510858 276049
rect 510802 275975 510858 275984
rect 510816 275890 510844 275975
rect 510816 275862 511106 275890
rect 514312 275876 514340 285806
rect 517520 277500 517572 277506
rect 517520 277442 517572 277448
rect 517532 275876 517560 277442
rect 520752 275876 520780 292538
rect 530596 284986 530624 590650
rect 536104 484424 536156 484430
rect 536104 484366 536156 484372
rect 536116 341562 536144 484366
rect 538864 360324 538916 360330
rect 538864 360266 538916 360272
rect 536104 341556 536156 341562
rect 536104 341498 536156 341504
rect 531964 334008 532016 334014
rect 531964 333950 532016 333956
rect 531976 284986 532004 333950
rect 533620 290012 533672 290018
rect 533620 289954 533672 289960
rect 527180 284980 527232 284986
rect 527180 284922 527232 284928
rect 530584 284980 530636 284986
rect 530584 284922 530636 284928
rect 531964 284980 532016 284986
rect 531964 284922 532016 284928
rect 523960 281784 524012 281790
rect 523960 281726 524012 281732
rect 523972 275876 524000 281726
rect 527192 275876 527220 284922
rect 530400 276276 530452 276282
rect 530400 276218 530452 276224
rect 530412 275876 530440 276218
rect 533632 275876 533660 289954
rect 536840 285796 536892 285802
rect 536840 285738 536892 285744
rect 536852 275876 536880 285738
rect 538876 278730 538904 360266
rect 542372 304298 542400 702406
rect 559668 700398 559696 702442
rect 559656 700392 559708 700398
rect 559656 700334 559708 700340
rect 582380 700392 582432 700398
rect 582380 700334 582432 700340
rect 565820 700324 565872 700330
rect 565820 700266 565872 700272
rect 561956 367124 562008 367130
rect 561956 367066 562008 367072
rect 552294 355328 552350 355337
rect 552294 355263 552350 355272
rect 542360 304292 542412 304298
rect 542360 304234 542412 304240
rect 546500 284980 546552 284986
rect 546500 284922 546552 284928
rect 540058 279032 540114 279041
rect 540058 278967 540114 278976
rect 538864 278724 538916 278730
rect 538864 278666 538916 278672
rect 540072 275876 540100 278967
rect 543280 278724 543332 278730
rect 543280 278666 543332 278672
rect 543292 275876 543320 278666
rect 546512 275876 546540 284922
rect 549076 277772 549128 277778
rect 549076 277714 549128 277720
rect 549088 275876 549116 277714
rect 552308 275876 552336 355263
rect 555516 283008 555568 283014
rect 555516 282950 555568 282956
rect 555528 275876 555556 282950
rect 558734 277536 558790 277545
rect 558734 277471 558790 277480
rect 558748 275876 558776 277471
rect 561968 275876 561996 367066
rect 563704 361616 563756 361622
rect 563704 361558 563756 361564
rect 563716 278730 563744 361558
rect 565832 284889 565860 700266
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 567844 683188 567896 683194
rect 567844 683130 567896 683136
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 566464 291236 566516 291242
rect 566464 291178 566516 291184
rect 565818 284880 565874 284889
rect 565818 284815 565874 284824
rect 563704 278724 563756 278730
rect 563704 278666 563756 278672
rect 565176 278724 565228 278730
rect 565176 278666 565228 278672
rect 565188 275876 565216 278666
rect 566476 277098 566504 291178
rect 566556 288516 566608 288522
rect 566556 288458 566608 288464
rect 566464 277092 566516 277098
rect 566464 277034 566516 277040
rect 566568 276690 566596 288458
rect 567856 281722 567884 683130
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 574744 643136 574796 643142
rect 574744 643078 574796 643084
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 573364 458856 573416 458862
rect 573364 458798 573416 458804
rect 571432 365764 571484 365770
rect 571432 365706 571484 365712
rect 570512 364404 570564 364410
rect 570512 364346 570564 364352
rect 570524 358086 570552 364346
rect 570512 358080 570564 358086
rect 570512 358022 570564 358028
rect 568578 354784 568634 354793
rect 568578 354719 568634 354728
rect 567844 281716 567896 281722
rect 567844 281658 567896 281664
rect 568396 281716 568448 281722
rect 568396 281658 568448 281664
rect 566556 276684 566608 276690
rect 566556 276626 566608 276632
rect 568408 275876 568436 281658
rect 568592 278769 568620 354719
rect 570052 313948 570104 313954
rect 570052 313890 570104 313896
rect 569960 282940 570012 282946
rect 569960 282882 570012 282888
rect 568578 278760 568634 278769
rect 568578 278695 568634 278704
rect 568672 277092 568724 277098
rect 568672 277034 568724 277040
rect 504362 275632 504418 275641
rect 409248 275596 409748 275602
rect 409248 275590 409696 275596
rect 390466 275567 390522 275576
rect 409696 275538 409748 275544
rect 452660 275596 452712 275602
rect 504418 275590 504666 275618
rect 504362 275567 504418 275576
rect 452660 275538 452712 275544
rect 389916 275256 389968 275262
rect 389916 275198 389968 275204
rect 568578 274952 568634 274961
rect 568578 274887 568634 274896
rect 568592 229094 568620 274887
rect 568684 267734 568712 277034
rect 568684 267706 569356 267734
rect 569328 257689 569356 267706
rect 569972 264625 570000 282882
rect 569958 264616 570014 264625
rect 569958 264551 570014 264560
rect 569314 257680 569370 257689
rect 569314 257615 569370 257624
rect 569958 237280 570014 237289
rect 569958 237215 570014 237224
rect 568592 229066 569356 229094
rect 569328 220833 569356 229066
rect 569314 220824 569370 220833
rect 569314 220759 569370 220768
rect 389822 162480 389878 162489
rect 389822 162415 389878 162424
rect 569314 156088 569370 156097
rect 569314 156023 569370 156032
rect 569328 142154 569356 156023
rect 568592 142126 569356 142154
rect 389086 132832 389142 132841
rect 389086 132767 389142 132776
rect 389824 124908 389876 124914
rect 389824 124850 389876 124856
rect 388720 111104 388772 111110
rect 388720 111046 388772 111052
rect 388732 95198 388760 111046
rect 389732 105596 389784 105602
rect 389732 105538 389784 105544
rect 389640 96824 389692 96830
rect 389640 96766 389692 96772
rect 388720 95192 388772 95198
rect 388720 95134 388772 95140
rect 388628 94852 388680 94858
rect 388628 94794 388680 94800
rect 389652 93809 389680 96766
rect 389744 96506 389772 105538
rect 389836 96830 389864 124850
rect 389824 96824 389876 96830
rect 389824 96766 389876 96772
rect 568592 96558 568620 142126
rect 569224 126268 569276 126274
rect 569224 126210 569276 126216
rect 568580 96552 568632 96558
rect 389744 96478 390034 96506
rect 568580 96494 568632 96500
rect 392596 95470 392624 96084
rect 392584 95464 392636 95470
rect 392584 95406 392636 95412
rect 395816 95130 395844 96084
rect 399036 95198 399064 96084
rect 399024 95192 399076 95198
rect 399024 95134 399076 95140
rect 395804 95124 395856 95130
rect 395804 95066 395856 95072
rect 389638 93800 389694 93809
rect 389638 93735 389694 93744
rect 402256 93634 402284 96084
rect 402244 93628 402296 93634
rect 402244 93570 402296 93576
rect 405476 92449 405504 96084
rect 405462 92440 405518 92449
rect 405462 92375 405518 92384
rect 408696 91089 408724 96084
rect 411916 93498 411944 96084
rect 415136 93566 415164 96084
rect 418356 95130 418384 96084
rect 418344 95124 418396 95130
rect 418344 95066 418396 95072
rect 415124 93560 415176 93566
rect 415124 93502 415176 93508
rect 411904 93492 411956 93498
rect 411904 93434 411956 93440
rect 418356 92206 418384 95066
rect 421576 94858 421604 96084
rect 424796 95062 424824 96084
rect 428016 95402 428044 96084
rect 428004 95396 428056 95402
rect 428004 95338 428056 95344
rect 424784 95056 424836 95062
rect 424784 94998 424836 95004
rect 421564 94852 421616 94858
rect 421564 94794 421616 94800
rect 418344 92200 418396 92206
rect 418344 92142 418396 92148
rect 431236 91798 431264 96084
rect 430488 91792 430540 91798
rect 430488 91734 430540 91740
rect 431224 91792 431276 91798
rect 431224 91734 431276 91740
rect 408682 91080 408738 91089
rect 408682 91015 408738 91024
rect 388536 90772 388588 90778
rect 388536 90714 388588 90720
rect 430500 89554 430528 91734
rect 434456 90846 434484 96084
rect 437032 94994 437060 96084
rect 437020 94988 437072 94994
rect 437020 94930 437072 94936
rect 434444 90840 434496 90846
rect 434444 90782 434496 90788
rect 429200 89548 429252 89554
rect 429200 89490 429252 89496
rect 430488 89548 430540 89554
rect 430488 89490 430540 89496
rect 429212 88330 429240 89490
rect 440252 89418 440280 96084
rect 443472 93770 443500 96084
rect 443460 93764 443512 93770
rect 443460 93706 443512 93712
rect 446692 92138 446720 96084
rect 449912 92206 449940 96084
rect 452672 96070 453146 96098
rect 449900 92200 449952 92206
rect 449900 92142 449952 92148
rect 446680 92132 446732 92138
rect 446680 92074 446732 92080
rect 440240 89412 440292 89418
rect 440240 89354 440292 89360
rect 429200 88324 429252 88330
rect 429200 88266 429252 88272
rect 452672 85338 452700 96070
rect 456352 93770 456380 96084
rect 456340 93764 456392 93770
rect 456340 93706 456392 93712
rect 459572 88194 459600 96084
rect 459560 88188 459612 88194
rect 459560 88130 459612 88136
rect 462792 88126 462820 96084
rect 465092 96070 466026 96098
rect 462780 88120 462832 88126
rect 462780 88062 462832 88068
rect 465092 86834 465120 96070
rect 469232 90982 469260 96084
rect 469220 90976 469272 90982
rect 469220 90918 469272 90924
rect 472452 90778 472480 96084
rect 475672 93702 475700 96084
rect 475660 93696 475712 93702
rect 475660 93638 475712 93644
rect 478892 90914 478920 96084
rect 478880 90908 478932 90914
rect 478880 90850 478932 90856
rect 472440 90772 472492 90778
rect 472440 90714 472492 90720
rect 482112 89486 482140 96084
rect 484412 96070 484702 96098
rect 487816 96070 487922 96098
rect 489932 96070 491142 96098
rect 494072 96070 494362 96098
rect 496832 96070 497582 96098
rect 482100 89480 482152 89486
rect 482100 89422 482152 89428
rect 465080 86828 465132 86834
rect 465080 86770 465132 86776
rect 452660 85332 452712 85338
rect 452660 85274 452712 85280
rect 484412 77246 484440 96070
rect 487816 93702 487844 96070
rect 487804 93696 487856 93702
rect 487804 93638 487856 93644
rect 487816 85474 487844 93638
rect 489932 86902 489960 96070
rect 489920 86896 489972 86902
rect 489920 86838 489972 86844
rect 487804 85468 487856 85474
rect 487804 85410 487856 85416
rect 494072 82686 494100 96070
rect 496832 85406 496860 96070
rect 500788 95334 500816 96084
rect 503732 96070 504022 96098
rect 500776 95328 500828 95334
rect 500776 95270 500828 95276
rect 496820 85400 496872 85406
rect 496820 85342 496872 85348
rect 503732 82754 503760 96070
rect 507228 95266 507256 96084
rect 509896 96070 510462 96098
rect 507216 95260 507268 95266
rect 507216 95202 507268 95208
rect 509896 92274 509924 96070
rect 513668 94926 513696 96084
rect 516152 96070 516902 96098
rect 518912 96070 520122 96098
rect 513656 94920 513708 94926
rect 513656 94862 513708 94868
rect 509884 92268 509936 92274
rect 509884 92210 509936 92216
rect 510528 92268 510580 92274
rect 510528 92210 510580 92216
rect 510540 84862 510568 92210
rect 510528 84856 510580 84862
rect 510528 84798 510580 84804
rect 516152 84114 516180 96070
rect 516140 84108 516192 84114
rect 516140 84050 516192 84056
rect 503720 82748 503772 82754
rect 503720 82690 503772 82696
rect 494060 82680 494112 82686
rect 494060 82622 494112 82628
rect 518912 81326 518940 96070
rect 523328 95266 523356 96084
rect 523316 95260 523368 95266
rect 523316 95202 523368 95208
rect 526548 89622 526576 96084
rect 529768 93634 529796 96084
rect 531332 96070 532358 96098
rect 535472 96070 535578 96098
rect 529756 93628 529808 93634
rect 529756 93570 529808 93576
rect 526536 89616 526588 89622
rect 526536 89558 526588 89564
rect 531332 85542 531360 96070
rect 535472 86873 535500 96070
rect 538784 93673 538812 96084
rect 542004 95062 542032 96084
rect 545132 96070 545238 96098
rect 541992 95056 542044 95062
rect 541992 94998 542044 95004
rect 538770 93664 538826 93673
rect 538770 93599 538826 93608
rect 535458 86864 535514 86873
rect 535458 86799 535514 86808
rect 531320 85536 531372 85542
rect 531320 85478 531372 85484
rect 522304 84856 522356 84862
rect 522304 84798 522356 84804
rect 518900 81320 518952 81326
rect 518900 81262 518952 81268
rect 484400 77240 484452 77246
rect 484400 77182 484452 77188
rect 387616 60716 387668 60722
rect 387616 60658 387668 60664
rect 373264 59356 373316 59362
rect 373264 59298 373316 59304
rect 522316 33114 522344 84798
rect 545132 77178 545160 96070
rect 548444 95198 548472 96084
rect 550652 96070 551678 96098
rect 548432 95192 548484 95198
rect 548432 95134 548484 95140
rect 548444 93854 548472 95134
rect 548444 93826 548564 93854
rect 548536 82822 548564 93826
rect 548524 82816 548576 82822
rect 548524 82758 548576 82764
rect 550652 81258 550680 96070
rect 554884 89690 554912 96084
rect 557552 96070 558118 96098
rect 560312 96070 561338 96098
rect 554872 89684 554924 89690
rect 554872 89626 554924 89632
rect 557552 84182 557580 96070
rect 560312 86970 560340 96070
rect 564544 93838 564572 96084
rect 564532 93832 564584 93838
rect 564532 93774 564584 93780
rect 567764 93566 567792 96084
rect 569236 95062 569264 126210
rect 569314 97200 569370 97209
rect 569314 97135 569370 97144
rect 569224 95056 569276 95062
rect 569224 94998 569276 95004
rect 569328 93634 569356 97135
rect 569316 93628 569368 93634
rect 569316 93570 569368 93576
rect 567752 93560 567804 93566
rect 567752 93502 567804 93508
rect 569972 91050 570000 237215
rect 570064 106865 570092 313890
rect 570236 307828 570288 307834
rect 570236 307770 570288 307776
rect 570144 276140 570196 276146
rect 570144 276082 570196 276088
rect 570156 223961 570184 276082
rect 570142 223952 570198 223961
rect 570142 223887 570198 223896
rect 570248 217161 570276 307770
rect 571340 276072 571392 276078
rect 571340 276014 571392 276020
rect 570234 217152 570290 217161
rect 570234 217087 570290 217096
rect 570142 180296 570198 180305
rect 570142 180231 570198 180240
rect 570050 106856 570106 106865
rect 570050 106791 570106 106800
rect 570050 99512 570106 99521
rect 570050 99447 570106 99456
rect 569960 91044 570012 91050
rect 569960 90986 570012 90992
rect 560300 86964 560352 86970
rect 560300 86906 560352 86912
rect 557540 84176 557592 84182
rect 557540 84118 557592 84124
rect 550640 81252 550692 81258
rect 550640 81194 550692 81200
rect 570064 78674 570092 99447
rect 570156 80034 570184 180231
rect 571352 163441 571380 276014
rect 571444 253881 571472 365706
rect 571616 287156 571668 287162
rect 571616 287098 571668 287104
rect 571524 276684 571576 276690
rect 571524 276626 571576 276632
rect 571536 267481 571564 276626
rect 571628 270881 571656 287098
rect 572718 274816 572774 274825
rect 572718 274751 572774 274760
rect 571614 270872 571670 270881
rect 571614 270807 571670 270816
rect 571522 267472 571578 267481
rect 571522 267407 571578 267416
rect 572628 260840 572680 260846
rect 572628 260782 572680 260788
rect 572640 260681 572668 260782
rect 572626 260672 572682 260681
rect 572626 260607 572682 260616
rect 571430 253872 571486 253881
rect 571430 253807 571486 253816
rect 572628 251184 572680 251190
rect 572626 251152 572628 251161
rect 572680 251152 572682 251161
rect 572626 251087 572682 251096
rect 572628 248260 572680 248266
rect 572628 248202 572680 248208
rect 572640 247761 572668 248202
rect 572626 247752 572682 247761
rect 572626 247687 572682 247696
rect 572628 241460 572680 241466
rect 572628 241402 572680 241408
rect 572640 240961 572668 241402
rect 572626 240952 572682 240961
rect 572626 240887 572682 240896
rect 572628 234592 572680 234598
rect 572628 234534 572680 234540
rect 572640 234161 572668 234534
rect 572626 234152 572682 234161
rect 572626 234087 572682 234096
rect 572626 230752 572682 230761
rect 572732 230738 572760 274751
rect 572682 230710 572760 230738
rect 572626 230687 572682 230696
rect 572628 227384 572680 227390
rect 572626 227352 572628 227361
rect 572680 227352 572682 227361
rect 572626 227287 572682 227296
rect 572626 213616 572682 213625
rect 572626 213551 572682 213560
rect 572640 212566 572668 213551
rect 572628 212560 572680 212566
rect 572628 212502 572680 212508
rect 572628 211132 572680 211138
rect 572628 211074 572680 211080
rect 572640 210361 572668 211074
rect 572626 210352 572682 210361
rect 572626 210287 572682 210296
rect 572444 206984 572496 206990
rect 572442 206952 572444 206961
rect 572496 206952 572498 206961
rect 572442 206887 572498 206896
rect 571524 203924 571576 203930
rect 571524 203866 571576 203872
rect 571536 203561 571564 203866
rect 571522 203552 571578 203561
rect 571522 203487 571578 203496
rect 572628 198688 572680 198694
rect 572628 198630 572680 198636
rect 572640 197441 572668 198630
rect 572626 197432 572682 197441
rect 572626 197367 572682 197376
rect 571708 191752 571760 191758
rect 571708 191694 571760 191700
rect 571720 190641 571748 191694
rect 571706 190632 571762 190641
rect 571706 190567 571762 190576
rect 572628 187672 572680 187678
rect 572628 187614 572680 187620
rect 572640 187241 572668 187614
rect 572626 187232 572682 187241
rect 572626 187167 572682 187176
rect 571432 184884 571484 184890
rect 571432 184826 571484 184832
rect 571444 183841 571472 184826
rect 571430 183832 571486 183841
rect 571430 183767 571486 183776
rect 572076 178016 572128 178022
rect 572076 177958 572128 177964
rect 572088 177041 572116 177958
rect 572074 177032 572130 177041
rect 572074 176967 572130 176976
rect 572626 170096 572682 170105
rect 572626 170031 572682 170040
rect 572640 169794 572668 170031
rect 572628 169788 572680 169794
rect 572628 169730 572680 169736
rect 572350 166696 572406 166705
rect 572350 166631 572406 166640
rect 572364 165646 572392 166631
rect 572352 165640 572404 165646
rect 572352 165582 572404 165588
rect 571338 163432 571394 163441
rect 571338 163367 571394 163376
rect 572626 159896 572682 159905
rect 572626 159831 572682 159840
rect 572640 158778 572668 159831
rect 572628 158772 572680 158778
rect 572628 158714 572680 158720
rect 572628 153264 572680 153270
rect 572626 153232 572628 153241
rect 572680 153232 572682 153241
rect 572626 153167 572682 153176
rect 572628 151088 572680 151094
rect 572628 151030 572680 151036
rect 572640 150521 572668 151030
rect 572626 150512 572682 150521
rect 572626 150447 572682 150456
rect 571708 147348 571760 147354
rect 571708 147290 571760 147296
rect 571720 147121 571748 147290
rect 571706 147112 571762 147121
rect 571706 147047 571762 147056
rect 572628 143608 572680 143614
rect 572626 143576 572628 143585
rect 572680 143576 572682 143585
rect 572626 143511 572682 143520
rect 572626 140176 572682 140185
rect 572626 140111 572682 140120
rect 572640 139466 572668 140111
rect 572628 139460 572680 139466
rect 572628 139402 572680 139408
rect 572628 137964 572680 137970
rect 572628 137906 572680 137912
rect 572640 136921 572668 137906
rect 572626 136912 572682 136921
rect 572626 136847 572682 136856
rect 572718 133376 572774 133385
rect 572718 133311 572774 133320
rect 572628 130212 572680 130218
rect 572628 130154 572680 130160
rect 572640 130121 572668 130154
rect 572626 130112 572682 130121
rect 572626 130047 572682 130056
rect 571338 126576 571394 126585
rect 571338 126511 571394 126520
rect 570604 111852 570656 111858
rect 570604 111794 570656 111800
rect 570616 92342 570644 111794
rect 571248 106344 571300 106350
rect 571246 106312 571248 106321
rect 571300 106312 571302 106321
rect 571246 106247 571302 106256
rect 571352 96257 571380 126511
rect 572628 124160 572680 124166
rect 572628 124102 572680 124108
rect 572640 123321 572668 124102
rect 572626 123312 572682 123321
rect 572626 123247 572682 123256
rect 571430 119776 571486 119785
rect 571430 119711 571486 119720
rect 571338 96248 571394 96257
rect 571338 96183 571394 96192
rect 571444 92410 571472 119711
rect 572628 117292 572680 117298
rect 572628 117234 572680 117240
rect 572640 116521 572668 117234
rect 572626 116512 572682 116521
rect 572626 116447 572682 116456
rect 571522 112976 571578 112985
rect 571522 112911 571578 112920
rect 571536 93809 571564 112911
rect 572626 102776 572682 102785
rect 572626 102711 572682 102720
rect 572640 102202 572668 102711
rect 572628 102196 572680 102202
rect 572628 102138 572680 102144
rect 571614 96656 571670 96665
rect 571614 96591 571670 96600
rect 571522 93800 571578 93809
rect 571522 93735 571578 93744
rect 571432 92404 571484 92410
rect 571432 92346 571484 92352
rect 570604 92336 570656 92342
rect 570604 92278 570656 92284
rect 571628 88262 571656 96591
rect 572732 93430 572760 133311
rect 573376 93702 573404 458798
rect 574100 377460 574152 377466
rect 574100 377402 574152 377408
rect 574112 376786 574140 377402
rect 574100 376780 574152 376786
rect 574100 376722 574152 376728
rect 573548 324352 573600 324358
rect 573548 324294 573600 324300
rect 573560 282946 573588 324294
rect 573548 282940 573600 282946
rect 573548 282882 573600 282888
rect 573456 280356 573508 280362
rect 573456 280298 573508 280304
rect 573364 93696 573416 93702
rect 573364 93638 573416 93644
rect 572720 93424 572772 93430
rect 572720 93366 572772 93372
rect 571616 88256 571668 88262
rect 571616 88198 571668 88204
rect 573468 86970 573496 280298
rect 574112 184890 574140 376722
rect 574756 283830 574784 643078
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 576124 536852 576176 536858
rect 576124 536794 576176 536800
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 575572 327140 575624 327146
rect 575572 327082 575624 327088
rect 575480 284436 575532 284442
rect 575480 284378 575532 284384
rect 574284 283824 574336 283830
rect 574284 283766 574336 283772
rect 574744 283824 574796 283830
rect 574744 283766 574796 283772
rect 574296 283150 574324 283766
rect 574284 283144 574336 283150
rect 574284 283086 574336 283092
rect 574192 280288 574244 280294
rect 574192 280230 574244 280236
rect 574204 191758 574232 280230
rect 574296 203930 574324 283086
rect 575492 206990 575520 284378
rect 575584 260778 575612 327082
rect 575572 260772 575624 260778
rect 575572 260714 575624 260720
rect 575480 206984 575532 206990
rect 575480 206926 575532 206932
rect 574284 203924 574336 203930
rect 574284 203866 574336 203872
rect 574192 191752 574244 191758
rect 574192 191694 574244 191700
rect 574100 184884 574152 184890
rect 574100 184826 574152 184832
rect 574100 165640 574152 165646
rect 574100 165582 574152 165588
rect 574112 96529 574140 165582
rect 575480 158772 575532 158778
rect 575480 158714 575532 158720
rect 574744 155236 574796 155242
rect 574744 155178 574796 155184
rect 574756 147354 574784 155178
rect 575388 153876 575440 153882
rect 575388 153818 575440 153824
rect 575400 153270 575428 153818
rect 575388 153264 575440 153270
rect 575388 153206 575440 153212
rect 574744 147348 574796 147354
rect 574744 147290 574796 147296
rect 574744 138032 574796 138038
rect 574744 137974 574796 137980
rect 574192 102196 574244 102202
rect 574192 102138 574244 102144
rect 574098 96520 574154 96529
rect 574098 96455 574154 96464
rect 573456 86964 573508 86970
rect 573456 86906 573508 86912
rect 570144 80028 570196 80034
rect 570144 79970 570196 79976
rect 574204 79966 574232 102138
rect 574756 95130 574784 137974
rect 575400 106962 575428 153206
rect 575388 106956 575440 106962
rect 575388 106898 575440 106904
rect 574836 106344 574888 106350
rect 574836 106286 574888 106292
rect 574744 95124 574796 95130
rect 574744 95066 574796 95072
rect 574192 79960 574244 79966
rect 574192 79902 574244 79908
rect 570052 78668 570104 78674
rect 570052 78610 570104 78616
rect 545120 77172 545172 77178
rect 545120 77114 545172 77120
rect 574848 73166 574876 106286
rect 575492 95033 575520 158714
rect 575572 143608 575624 143614
rect 575572 143550 575624 143556
rect 575584 96626 575612 143550
rect 575572 96620 575624 96626
rect 575572 96562 575624 96568
rect 576136 95198 576164 536794
rect 580262 524512 580318 524521
rect 580262 524447 580318 524456
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 580184 470626 580212 471407
rect 580172 470620 580224 470626
rect 580172 470562 580224 470568
rect 580276 458862 580304 524447
rect 580264 458856 580316 458862
rect 580264 458798 580316 458804
rect 578882 458144 578938 458153
rect 578882 458079 578938 458088
rect 577504 418192 577556 418198
rect 577504 418134 577556 418140
rect 577516 281654 577544 418134
rect 578896 368558 578924 458079
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 579618 418296 579674 418305
rect 579618 418231 579674 418240
rect 579632 418198 579660 418231
rect 579620 418192 579672 418198
rect 579620 418134 579672 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 377466 580212 378383
rect 580172 377460 580224 377466
rect 580172 377402 580224 377408
rect 578240 368552 578292 368558
rect 578240 368494 578292 368500
rect 578884 368552 578936 368558
rect 578884 368494 578936 368500
rect 576952 281648 577004 281654
rect 576952 281590 577004 281596
rect 577504 281648 577556 281654
rect 577504 281590 577556 281596
rect 576858 280392 576914 280401
rect 576858 280327 576914 280336
rect 576216 277636 576268 277642
rect 576216 277578 576268 277584
rect 576228 219434 576256 277578
rect 576308 260772 576360 260778
rect 576308 260714 576360 260720
rect 576320 258738 576348 260714
rect 576308 258732 576360 258738
rect 576308 258674 576360 258680
rect 576216 219428 576268 219434
rect 576216 219370 576268 219376
rect 576216 205692 576268 205698
rect 576216 205634 576268 205640
rect 576124 95192 576176 95198
rect 576124 95134 576176 95140
rect 575478 95024 575534 95033
rect 575478 94959 575534 94968
rect 576228 92206 576256 205634
rect 576320 178022 576348 258674
rect 576872 227390 576900 280327
rect 576964 248266 576992 281590
rect 577596 278724 577648 278730
rect 577596 278666 577648 278672
rect 576952 248260 577004 248266
rect 576952 248202 577004 248208
rect 577504 244316 577556 244322
rect 577504 244258 577556 244264
rect 576860 227384 576912 227390
rect 576860 227326 576912 227332
rect 576308 178016 576360 178022
rect 576308 177958 576360 177964
rect 576860 169788 576912 169794
rect 576860 169730 576912 169736
rect 576872 92478 576900 169730
rect 576860 92472 576912 92478
rect 576860 92414 576912 92420
rect 576216 92200 576268 92206
rect 576216 92142 576268 92148
rect 577516 90982 577544 244258
rect 577608 130218 577636 278666
rect 577596 130212 577648 130218
rect 577596 130154 577648 130160
rect 578252 95266 578280 368494
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580184 364410 580212 365055
rect 580172 364404 580224 364410
rect 580172 364346 580224 364352
rect 580356 362976 580408 362982
rect 580356 362918 580408 362924
rect 578332 360256 578384 360262
rect 578332 360198 578384 360204
rect 578344 126274 578372 360198
rect 580262 354512 580318 354521
rect 580262 354447 580318 354456
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 324358 580212 325207
rect 580172 324352 580224 324358
rect 580172 324294 580224 324300
rect 580276 312089 580304 354447
rect 580368 351937 580396 362918
rect 580354 351928 580410 351937
rect 580354 351863 580410 351872
rect 580368 349858 580396 351863
rect 580356 349852 580408 349858
rect 580356 349794 580408 349800
rect 580262 312080 580318 312089
rect 580262 312015 580318 312024
rect 579618 298752 579674 298761
rect 579618 298687 579674 298696
rect 579632 294545 579660 298687
rect 579618 294536 579674 294545
rect 579618 294471 579674 294480
rect 579618 278896 579674 278905
rect 579618 278831 579674 278840
rect 579632 151094 579660 278831
rect 580276 278730 580304 312015
rect 581184 283076 581236 283082
rect 581184 283018 581236 283024
rect 580998 280528 581054 280537
rect 580998 280463 581054 280472
rect 580448 278860 580500 278866
rect 580448 278802 580500 278808
rect 580264 278724 580316 278730
rect 580264 278666 580316 278672
rect 579710 276176 579766 276185
rect 579710 276111 579766 276120
rect 579724 198694 579752 276111
rect 580172 275324 580224 275330
rect 580172 275266 580224 275272
rect 580184 272241 580212 275266
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580184 258738 580212 258839
rect 580172 258732 580224 258738
rect 580172 258674 580224 258680
rect 580080 219428 580132 219434
rect 580080 219370 580132 219376
rect 580092 219065 580120 219370
rect 580078 219056 580134 219065
rect 580078 218991 580134 219000
rect 579712 198688 579764 198694
rect 579712 198630 579764 198636
rect 580354 192536 580410 192545
rect 580354 192471 580410 192480
rect 580368 155242 580396 192471
rect 580460 179217 580488 278802
rect 580906 205728 580962 205737
rect 580906 205663 580908 205672
rect 580960 205663 580962 205672
rect 580908 205634 580960 205640
rect 580446 179208 580502 179217
rect 580446 179143 580502 179152
rect 580356 155236 580408 155242
rect 580356 155178 580408 155184
rect 581012 153882 581040 280463
rect 581092 280220 581144 280226
rect 581092 280162 581144 280168
rect 581104 234598 581132 280162
rect 581196 260846 581224 283018
rect 581644 278928 581696 278934
rect 581644 278870 581696 278876
rect 581184 260840 581236 260846
rect 581184 260782 581236 260788
rect 581092 234592 581144 234598
rect 581092 234534 581144 234540
rect 581000 153876 581052 153882
rect 581000 153818 581052 153824
rect 581656 152697 581684 278870
rect 581642 152688 581698 152697
rect 581642 152623 581698 152632
rect 579620 151088 579672 151094
rect 579620 151030 579672 151036
rect 579632 150482 579660 151030
rect 579620 150476 579672 150482
rect 579620 150418 579672 150424
rect 580264 150476 580316 150482
rect 580264 150418 580316 150424
rect 580170 139360 580226 139369
rect 580170 139295 580226 139304
rect 580184 138038 580212 139295
rect 580172 138032 580224 138038
rect 580172 137974 580224 137980
rect 578332 126268 578384 126274
rect 578332 126210 578384 126216
rect 579620 126268 579672 126274
rect 579620 126210 579672 126216
rect 579632 126041 579660 126210
rect 579618 126032 579674 126041
rect 579618 125967 579674 125976
rect 579894 112840 579950 112849
rect 579894 112775 579950 112784
rect 579908 111858 579936 112775
rect 579896 111852 579948 111858
rect 579896 111794 579948 111800
rect 578240 95260 578292 95266
rect 578240 95202 578292 95208
rect 577504 90976 577556 90982
rect 577504 90918 577556 90924
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 574836 73160 574888 73166
rect 574836 73102 574888 73108
rect 579988 73160 580040 73166
rect 579988 73102 580040 73108
rect 580000 73001 580028 73102
rect 579986 72992 580042 73001
rect 579986 72927 580042 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580170 33144 580226 33153
rect 522304 33108 522356 33114
rect 580170 33079 580172 33088
rect 522304 33050 522356 33056
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 579618 15872 579674 15881
rect 579618 15807 579674 15816
rect 351920 2984 351972 2990
rect 351920 2926 351972 2932
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579632 354 579660 15807
rect 580276 6633 580304 150418
rect 580356 106956 580408 106962
rect 580356 106898 580408 106904
rect 580368 99521 580396 106898
rect 580354 99512 580410 99521
rect 580354 99447 580410 99456
rect 582392 93770 582420 700334
rect 582562 697232 582618 697241
rect 582562 697167 582618 697176
rect 582576 281625 582604 697167
rect 582654 670712 582710 670721
rect 582654 670647 582710 670656
rect 582562 281616 582618 281625
rect 582472 281580 582524 281586
rect 582562 281551 582618 281560
rect 582472 281522 582524 281528
rect 582484 251190 582512 281522
rect 582472 251184 582524 251190
rect 582472 251126 582524 251132
rect 582576 241466 582604 281551
rect 582668 281489 582696 670647
rect 582746 617536 582802 617545
rect 582746 617471 582802 617480
rect 582760 285734 582788 617471
rect 583850 563816 583906 563825
rect 583850 563751 583906 563760
rect 583024 369912 583076 369918
rect 583024 369854 583076 369860
rect 582840 356108 582892 356114
rect 582840 356050 582892 356056
rect 582748 285728 582800 285734
rect 582748 285670 582800 285676
rect 582654 281480 582710 281489
rect 582654 281415 582710 281424
rect 582656 276412 582708 276418
rect 582656 276354 582708 276360
rect 582564 241460 582616 241466
rect 582564 241402 582616 241408
rect 582668 165889 582696 276354
rect 582760 245614 582788 245645
rect 582748 245608 582800 245614
rect 582746 245576 582748 245585
rect 582800 245576 582802 245585
rect 582746 245511 582802 245520
rect 582760 244322 582788 245511
rect 582748 244316 582800 244322
rect 582748 244258 582800 244264
rect 582748 212560 582800 212566
rect 582748 212502 582800 212508
rect 582654 165880 582710 165889
rect 582654 165815 582710 165824
rect 582656 139460 582708 139466
rect 582656 139402 582708 139408
rect 582668 95169 582696 139402
rect 582654 95160 582710 95169
rect 582654 95095 582710 95104
rect 582380 93764 582432 93770
rect 582380 93706 582432 93712
rect 582760 81394 582788 212502
rect 582852 93566 582880 356050
rect 582932 336048 582984 336054
rect 582932 335990 582984 335996
rect 582944 93838 582972 335990
rect 583036 137970 583064 369854
rect 583864 296714 583892 563751
rect 583680 296686 583892 296714
rect 583680 291122 583708 296686
rect 583864 291378 583984 291394
rect 583852 291372 583984 291378
rect 583904 291366 583984 291372
rect 583852 291314 583904 291320
rect 583680 291094 583892 291122
rect 583668 289944 583720 289950
rect 583668 289886 583720 289892
rect 583576 288448 583628 288454
rect 583576 288390 583628 288396
rect 583116 287088 583168 287094
rect 583116 287030 583168 287036
rect 583128 205737 583156 287030
rect 583300 285728 583352 285734
rect 583300 285670 583352 285676
rect 583206 281480 583262 281489
rect 583206 281415 583262 281424
rect 583220 280265 583248 281415
rect 583206 280256 583262 280265
rect 583206 280191 583262 280200
rect 583114 205728 583170 205737
rect 583114 205663 583170 205672
rect 583024 137964 583076 137970
rect 583024 137906 583076 137912
rect 583220 117298 583248 280191
rect 583312 124166 583340 285670
rect 583484 284368 583536 284374
rect 583484 284310 583536 284316
rect 583392 278792 583444 278798
rect 583392 278734 583444 278740
rect 583404 232393 583432 278734
rect 583390 232384 583446 232393
rect 583390 232319 583446 232328
rect 583496 187678 583524 284310
rect 583588 211138 583616 288390
rect 583680 245614 583708 289886
rect 583760 278996 583812 279002
rect 583760 278938 583812 278944
rect 583668 245608 583720 245614
rect 583668 245550 583720 245556
rect 583576 211132 583628 211138
rect 583576 211074 583628 211080
rect 583772 195242 583800 278938
rect 583588 195214 583800 195242
rect 583588 190454 583616 195214
rect 583864 193186 583892 291094
rect 583852 193180 583904 193186
rect 583852 193122 583904 193128
rect 583850 193080 583906 193089
rect 583956 193066 583984 291366
rect 583906 193038 583984 193066
rect 583850 193015 583906 193024
rect 583852 192976 583904 192982
rect 583852 192918 583904 192924
rect 583588 190426 583800 190454
rect 583484 187672 583536 187678
rect 583484 187614 583536 187620
rect 583300 124160 583352 124166
rect 583300 124102 583352 124108
rect 583208 117292 583260 117298
rect 583208 117234 583260 117240
rect 582932 93832 582984 93838
rect 582932 93774 582984 93780
rect 582840 93560 582892 93566
rect 582840 93502 582892 93508
rect 582748 81388 582800 81394
rect 582748 81330 582800 81336
rect 583772 46889 583800 190426
rect 583864 89554 583892 192918
rect 583852 89548 583904 89554
rect 583852 89490 583904 89496
rect 583758 46880 583814 46889
rect 583758 46815 583814 46824
rect 580262 6624 580318 6633
rect 580262 6559 580318 6568
rect 579774 354 579886 480
rect 579632 326 579886 354
rect 579774 -960 579886 326
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3422 566888 3478 566944
rect 3422 553832 3478 553888
rect 3422 527856 3478 527912
rect 3422 514820 3478 514856
rect 3422 514800 3424 514820
rect 3424 514800 3476 514820
rect 3476 514800 3478 514820
rect 3054 501744 3110 501800
rect 3422 475632 3478 475688
rect 3238 462576 3294 462632
rect 3146 449520 3202 449576
rect 3422 423544 3478 423600
rect 3146 410488 3202 410544
rect 3422 397468 3424 397488
rect 3424 397468 3476 397488
rect 3476 397468 3478 397488
rect 3422 397432 3478 397468
rect 3422 371320 3478 371376
rect 3422 358400 3478 358456
rect 3514 345344 3570 345400
rect 3422 319232 3478 319288
rect 3238 306176 3294 306232
rect 3422 293120 3478 293176
rect 3054 267144 3110 267200
rect 2778 254108 2834 254144
rect 2778 254088 2780 254108
rect 2780 254088 2832 254108
rect 2832 254088 2834 254108
rect 3422 241032 3478 241088
rect 3330 214920 3386 214976
rect 3422 201864 3478 201920
rect 3422 188808 3478 188864
rect 3698 162832 3754 162888
rect 3422 149776 3478 149832
rect 3238 136720 3294 136776
rect 2778 110608 2834 110664
rect 3422 97588 3424 97608
rect 3424 97588 3476 97608
rect 3476 97588 3478 97608
rect 3422 97552 3478 97588
rect 3146 84632 3202 84688
rect 3422 71576 3478 71632
rect 2778 64096 2834 64152
rect 3054 58520 3110 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3514 32408 3570 32464
rect 3422 19352 3478 19408
rect 8298 40568 8354 40624
rect 3422 6432 3478 6488
rect 11058 46144 11114 46200
rect 17958 75112 18014 75168
rect 13818 66816 13874 66872
rect 35162 239400 35218 239456
rect 35806 239400 35862 239456
rect 32402 4800 32458 4856
rect 46202 242936 46258 242992
rect 41326 182960 41382 183016
rect 54942 203496 54998 203552
rect 50986 187040 51042 187096
rect 57610 239808 57666 239864
rect 59174 263628 59230 263664
rect 59174 263608 59176 263628
rect 59176 263608 59228 263628
rect 59228 263608 59230 263628
rect 59266 195200 59322 195256
rect 59174 188264 59230 188320
rect 61842 240080 61898 240136
rect 64602 298152 64658 298208
rect 61934 218592 61990 218648
rect 66902 292984 66958 293040
rect 66902 286320 66958 286376
rect 67638 290400 67694 290456
rect 67730 289720 67786 289776
rect 67638 289040 67694 289096
rect 67638 287680 67694 287736
rect 67730 287000 67786 287056
rect 67638 285676 67640 285696
rect 67640 285676 67692 285696
rect 67692 285676 67694 285696
rect 67638 285640 67694 285676
rect 68742 291080 68798 291136
rect 68834 288360 68890 288416
rect 68558 284960 68614 285016
rect 67638 284316 67640 284336
rect 67640 284316 67692 284336
rect 67692 284316 67694 284336
rect 67638 284280 67694 284316
rect 67730 283600 67786 283656
rect 67822 282920 67878 282976
rect 67638 281560 67694 281616
rect 68282 280880 68338 280936
rect 67638 280220 67694 280256
rect 67638 280200 67640 280220
rect 67640 280200 67692 280220
rect 67692 280200 67694 280220
rect 67638 279520 67694 279576
rect 67546 278840 67602 278896
rect 68098 278160 68154 278216
rect 67638 277480 67694 277536
rect 67730 276800 67786 276856
rect 67638 276120 67694 276176
rect 67638 275440 67694 275496
rect 67454 274760 67510 274816
rect 67362 269320 67418 269376
rect 64786 181464 64842 181520
rect 67270 251640 67326 251696
rect 66074 129240 66130 129296
rect 66166 126248 66222 126304
rect 66166 125160 66222 125216
rect 64786 124208 64842 124264
rect 66166 124208 66222 124264
rect 60646 94832 60702 94888
rect 57886 89664 57942 89720
rect 64694 102176 64750 102232
rect 66074 123528 66130 123584
rect 66166 122576 66222 122632
rect 55126 85448 55182 85504
rect 67730 274080 67786 274136
rect 67638 273400 67694 273456
rect 67638 272720 67694 272776
rect 67638 271360 67694 271416
rect 67730 270680 67786 270736
rect 67638 270000 67694 270056
rect 68190 268640 68246 268696
rect 67638 267960 67694 268016
rect 67638 266600 67694 266656
rect 67730 265920 67786 265976
rect 67638 265240 67694 265296
rect 67638 264560 67694 264616
rect 67638 263880 67694 263936
rect 67730 263200 67786 263256
rect 67638 262520 67694 262576
rect 67730 261840 67786 261896
rect 68190 261160 68246 261216
rect 67638 260480 67694 260536
rect 67638 259800 67694 259856
rect 67730 259120 67786 259176
rect 67638 258440 67694 258496
rect 67638 257760 67694 257816
rect 67638 257080 67694 257136
rect 67638 255720 67694 255776
rect 67730 254360 67786 254416
rect 67638 253680 67694 253736
rect 68374 272040 68430 272096
rect 70674 292576 70730 292632
rect 71686 292304 71742 292360
rect 73894 294480 73950 294536
rect 77758 292712 77814 292768
rect 94594 296928 94650 296984
rect 95146 295976 95202 296032
rect 95790 294072 95846 294128
rect 97722 298288 97778 298344
rect 98734 294480 98790 294536
rect 103518 294208 103574 294264
rect 106738 293936 106794 293992
rect 108026 292848 108082 292904
rect 111246 295296 111302 295352
rect 114190 291896 114246 291952
rect 117226 294072 117282 294128
rect 117686 294072 117742 294128
rect 68926 267280 68982 267336
rect 69202 256400 69258 256456
rect 69018 253000 69074 253056
rect 68926 252320 68982 252376
rect 67730 250960 67786 251016
rect 67638 250280 67694 250336
rect 67638 249600 67694 249656
rect 67638 248920 67694 248976
rect 67730 248240 67786 248296
rect 67638 247560 67694 247616
rect 68098 245556 68100 245576
rect 68100 245556 68152 245576
rect 68152 245556 68154 245576
rect 68098 245520 68154 245556
rect 68006 244840 68062 244896
rect 67546 244160 67602 244216
rect 67638 242120 67694 242176
rect 67454 188400 67510 188456
rect 69294 245520 69350 245576
rect 73158 186904 73214 186960
rect 75826 230424 75882 230480
rect 98366 238176 98422 238232
rect 74538 181328 74594 181384
rect 98642 178608 98698 178664
rect 102046 177656 102102 177712
rect 106738 238312 106794 238368
rect 115110 238448 115166 238504
rect 117042 239672 117098 239728
rect 118974 238584 119030 238640
rect 117226 237088 117282 237144
rect 120906 294208 120962 294264
rect 120814 292712 120870 292768
rect 120814 282240 120870 282296
rect 120722 268640 120778 268696
rect 120170 250960 120226 251016
rect 120722 250996 120724 251016
rect 120724 250996 120776 251016
rect 120776 250996 120778 251016
rect 120722 250960 120778 250996
rect 120078 241440 120134 241496
rect 121458 291760 121514 291816
rect 121458 291080 121514 291136
rect 121550 290400 121606 290456
rect 121458 289756 121460 289776
rect 121460 289756 121512 289776
rect 121512 289756 121514 289776
rect 121458 289720 121514 289756
rect 122010 289040 122066 289096
rect 121550 288360 121606 288416
rect 121458 287680 121514 287736
rect 121642 287000 121698 287056
rect 121458 286320 121514 286376
rect 121550 284960 121606 285016
rect 121458 284280 121514 284336
rect 121458 282940 121514 282976
rect 121458 282920 121460 282940
rect 121460 282920 121512 282940
rect 121512 282920 121514 282940
rect 121458 281580 121514 281616
rect 121458 281560 121460 281580
rect 121460 281560 121512 281580
rect 121512 281560 121514 281580
rect 121458 280220 121514 280256
rect 121458 280200 121460 280220
rect 121460 280200 121512 280220
rect 121512 280200 121514 280220
rect 121550 279520 121606 279576
rect 121458 278860 121514 278896
rect 121458 278840 121460 278860
rect 121460 278840 121512 278860
rect 121512 278840 121514 278860
rect 121550 278160 121606 278216
rect 121458 277480 121514 277536
rect 122102 285640 122158 285696
rect 122378 280880 122434 280936
rect 121550 276800 121606 276856
rect 121458 276120 121514 276176
rect 121550 275440 121606 275496
rect 121458 274780 121514 274816
rect 121458 274760 121460 274780
rect 121460 274760 121512 274780
rect 121512 274760 121514 274780
rect 121458 274080 121514 274136
rect 121458 273400 121514 273456
rect 121458 272060 121514 272096
rect 121458 272040 121460 272060
rect 121460 272040 121512 272060
rect 121512 272040 121514 272060
rect 121458 271360 121514 271416
rect 121550 270000 121606 270056
rect 121458 269320 121514 269376
rect 122102 267280 122158 267336
rect 121458 266600 121514 266656
rect 121458 265920 121514 265976
rect 121550 264560 121606 264616
rect 121458 263880 121514 263936
rect 121458 263200 121514 263256
rect 121458 262520 121514 262576
rect 121550 261840 121606 261896
rect 121458 261160 121514 261216
rect 121550 260480 121606 260536
rect 121458 259800 121514 259856
rect 121550 259120 121606 259176
rect 121458 258440 121514 258496
rect 121550 257760 121606 257816
rect 121458 257080 121514 257136
rect 121550 256400 121606 256456
rect 121458 255720 121514 255776
rect 121458 254360 121514 254416
rect 121550 253680 121606 253736
rect 121458 253000 121514 253056
rect 121550 252320 121606 252376
rect 121458 251640 121514 251696
rect 121458 250280 121514 250336
rect 121458 248920 121514 248976
rect 121458 248240 121514 248296
rect 121550 246880 121606 246936
rect 121458 246200 121514 246256
rect 121550 245520 121606 245576
rect 121458 244840 121514 244896
rect 121550 244160 121606 244216
rect 121458 243480 121514 243536
rect 121458 242800 121514 242856
rect 121642 242120 121698 242176
rect 121458 240760 121514 240816
rect 121550 240080 121606 240136
rect 122286 272720 122342 272776
rect 122102 232464 122158 232520
rect 100666 177520 100722 177576
rect 103426 177520 103482 177576
rect 110418 179424 110474 179480
rect 110234 176976 110290 177032
rect 104622 176704 104678 176760
rect 107014 176740 107016 176760
rect 107016 176740 107068 176760
rect 107068 176740 107070 176760
rect 107014 176704 107070 176740
rect 108118 176704 108174 176760
rect 110694 177520 110750 177576
rect 112994 177520 113050 177576
rect 115846 177520 115902 177576
rect 114374 176976 114430 177032
rect 119986 177520 120042 177576
rect 121090 177520 121146 177576
rect 123574 240760 123630 240816
rect 124126 242528 124182 242584
rect 123482 182824 123538 182880
rect 127622 295296 127678 295352
rect 125046 181600 125102 181656
rect 129646 295976 129702 296032
rect 130474 357448 130530 357504
rect 131762 204856 131818 204912
rect 133142 190984 133198 191040
rect 145654 291896 145710 291952
rect 145654 227568 145710 227624
rect 127622 184184 127678 184240
rect 126886 177520 126942 177576
rect 128082 177520 128138 177576
rect 130750 177520 130806 177576
rect 147218 226208 147274 226264
rect 152462 365744 152518 365800
rect 149702 299376 149758 299432
rect 156510 257216 156566 257272
rect 158442 296792 158498 296848
rect 157338 254224 157394 254280
rect 157246 237224 157302 237280
rect 132038 176976 132094 177032
rect 160558 311908 160614 311944
rect 160558 311888 160560 311908
rect 160560 311888 160612 311908
rect 160612 311888 160614 311908
rect 159454 231784 159510 231840
rect 160098 244840 160154 244896
rect 161294 244840 161350 244896
rect 161294 213832 161350 213888
rect 157982 177248 158038 177304
rect 118422 176704 118478 176760
rect 122746 176704 122802 176760
rect 123022 176704 123078 176760
rect 128174 176704 128230 176760
rect 129462 176704 129518 176760
rect 133142 176704 133198 176760
rect 135718 176704 135774 176760
rect 148230 176704 148286 176760
rect 158994 176724 159050 176760
rect 158994 176704 158996 176724
rect 158996 176704 159048 176724
rect 159048 176704 159050 176724
rect 162306 229744 162362 229800
rect 164146 179968 164202 180024
rect 165618 266348 165674 266384
rect 165618 266328 165620 266348
rect 165620 266328 165672 266348
rect 165672 266328 165674 266348
rect 165066 241168 165122 241224
rect 164974 189624 165030 189680
rect 116950 175616 117006 175672
rect 124494 175616 124550 175672
rect 134430 175616 134486 175672
rect 98366 175344 98422 175400
rect 67638 128016 67694 128072
rect 67454 120808 67510 120864
rect 67730 100680 67786 100736
rect 67454 90888 67510 90944
rect 166262 178744 166318 178800
rect 169758 297336 169814 297392
rect 170494 293936 170550 293992
rect 168378 242120 168434 242176
rect 167734 184320 167790 184376
rect 166998 176840 167054 176896
rect 167642 171536 167698 171592
rect 172334 160112 172390 160168
rect 112350 94696 112406 94752
rect 113178 94696 113234 94752
rect 123206 94696 123262 94752
rect 151910 94696 151966 94752
rect 125598 94424 125654 94480
rect 121734 93608 121790 93664
rect 93950 93472 94006 93528
rect 107750 93472 107806 93528
rect 110142 93200 110198 93256
rect 85762 92384 85818 92440
rect 87234 92384 87290 92440
rect 88982 92420 88984 92440
rect 88984 92420 89036 92440
rect 89036 92420 89038 92440
rect 88982 92384 89038 92420
rect 100482 92384 100538 92440
rect 107474 92384 107530 92440
rect 109682 92384 109738 92440
rect 75826 91160 75882 91216
rect 85486 91160 85542 91216
rect 99286 91432 99342 91488
rect 99102 91296 99158 91352
rect 86866 91160 86922 91216
rect 90730 91160 90786 91216
rect 92386 91160 92442 91216
rect 93766 91160 93822 91216
rect 95146 91160 95202 91216
rect 96526 91160 96582 91216
rect 97078 91160 97134 91216
rect 97906 91160 97962 91216
rect 97078 86808 97134 86864
rect 99194 91160 99250 91216
rect 104254 91568 104310 91624
rect 101862 91432 101918 91488
rect 100574 91160 100630 91216
rect 102046 91296 102102 91352
rect 103334 91296 103390 91352
rect 101954 91160 102010 91216
rect 101954 82728 102010 82784
rect 103426 91160 103482 91216
rect 106186 91296 106242 91352
rect 104806 91160 104862 91216
rect 106094 91160 106150 91216
rect 103426 81368 103482 81424
rect 106094 84088 106150 84144
rect 107566 91160 107622 91216
rect 108486 91160 108542 91216
rect 111614 92384 111670 92440
rect 114190 92384 114246 92440
rect 118054 92404 118110 92440
rect 118054 92384 118056 92404
rect 118056 92384 118108 92404
rect 118108 92384 118110 92404
rect 110234 91160 110290 91216
rect 124494 92384 124550 92440
rect 125414 92384 125470 92440
rect 115386 91704 115442 91760
rect 111706 91160 111762 91216
rect 113086 91160 113142 91216
rect 113914 91160 113970 91216
rect 110234 88168 110290 88224
rect 124126 91432 124182 91488
rect 119894 91296 119950 91352
rect 120722 91296 120778 91352
rect 115846 91160 115902 91216
rect 117134 91160 117190 91216
rect 118238 91160 118294 91216
rect 119986 91160 120042 91216
rect 121366 91160 121422 91216
rect 122746 91160 122802 91216
rect 124034 91160 124090 91216
rect 55218 36488 55274 36544
rect 67638 59880 67694 59936
rect 69018 54440 69074 54496
rect 77390 17176 77446 17232
rect 117318 26832 117374 26888
rect 125782 92384 125838 92440
rect 151542 93472 151598 93528
rect 128174 93200 128230 93256
rect 126886 91296 126942 91352
rect 126794 91160 126850 91216
rect 128358 93064 128414 93120
rect 129462 92384 129518 92440
rect 135718 92384 135774 92440
rect 151726 92112 151782 92168
rect 132222 91568 132278 91624
rect 151358 91568 151414 91624
rect 130750 91160 130806 91216
rect 133142 91160 133198 91216
rect 134706 91160 134762 91216
rect 167918 111696 167974 111752
rect 167826 110064 167882 110120
rect 168102 108704 168158 108760
rect 173162 95104 173218 95160
rect 176658 354320 176714 354376
rect 176566 352144 176622 352200
rect 176474 309984 176530 310040
rect 176382 292304 176438 292360
rect 176474 252864 176530 252920
rect 176658 345344 176714 345400
rect 176842 343304 176898 343360
rect 176842 334464 176898 334520
rect 176658 332560 176714 332616
rect 176658 327664 176714 327720
rect 176658 325760 176714 325816
rect 177946 321544 178002 321600
rect 177854 318824 177910 318880
rect 176658 314744 176714 314800
rect 176658 312704 176714 312760
rect 176658 305904 176714 305960
rect 176658 301144 176714 301200
rect 176658 299104 176714 299160
rect 176658 297200 176714 297256
rect 176658 295024 176714 295080
rect 176658 290264 176714 290320
rect 176658 286184 176714 286240
rect 176658 283464 176714 283520
rect 176658 281580 176714 281616
rect 176658 281560 176660 281580
rect 176660 281560 176712 281580
rect 176712 281560 176714 281580
rect 176658 279520 176714 279576
rect 176658 277480 176714 277536
rect 177486 274760 177542 274816
rect 176658 272584 176714 272640
rect 177762 270544 177818 270600
rect 176658 268504 176714 268560
rect 176658 265920 176714 265976
rect 176658 261704 176714 261760
rect 176658 259664 176714 259720
rect 176658 254904 176714 254960
rect 177670 250824 177726 250880
rect 176658 246064 176714 246120
rect 177578 241984 177634 242040
rect 178682 288360 178738 288416
rect 179786 357720 179842 357776
rect 193218 357584 193274 357640
rect 193862 357584 193918 357640
rect 201498 355272 201554 355328
rect 206282 357448 206338 357504
rect 213918 364384 213974 364440
rect 211802 357720 211858 357776
rect 209962 354864 210018 354920
rect 243634 363024 243690 363080
rect 242162 357448 242218 357504
rect 258906 358808 258962 358864
rect 269026 357720 269082 357776
rect 256790 354864 256846 354920
rect 274546 356088 274602 356144
rect 247038 354728 247094 354784
rect 248142 354728 248198 354784
rect 282090 356224 282146 356280
rect 291750 354592 291806 354648
rect 292210 354592 292266 354648
rect 179510 348132 179566 348188
rect 179510 341332 179566 341388
rect 179142 336504 179198 336560
rect 179050 257080 179106 257136
rect 179050 246064 179106 246120
rect 179050 224576 179106 224632
rect 293130 338680 293186 338736
rect 293866 338680 293922 338736
rect 293958 334600 294014 334656
rect 295338 349560 295394 349616
rect 296166 357584 296222 357640
rect 296074 354320 296130 354376
rect 295982 345480 296038 345536
rect 295338 340720 295394 340776
rect 295338 336676 295340 336696
rect 295340 336676 295392 336696
rect 295392 336676 295394 336696
rect 295338 336640 295394 336676
rect 295338 331900 295394 331936
rect 295338 331880 295340 331900
rect 295340 331880 295392 331900
rect 295392 331880 295394 331900
rect 294050 329840 294106 329896
rect 294326 329860 294382 329896
rect 294326 329840 294328 329860
rect 294328 329840 294380 329860
rect 294380 329840 294382 329860
rect 293038 328344 293094 328400
rect 294142 325760 294198 325816
rect 179510 308012 179566 308068
rect 179234 303864 179290 303920
rect 179326 263744 179382 263800
rect 179418 248104 179474 248160
rect 293222 301280 293278 301336
rect 293130 287680 293186 287736
rect 293038 268096 293094 268152
rect 179786 244092 179842 244148
rect 179510 242936 179566 242992
rect 204258 240624 204314 240680
rect 180890 234368 180946 234424
rect 186962 187176 187018 187232
rect 192206 237088 192262 237144
rect 191194 94832 191250 94888
rect 192482 84768 192538 84824
rect 194046 89664 194102 89720
rect 198002 191120 198058 191176
rect 276294 240624 276350 240680
rect 207386 237360 207442 237416
rect 202142 235184 202198 235240
rect 206282 232600 206338 232656
rect 206374 171672 206430 171728
rect 211802 179968 211858 180024
rect 215206 239400 215262 239456
rect 213918 175616 213974 175672
rect 213918 174936 213974 174992
rect 214010 174256 214066 174312
rect 213918 173576 213974 173632
rect 214010 172896 214066 172952
rect 214194 172216 214250 172272
rect 214102 171536 214158 171592
rect 213918 170312 213974 170368
rect 213918 169668 213920 169688
rect 213920 169668 213972 169688
rect 213972 169668 213974 169688
rect 213918 169632 213974 169668
rect 214010 168952 214066 169008
rect 214010 168292 214066 168328
rect 214010 168272 214012 168292
rect 214012 168272 214064 168292
rect 214064 168272 214066 168292
rect 213918 167592 213974 167648
rect 213918 166912 213974 166968
rect 214102 166368 214158 166424
rect 214010 165688 214066 165744
rect 213918 165008 213974 165064
rect 214010 163648 214066 163704
rect 213918 162968 213974 163024
rect 214562 162288 214618 162344
rect 213918 161744 213974 161800
rect 214746 170992 214802 171048
rect 213918 161064 213974 161120
rect 214010 160384 214066 160440
rect 213918 159024 213974 159080
rect 213918 158344 213974 158400
rect 214930 157664 214986 157720
rect 213918 157120 213974 157176
rect 214010 156440 214066 156496
rect 213918 155760 213974 155816
rect 214010 154400 214066 154456
rect 213918 153720 213974 153776
rect 213918 153040 213974 153096
rect 214010 152496 214066 152552
rect 214654 151816 214710 151872
rect 214010 151136 214066 151192
rect 213918 150476 213974 150512
rect 213918 150456 213920 150476
rect 213920 150456 213972 150476
rect 213972 150456 213974 150476
rect 214010 149776 214066 149832
rect 213918 149096 213974 149152
rect 213918 148416 213974 148472
rect 214102 147872 214158 147928
rect 214010 147192 214066 147248
rect 213918 146512 213974 146568
rect 214010 145832 214066 145888
rect 213918 145152 213974 145208
rect 213918 144472 213974 144528
rect 214654 143792 214710 143848
rect 213918 143248 213974 143304
rect 214562 142568 214618 142624
rect 214010 141888 214066 141944
rect 213918 141208 213974 141264
rect 213918 140528 213974 140584
rect 214010 139168 214066 139224
rect 213918 138624 213974 138680
rect 214010 135904 214066 135960
rect 213918 135224 213974 135280
rect 213918 134544 213974 134600
rect 213918 133320 213974 133376
rect 213918 131280 213974 131336
rect 214010 129240 214066 129296
rect 213918 128696 213974 128752
rect 213918 128016 213974 128072
rect 214010 126656 214066 126712
rect 213918 125976 213974 126032
rect 214010 125296 214066 125352
rect 213918 124616 213974 124672
rect 214010 124072 214066 124128
rect 213918 123392 213974 123448
rect 214010 122712 214066 122768
rect 213918 122032 213974 122088
rect 214010 121352 214066 121408
rect 213918 120672 213974 120728
rect 214102 119992 214158 120048
rect 214010 119448 214066 119504
rect 213918 118768 213974 118824
rect 214010 118088 214066 118144
rect 213918 117428 213974 117464
rect 213918 117408 213920 117428
rect 213920 117408 213972 117428
rect 213972 117408 213974 117428
rect 213182 116728 213238 116784
rect 213918 116048 213974 116104
rect 214010 115368 214066 115424
rect 213918 114824 213974 114880
rect 214010 114144 214066 114200
rect 213918 113464 213974 113520
rect 214010 112784 214066 112840
rect 213918 112104 213974 112160
rect 214010 111424 214066 111480
rect 213918 110744 213974 110800
rect 214010 110200 214066 110256
rect 213918 109520 213974 109576
rect 214010 108840 214066 108896
rect 213918 108160 213974 108216
rect 214010 107480 214066 107536
rect 213918 106800 213974 106856
rect 214010 106120 214066 106176
rect 214102 105576 214158 105632
rect 213918 104896 213974 104952
rect 214010 104216 214066 104272
rect 213918 103572 213920 103592
rect 213920 103572 213972 103592
rect 213972 103572 213974 103592
rect 213918 103536 213974 103572
rect 214654 139848 214710 139904
rect 214654 137264 214710 137320
rect 214746 136584 214802 136640
rect 214010 102856 214066 102912
rect 213918 102196 213974 102232
rect 213918 102176 213920 102196
rect 213920 102176 213972 102196
rect 213972 102176 213974 102196
rect 213918 100952 213974 101008
rect 214010 100272 214066 100328
rect 213918 98912 213974 98968
rect 213918 97552 213974 97608
rect 213918 96328 213974 96384
rect 214102 99592 214158 99648
rect 214562 98232 214618 98288
rect 214930 97144 214986 97200
rect 214838 96872 214894 96928
rect 229098 189760 229154 189816
rect 236274 238448 236330 238504
rect 233882 238176 233938 238232
rect 229742 182960 229798 183016
rect 233882 177520 233938 177576
rect 240506 238584 240562 238640
rect 238022 181600 238078 181656
rect 232502 175888 232558 175944
rect 244278 177384 244334 177440
rect 246394 179152 246450 179208
rect 254674 238448 254730 238504
rect 247682 176024 247738 176080
rect 248050 175752 248106 175808
rect 249154 175208 249210 175264
rect 249338 173304 249394 173360
rect 249430 172760 249486 172816
rect 249246 171808 249302 171864
rect 249154 160520 249210 160576
rect 249798 153448 249854 153504
rect 250166 164328 250222 164384
rect 251178 157800 251234 157856
rect 251178 156304 251234 156360
rect 249890 151136 249946 151192
rect 251178 149776 251234 149832
rect 251822 172352 251878 172408
rect 252558 171400 252614 171456
rect 251730 170856 251786 170912
rect 251822 170448 251878 170504
rect 252466 169088 252522 169144
rect 252466 168172 252468 168192
rect 252468 168172 252520 168192
rect 252520 168172 252522 168192
rect 252466 168136 252522 168172
rect 252466 167592 252522 167648
rect 252374 167184 252430 167240
rect 252374 166640 252430 166696
rect 252466 166232 252522 166288
rect 252282 165688 252338 165744
rect 252466 165280 252522 165336
rect 252466 164736 252522 164792
rect 252190 162968 252246 163024
rect 252098 162424 252154 162480
rect 252466 162016 252522 162072
rect 251546 161472 251602 161528
rect 251546 160112 251602 160168
rect 251454 159160 251510 159216
rect 251362 158752 251418 158808
rect 252466 158208 252522 158264
rect 251914 157936 251970 157992
rect 251362 156848 251418 156904
rect 251822 154944 251878 155000
rect 252374 155896 252430 155952
rect 252466 155352 252522 155408
rect 252742 169496 252798 169552
rect 253202 163920 253258 163976
rect 253202 162968 253258 163024
rect 252650 154400 252706 154456
rect 252466 153992 252522 154048
rect 252466 153076 252468 153096
rect 252468 153076 252520 153096
rect 252520 153076 252522 153096
rect 252466 153040 252522 153076
rect 252374 152632 252430 152688
rect 252282 152088 252338 152144
rect 251270 149232 251326 149288
rect 251914 150728 251970 150784
rect 251822 148824 251878 148880
rect 251730 146920 251786 146976
rect 251546 144608 251602 144664
rect 251914 144064 251970 144120
rect 250626 143112 250682 143168
rect 251086 142568 251142 142624
rect 218058 95920 218114 95976
rect 242898 3168 242954 3224
rect 249246 97008 249302 97064
rect 250994 95648 251050 95704
rect 251730 139848 251786 139904
rect 251730 139440 251786 139496
rect 251362 138488 251418 138544
rect 251730 135632 251786 135688
rect 251730 132776 251786 132832
rect 251730 129104 251786 129160
rect 251178 125332 251180 125352
rect 251180 125332 251232 125352
rect 251232 125332 251234 125352
rect 251178 125296 251234 125332
rect 251546 120536 251602 120592
rect 251546 114008 251602 114064
rect 251546 112104 251602 112160
rect 251546 106936 251602 106992
rect 251638 105984 251694 106040
rect 251270 104080 251326 104136
rect 251178 98948 251180 98968
rect 251180 98948 251232 98968
rect 251232 98948 251234 98968
rect 251178 98912 251234 98948
rect 251178 96600 251234 96656
rect 252466 151716 252468 151736
rect 252468 151716 252520 151736
rect 252520 151716 252522 151736
rect 252466 151680 252522 151716
rect 253202 149640 253258 149696
rect 252466 148280 252522 148336
rect 252466 147500 252468 147520
rect 252468 147500 252520 147520
rect 252520 147500 252522 147520
rect 252466 147464 252522 147500
rect 252374 146512 252430 146568
rect 252098 145968 252154 146024
rect 252282 145016 252338 145072
rect 252466 143656 252522 143712
rect 252466 142704 252522 142760
rect 252374 142160 252430 142216
rect 252466 141344 252522 141400
rect 252098 140392 252154 140448
rect 252098 137536 252154 137592
rect 251914 131416 251970 131472
rect 252098 136176 252154 136232
rect 252466 136992 252522 137048
rect 252374 135224 252430 135280
rect 252466 134680 252522 134736
rect 252282 134272 252338 134328
rect 252466 133748 252522 133784
rect 252466 133728 252468 133748
rect 252468 133728 252520 133748
rect 252520 133728 252522 133748
rect 252374 133320 252430 133376
rect 252466 132404 252468 132424
rect 252468 132404 252520 132424
rect 252520 132404 252522 132424
rect 252466 132368 252522 132404
rect 252466 131824 252522 131880
rect 252466 130872 252522 130928
rect 252374 130464 252430 130520
rect 252190 130056 252246 130112
rect 252466 129512 252522 129568
rect 252374 128560 252430 128616
rect 252466 128152 252522 128208
rect 252374 127200 252430 127256
rect 251822 117816 251878 117872
rect 252466 126656 252522 126712
rect 252466 126248 252522 126304
rect 252374 125704 252430 125760
rect 252466 124752 252522 124808
rect 252374 124344 252430 124400
rect 252466 123936 252522 123992
rect 252374 123392 252430 123448
rect 252282 122984 252338 123040
rect 252466 122440 252522 122496
rect 252374 122032 252430 122088
rect 252466 121488 252522 121544
rect 252466 121080 252522 121136
rect 252374 120128 252430 120184
rect 252098 119176 252154 119232
rect 252466 119584 252522 119640
rect 252374 118768 252430 118824
rect 252006 116356 252008 116376
rect 252008 116356 252060 116376
rect 252060 116356 252062 116376
rect 252006 116320 252062 116356
rect 251914 115912 251970 115968
rect 252006 114960 252062 115016
rect 251822 113464 251878 113520
rect 252466 118224 252522 118280
rect 252374 117272 252430 117328
rect 252466 116864 252522 116920
rect 252282 115368 252338 115424
rect 252466 114436 252522 114472
rect 252466 114416 252468 114436
rect 252468 114416 252520 114436
rect 252520 114416 252522 114436
rect 252098 109792 252154 109848
rect 252098 107888 252154 107944
rect 251822 104624 251878 104680
rect 251914 102720 251970 102776
rect 251822 101360 251878 101416
rect 252098 105032 252154 105088
rect 252098 103672 252154 103728
rect 252374 113056 252430 113112
rect 252466 112648 252522 112704
rect 252374 111716 252430 111752
rect 252374 111696 252376 111716
rect 252376 111696 252428 111716
rect 252428 111696 252430 111716
rect 252466 110744 252522 110800
rect 252466 110200 252522 110256
rect 252374 109248 252430 109304
rect 252466 108840 252522 108896
rect 252374 108296 252430 108352
rect 252466 107480 252522 107536
rect 252374 106528 252430 106584
rect 252466 105576 252522 105632
rect 252282 104216 252338 104272
rect 252190 103128 252246 103184
rect 252466 102176 252522 102232
rect 252374 101768 252430 101824
rect 252466 101360 252522 101416
rect 252098 100816 252154 100872
rect 252006 100408 252062 100464
rect 251914 99864 251970 99920
rect 252098 99456 252154 99512
rect 251822 97824 251878 97880
rect 252374 98504 252430 98560
rect 252282 97960 252338 98016
rect 251914 97552 251970 97608
rect 251822 97008 251878 97064
rect 254214 177248 254270 177304
rect 255318 176432 255374 176488
rect 254122 146240 254178 146296
rect 252466 96600 252522 96656
rect 256238 146240 256294 146296
rect 259458 6296 259514 6352
rect 255870 3440 255926 3496
rect 257066 3440 257122 3496
rect 265622 228928 265678 228984
rect 265622 227704 265678 227760
rect 262954 148144 263010 148200
rect 271234 3440 271290 3496
rect 278318 3304 278374 3360
rect 283930 134408 283986 134464
rect 287702 238856 287758 238912
rect 287886 238720 287942 238776
rect 287058 26968 287114 27024
rect 285770 26832 285826 26888
rect 287978 145560 288034 145616
rect 291106 238720 291162 238776
rect 293958 299240 294014 299296
rect 293314 241440 293370 241496
rect 294050 263880 294106 263936
rect 294234 323040 294290 323096
rect 295338 321000 295394 321056
rect 295338 318960 295394 319016
rect 295338 316920 295394 316976
rect 295338 314200 295394 314256
rect 295338 311908 295394 311944
rect 295338 311888 295340 311908
rect 295340 311888 295392 311908
rect 295392 311888 295394 311908
rect 295338 310120 295394 310176
rect 295338 308080 295394 308136
rect 295338 305360 295394 305416
rect 295338 303320 295394 303376
rect 295338 296520 295394 296576
rect 295338 294480 295394 294536
rect 296626 292440 296682 292496
rect 296074 290400 296130 290456
rect 295338 285676 295340 285696
rect 295340 285676 295392 285696
rect 295392 285676 295394 285696
rect 295338 285640 295394 285676
rect 295338 283600 295394 283656
rect 295338 281580 295394 281616
rect 295338 281560 295340 281580
rect 295340 281560 295392 281580
rect 295392 281560 295394 281580
rect 295338 278860 295394 278896
rect 295338 278840 295340 278860
rect 295340 278840 295392 278860
rect 295392 278840 295394 278860
rect 295338 276800 295394 276856
rect 295338 274760 295394 274816
rect 295338 272720 295394 272776
rect 295338 270000 295394 270056
rect 295338 265920 295394 265976
rect 295338 261180 295394 261216
rect 295338 261160 295340 261180
rect 295340 261160 295392 261180
rect 295392 261160 295394 261180
rect 295338 259120 295394 259176
rect 295982 257080 296038 257136
rect 295614 255040 295670 255096
rect 295522 248240 295578 248296
rect 295522 246200 295578 246256
rect 295798 243480 295854 243536
rect 296534 252048 296590 252104
rect 297178 252048 297234 252104
rect 296626 250280 296682 250336
rect 296534 248376 296590 248432
rect 296074 3304 296130 3360
rect 299478 240760 299534 240816
rect 297730 139984 297786 140040
rect 305734 510584 305790 510640
rect 300950 231784 301006 231840
rect 301042 224712 301098 224768
rect 300858 128968 300914 129024
rect 303618 193840 303674 193896
rect 306470 233144 306526 233200
rect 306378 175888 306434 175944
rect 306746 174800 306802 174856
rect 307666 174392 307722 174448
rect 307298 174020 307300 174040
rect 307300 174020 307352 174040
rect 307352 174020 307354 174040
rect 307298 173984 307354 174020
rect 307574 173576 307630 173632
rect 307298 173168 307354 173224
rect 307666 172624 307722 172680
rect 306930 172216 306986 172272
rect 306562 171808 306618 171864
rect 307666 171400 307722 171456
rect 307390 170992 307446 171048
rect 306746 170584 306802 170640
rect 307298 169804 307300 169824
rect 307300 169804 307352 169824
rect 307352 169804 307354 169824
rect 307298 169768 307354 169804
rect 306746 169224 306802 169280
rect 307298 168428 307354 168464
rect 307298 168408 307300 168428
rect 307300 168408 307352 168428
rect 307352 168408 307354 168428
rect 307298 168000 307354 168056
rect 306562 166368 306618 166424
rect 307114 165008 307170 165064
rect 306746 162424 306802 162480
rect 306746 161200 306802 161256
rect 306746 156984 306802 157040
rect 306930 156168 306986 156224
rect 306562 153992 306618 154048
rect 307022 153584 307078 153640
rect 306562 152632 306618 152688
rect 306930 149232 306986 149288
rect 306562 145832 306618 145888
rect 305734 145424 305790 145480
rect 305642 124616 305698 124672
rect 306930 145052 306932 145072
rect 306932 145052 306984 145072
rect 306984 145052 306986 145072
rect 306930 145016 306986 145052
rect 306930 144608 306986 144664
rect 306562 144200 306618 144256
rect 306010 140800 306066 140856
rect 305826 106256 305882 106312
rect 305734 99456 305790 99512
rect 305918 103808 305974 103864
rect 306746 142432 306802 142488
rect 306930 139032 306986 139088
rect 306930 137808 306986 137864
rect 306930 136584 306986 136640
rect 306746 134816 306802 134872
rect 306930 133592 306986 133648
rect 306746 131008 306802 131064
rect 306746 125432 306802 125488
rect 307298 164192 307354 164248
rect 307206 162968 307262 163024
rect 307666 170176 307722 170232
rect 307574 168816 307630 168872
rect 307666 167592 307722 167648
rect 307482 167184 307538 167240
rect 307666 166776 307722 166832
rect 307482 165824 307538 165880
rect 307574 165416 307630 165472
rect 307666 164600 307722 164656
rect 307482 163784 307538 163840
rect 307666 163376 307722 163432
rect 307666 162016 307722 162072
rect 307482 161608 307538 161664
rect 307574 160792 307630 160848
rect 307666 160384 307722 160440
rect 307574 159976 307630 160032
rect 307482 159568 307538 159624
rect 307666 159024 307722 159080
rect 307666 158616 307722 158672
rect 307482 158208 307538 158264
rect 307574 157800 307630 157856
rect 307666 156576 307722 156632
rect 307666 155624 307722 155680
rect 307482 155216 307538 155272
rect 307298 154808 307354 154864
rect 307574 154400 307630 154456
rect 307666 153176 307722 153232
rect 307574 152224 307630 152280
rect 307666 151816 307722 151872
rect 307482 151408 307538 151464
rect 307574 151000 307630 151056
rect 307666 150612 307722 150648
rect 307666 150592 307668 150612
rect 307668 150592 307720 150612
rect 307720 150592 307722 150612
rect 307482 149776 307538 149832
rect 307574 148824 307630 148880
rect 307482 148416 307538 148472
rect 307666 148008 307722 148064
rect 307390 147600 307446 147656
rect 307482 147192 307538 147248
rect 307574 146784 307630 146840
rect 307666 146412 307668 146432
rect 307668 146412 307720 146432
rect 307720 146412 307722 146432
rect 307666 146376 307722 146412
rect 307666 143792 307722 143848
rect 307666 143384 307722 143440
rect 307482 142976 307538 143032
rect 307390 141616 307446 141672
rect 307206 138216 307262 138272
rect 307114 129820 307116 129840
rect 307116 129820 307168 129840
rect 307168 129820 307170 129840
rect 307114 129784 307170 129820
rect 307114 123004 307170 123040
rect 307114 122984 307116 123004
rect 307116 122984 307168 123004
rect 307168 122984 307170 123004
rect 306746 121216 306802 121272
rect 306562 119584 306618 119640
rect 307114 119040 307170 119096
rect 306930 118632 306986 118688
rect 306562 118224 306618 118280
rect 307022 115640 307078 115696
rect 306562 114008 306618 114064
rect 307114 114824 307170 114880
rect 306930 110200 306986 110256
rect 306746 103400 306802 103456
rect 306746 102040 306802 102096
rect 306562 99048 306618 99104
rect 307022 97824 307078 97880
rect 304354 6160 304410 6216
rect 307298 136992 307354 137048
rect 307666 141208 307722 141264
rect 307574 140392 307630 140448
rect 307666 139576 307722 139632
rect 307666 137400 307722 137456
rect 307482 136176 307538 136232
rect 307574 135632 307630 135688
rect 307666 135260 307668 135280
rect 307668 135260 307720 135280
rect 307720 135260 307722 135280
rect 307666 135224 307722 135260
rect 307666 134408 307722 134464
rect 307482 133184 307538 133240
rect 307482 132232 307538 132288
rect 307574 131824 307630 131880
rect 307666 131416 307722 131472
rect 307574 130600 307630 130656
rect 307666 130192 307722 130248
rect 307482 129240 307538 129296
rect 307666 128832 307722 128888
rect 307482 128016 307538 128072
rect 307666 127608 307722 127664
rect 307574 127200 307630 127256
rect 307574 126384 307630 126440
rect 307666 125840 307722 125896
rect 307482 125024 307538 125080
rect 307666 124244 307668 124264
rect 307668 124244 307720 124264
rect 307720 124244 307722 124264
rect 307666 124208 307722 124244
rect 307482 123800 307538 123856
rect 307666 123392 307722 123448
rect 307482 122440 307538 122496
rect 307574 122032 307630 122088
rect 307666 121644 307722 121680
rect 307666 121624 307668 121644
rect 307668 121624 307720 121644
rect 307720 121624 307722 121644
rect 307574 120808 307630 120864
rect 307666 120400 307722 120456
rect 307666 119992 307722 120048
rect 307666 117428 307722 117464
rect 307666 117408 307668 117428
rect 307668 117408 307720 117428
rect 307720 117408 307722 117428
rect 307574 117000 307630 117056
rect 307482 116592 307538 116648
rect 307666 116184 307722 116240
rect 307482 115232 307538 115288
rect 307574 114416 307630 114472
rect 307666 113192 307722 113248
rect 307574 112240 307630 112296
rect 307666 111852 307722 111888
rect 307666 111832 307668 111852
rect 307668 111832 307720 111852
rect 307720 111832 307722 111852
rect 307482 111424 307538 111480
rect 307666 111016 307722 111072
rect 307574 110608 307630 110664
rect 307666 109792 307722 109848
rect 307574 109248 307630 109304
rect 307390 108840 307446 108896
rect 307482 108432 307538 108488
rect 307666 108024 307722 108080
rect 307574 107616 307630 107672
rect 307482 107208 307538 107264
rect 307574 106800 307630 106856
rect 307666 106428 307668 106448
rect 307668 106428 307720 106448
rect 307720 106428 307722 106448
rect 307666 106392 307722 106428
rect 307482 106256 307538 106312
rect 307574 105440 307630 105496
rect 307666 105032 307722 105088
rect 307482 104624 307538 104680
rect 307666 104216 307722 104272
rect 307482 102992 307538 103048
rect 307666 102448 307722 102504
rect 307482 101632 307538 101688
rect 307574 101224 307630 101280
rect 307666 100836 307722 100872
rect 307666 100816 307668 100836
rect 307668 100816 307720 100836
rect 307720 100816 307722 100836
rect 307666 100408 307722 100464
rect 307482 100000 307538 100056
rect 307666 99456 307722 99512
rect 307574 98640 307630 98696
rect 307666 98232 307722 98288
rect 307482 97416 307538 97472
rect 307666 96600 307722 96656
rect 307666 96192 307722 96248
rect 310610 216552 310666 216608
rect 310610 215328 310666 215384
rect 313278 239808 313334 239864
rect 311254 215328 311310 215384
rect 310426 179968 310482 180024
rect 316038 352552 316094 352608
rect 313922 177248 313978 177304
rect 316038 178064 316094 178120
rect 317326 178064 317382 178120
rect 315486 175888 315542 175944
rect 324962 357720 325018 357776
rect 319442 195200 319498 195256
rect 320178 176704 320234 176760
rect 318154 176024 318210 176080
rect 321282 165688 321338 165744
rect 321834 148280 321890 148336
rect 322846 147736 322902 147792
rect 321742 139032 321798 139088
rect 322846 138488 322902 138544
rect 321650 122168 321706 122224
rect 321558 106800 321614 106856
rect 321742 106800 321798 106856
rect 321650 101088 321706 101144
rect 321558 96600 321614 96656
rect 321558 95104 321614 95160
rect 313278 50224 313334 50280
rect 324410 189080 324466 189136
rect 323674 185000 323730 185056
rect 324318 175480 324374 175536
rect 324318 173984 324374 174040
rect 324318 171672 324374 171728
rect 324318 170856 324374 170912
rect 324318 170040 324374 170096
rect 324318 169360 324374 169416
rect 324502 168544 324558 168600
rect 324870 172080 324926 172136
rect 324410 167728 324466 167784
rect 324318 167048 324374 167104
rect 324318 166232 324374 166288
rect 324318 165416 324374 165472
rect 323122 164736 323178 164792
rect 323398 164736 323454 164792
rect 324318 163920 324374 163976
rect 324410 163104 324466 163160
rect 324318 160792 324374 160848
rect 324318 159332 324320 159352
rect 324320 159332 324372 159352
rect 324372 159332 324374 159352
rect 324318 159296 324374 159332
rect 324318 158480 324374 158536
rect 324410 157800 324466 157856
rect 324318 156984 324374 157040
rect 324410 156304 324466 156360
rect 324318 154672 324374 154728
rect 324318 153992 324374 154048
rect 325054 174664 325110 174720
rect 325606 160112 325662 160168
rect 324410 153176 324466 153232
rect 324962 152360 325018 152416
rect 324410 151680 324466 151736
rect 324318 150864 324374 150920
rect 324318 150048 324374 150104
rect 324410 149368 324466 149424
rect 324318 147056 324374 147112
rect 324318 145424 324374 145480
rect 324318 144780 324320 144800
rect 324320 144780 324372 144800
rect 324372 144780 324374 144800
rect 324318 144744 324374 144780
rect 324410 143928 324466 143984
rect 324318 143112 324374 143168
rect 324410 142432 324466 142488
rect 324318 141616 324374 141672
rect 324410 140800 324466 140856
rect 324318 140120 324374 140176
rect 324318 137808 324374 137864
rect 324410 136992 324466 137048
rect 324318 136312 324374 136368
rect 324410 135496 324466 135552
rect 324318 134680 324374 134736
rect 324410 134000 324466 134056
rect 324318 133184 324374 133240
rect 324318 132404 324320 132424
rect 324320 132404 324372 132424
rect 324372 132404 324374 132424
rect 324318 132368 324374 132404
rect 324410 131688 324466 131744
rect 324318 130872 324374 130928
rect 324410 130056 324466 130112
rect 323030 129376 323086 129432
rect 325054 129376 325110 129432
rect 324318 128560 324374 128616
rect 324318 127744 324374 127800
rect 324502 127064 324558 127120
rect 324318 126248 324374 126304
rect 324318 125432 324374 125488
rect 324410 124752 324466 124808
rect 324318 123936 324374 123992
rect 324410 123120 324466 123176
rect 324318 122476 324320 122496
rect 324320 122476 324372 122496
rect 324372 122476 324374 122496
rect 324318 122440 324374 122476
rect 324318 120808 324374 120864
rect 324410 120128 324466 120184
rect 324318 119312 324374 119368
rect 324318 118532 324320 118552
rect 324320 118532 324372 118552
rect 324372 118532 324374 118552
rect 324318 118496 324374 118532
rect 324410 117816 324466 117872
rect 324318 117000 324374 117056
rect 324502 116320 324558 116376
rect 324318 115504 324374 115560
rect 324410 114688 324466 114744
rect 324318 114008 324374 114064
rect 324410 113192 324466 113248
rect 324318 112376 324374 112432
rect 324410 111696 324466 111752
rect 324318 110880 324374 110936
rect 324778 110064 324834 110120
rect 324318 109384 324374 109440
rect 324410 108568 324466 108624
rect 324318 107752 324374 107808
rect 324318 105440 324374 105496
rect 326434 178608 326490 178664
rect 325882 161608 325938 161664
rect 327538 121372 327594 121408
rect 327538 121352 327540 121372
rect 327540 121352 327592 121372
rect 327592 121352 327594 121372
rect 325514 107072 325570 107128
rect 322938 103944 322994 104000
rect 325606 103128 325662 103184
rect 324410 102448 324466 102504
rect 324594 100816 324650 100872
rect 322938 100136 322994 100192
rect 324318 99340 324374 99376
rect 324318 99320 324320 99340
rect 324320 99320 324372 99340
rect 324372 99320 324374 99340
rect 324410 98504 324466 98560
rect 324318 96328 324374 96384
rect 324318 93200 324374 93256
rect 324594 97824 324650 97880
rect 324502 93744 324558 93800
rect 327906 85448 327962 85504
rect 329930 109656 329986 109712
rect 331494 161200 331550 161256
rect 333242 274760 333298 274816
rect 340142 273808 340198 273864
rect 338118 211792 338174 211848
rect 340786 129004 340788 129024
rect 340788 129004 340840 129024
rect 340840 129004 340842 129024
rect 340786 128968 340842 129004
rect 339498 51720 339554 51776
rect 336738 42064 336794 42120
rect 338670 3440 338726 3496
rect 342442 207576 342498 207632
rect 346306 115096 346362 115152
rect 347686 285640 347742 285696
rect 347686 227568 347742 227624
rect 345018 24112 345074 24168
rect 349250 200640 349306 200696
rect 355322 357448 355378 357504
rect 353298 222808 353354 222864
rect 354770 184320 354826 184376
rect 358082 272448 358138 272504
rect 356794 228792 356850 228848
rect 357346 116456 357402 116512
rect 359554 280200 359610 280256
rect 360934 281560 360990 281616
rect 359554 234504 359610 234560
rect 359554 178744 359610 178800
rect 363694 284824 363750 284880
rect 362222 96328 362278 96384
rect 365166 278976 365222 279032
rect 368478 241440 368534 241496
rect 368478 241168 368534 241224
rect 369306 241440 369362 241496
rect 370594 237088 370650 237144
rect 371974 238584 372030 238640
rect 373998 224848 374054 224904
rect 373354 200776 373410 200832
rect 373446 128968 373502 129024
rect 377402 341400 377458 341456
rect 374734 224848 374790 224904
rect 374642 92384 374698 92440
rect 377586 280336 377642 280392
rect 376114 95104 376170 95160
rect 380346 278840 380402 278896
rect 380254 274896 380310 274952
rect 380346 237224 380402 237280
rect 380162 94968 380218 95024
rect 382278 234640 382334 234696
rect 383106 274624 383162 274680
rect 383106 235864 383162 235920
rect 383106 234640 383162 234696
rect 383014 179424 383070 179480
rect 382922 173848 382978 173904
rect 385038 279112 385094 279168
rect 384302 277616 384358 277672
rect 384486 277480 384542 277536
rect 384486 161336 384542 161392
rect 383566 91024 383622 91080
rect 386878 273400 386934 273456
rect 387154 270000 387210 270056
rect 387062 266600 387118 266656
rect 386878 263200 386934 263256
rect 386878 259936 386934 259992
rect 386878 256400 386934 256456
rect 386878 253000 386934 253056
rect 386878 246336 386934 246392
rect 386602 243516 386604 243536
rect 386604 243516 386656 243536
rect 386656 243516 386658 243536
rect 386602 243480 386658 243516
rect 386878 240216 386934 240272
rect 387522 249600 387578 249656
rect 386786 236680 386842 236736
rect 386510 233416 386566 233472
rect 386418 226616 386474 226672
rect 386970 223216 387026 223272
rect 387154 230016 387210 230072
rect 387154 223216 387210 223272
rect 387062 222128 387118 222184
rect 386878 219816 386934 219872
rect 386878 212880 386934 212936
rect 387522 216416 387578 216472
rect 386878 209480 386934 209536
rect 386878 206080 386934 206136
rect 386878 202680 386934 202736
rect 387062 199280 387118 199336
rect 386878 196016 386934 196072
rect 386418 193296 386474 193352
rect 386878 189760 386934 189816
rect 386786 186496 386842 186552
rect 386418 182960 386474 183016
rect 386878 179560 386934 179616
rect 387706 270000 387762 270056
rect 387154 172896 387210 172952
rect 386878 169496 386934 169552
rect 386878 166096 386934 166152
rect 386878 162696 386934 162752
rect 387062 159160 387118 159216
rect 386878 152496 386934 152552
rect 386602 149096 386658 149152
rect 386602 145560 386658 145616
rect 387614 142840 387670 142896
rect 387154 139440 387210 139496
rect 386694 136040 386750 136096
rect 386602 129376 386658 129432
rect 386786 122576 386842 122632
rect 386878 119176 386934 119232
rect 386878 115640 386934 115696
rect 386602 108996 386658 109032
rect 386602 108976 386604 108996
rect 386604 108976 386656 108996
rect 386656 108976 386658 108996
rect 387614 125976 387670 126032
rect 387062 106120 387118 106176
rect 386878 98776 386934 98832
rect 387614 106120 387670 106176
rect 387614 105576 387670 105632
rect 388534 277752 388590 277808
rect 388442 213832 388498 213888
rect 387798 175888 387854 175944
rect 388442 155896 388498 155952
rect 388994 216416 389050 216472
rect 391202 301416 391258 301472
rect 390466 275576 390522 275632
rect 494794 702480 494850 702536
rect 462318 311072 462374 311128
rect 444746 276256 444802 276312
rect 460202 277752 460258 277808
rect 476302 279112 476358 279168
rect 479522 277616 479578 277672
rect 510802 275984 510858 276040
rect 552294 355272 552350 355328
rect 540058 278976 540114 279032
rect 558734 277480 558790 277536
rect 580170 683848 580226 683904
rect 565818 284824 565874 284880
rect 580170 644000 580226 644056
rect 568578 354728 568634 354784
rect 568578 278704 568634 278760
rect 504362 275576 504418 275632
rect 568578 274896 568634 274952
rect 569958 264560 570014 264616
rect 569314 257624 569370 257680
rect 569958 237224 570014 237280
rect 569314 220768 569370 220824
rect 389822 162424 389878 162480
rect 569314 156032 569370 156088
rect 389086 132776 389142 132832
rect 389638 93744 389694 93800
rect 405462 92384 405518 92440
rect 408682 91024 408738 91080
rect 538770 93608 538826 93664
rect 535458 86808 535514 86864
rect 569314 97144 569370 97200
rect 570142 223896 570198 223952
rect 570234 217096 570290 217152
rect 570142 180240 570198 180296
rect 570050 106800 570106 106856
rect 570050 99456 570106 99512
rect 572718 274760 572774 274816
rect 571614 270816 571670 270872
rect 571522 267416 571578 267472
rect 572626 260616 572682 260672
rect 571430 253816 571486 253872
rect 572626 251132 572628 251152
rect 572628 251132 572680 251152
rect 572680 251132 572682 251152
rect 572626 251096 572682 251132
rect 572626 247696 572682 247752
rect 572626 240896 572682 240952
rect 572626 234096 572682 234152
rect 572626 230696 572682 230752
rect 572626 227332 572628 227352
rect 572628 227332 572680 227352
rect 572680 227332 572682 227352
rect 572626 227296 572682 227332
rect 572626 213560 572682 213616
rect 572626 210296 572682 210352
rect 572442 206932 572444 206952
rect 572444 206932 572496 206952
rect 572496 206932 572498 206952
rect 572442 206896 572498 206932
rect 571522 203496 571578 203552
rect 572626 197376 572682 197432
rect 571706 190576 571762 190632
rect 572626 187176 572682 187232
rect 571430 183776 571486 183832
rect 572074 176976 572130 177032
rect 572626 170040 572682 170096
rect 572350 166640 572406 166696
rect 571338 163376 571394 163432
rect 572626 159840 572682 159896
rect 572626 153212 572628 153232
rect 572628 153212 572680 153232
rect 572680 153212 572682 153232
rect 572626 153176 572682 153212
rect 572626 150456 572682 150512
rect 571706 147056 571762 147112
rect 572626 143556 572628 143576
rect 572628 143556 572680 143576
rect 572680 143556 572682 143576
rect 572626 143520 572682 143556
rect 572626 140120 572682 140176
rect 572626 136856 572682 136912
rect 572718 133320 572774 133376
rect 572626 130056 572682 130112
rect 571338 126520 571394 126576
rect 571246 106292 571248 106312
rect 571248 106292 571300 106312
rect 571300 106292 571302 106312
rect 571246 106256 571302 106292
rect 572626 123256 572682 123312
rect 571430 119720 571486 119776
rect 571338 96192 571394 96248
rect 572626 116456 572682 116512
rect 571522 112920 571578 112976
rect 572626 102720 572682 102776
rect 571614 96600 571670 96656
rect 571522 93744 571578 93800
rect 580170 630808 580226 630864
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 580170 537784 580226 537840
rect 574098 96464 574154 96520
rect 580262 524456 580318 524512
rect 580170 484608 580226 484664
rect 580170 471416 580226 471472
rect 578882 458088 578938 458144
rect 580170 431568 580226 431624
rect 579618 418240 579674 418296
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 576858 280336 576914 280392
rect 575478 94968 575534 95024
rect 580170 365064 580226 365120
rect 580262 354456 580318 354512
rect 580170 325216 580226 325272
rect 580354 351872 580410 351928
rect 580262 312024 580318 312080
rect 579618 298696 579674 298752
rect 579618 294480 579674 294536
rect 579618 278840 579674 278896
rect 580998 280472 581054 280528
rect 579710 276120 579766 276176
rect 580170 272176 580226 272232
rect 580170 258848 580226 258904
rect 580078 219000 580134 219056
rect 580354 192480 580410 192536
rect 580906 205692 580962 205728
rect 580906 205672 580908 205692
rect 580908 205672 580960 205692
rect 580960 205672 580962 205692
rect 580446 179152 580502 179208
rect 581642 152632 581698 152688
rect 580170 139304 580226 139360
rect 579618 125976 579674 126032
rect 579894 112784 579950 112840
rect 580170 86128 580226 86184
rect 579986 72936 580042 72992
rect 580170 59608 580226 59664
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 579618 15816 579674 15872
rect 580354 99456 580410 99512
rect 582562 697176 582618 697232
rect 582654 670656 582710 670712
rect 582562 281560 582618 281616
rect 582746 617480 582802 617536
rect 583850 563760 583906 563816
rect 582654 281424 582710 281480
rect 582746 245556 582748 245576
rect 582748 245556 582800 245576
rect 582800 245556 582802 245576
rect 582746 245520 582802 245556
rect 582654 165824 582710 165880
rect 582654 95104 582710 95160
rect 583206 281424 583262 281480
rect 583206 280200 583262 280256
rect 583114 205672 583170 205728
rect 583390 232328 583446 232384
rect 583850 193024 583906 193080
rect 583758 46824 583814 46880
rect 580262 6568 580318 6624
<< obsm2 >>
rect 68800 95100 164756 174600
<< metal3 >>
rect 295926 702476 295932 702540
rect 295996 702538 296002 702540
rect 494789 702538 494855 702541
rect 295996 702536 494855 702538
rect 295996 702480 494794 702536
rect 494850 702480 494855 702536
rect 295996 702478 494855 702480
rect 295996 702476 296002 702478
rect 494789 702475 494855 702478
rect -960 697220 480 697460
rect 582557 697234 582623 697237
rect 583520 697234 584960 697324
rect 582557 697232 584960 697234
rect 582557 697176 582562 697232
rect 582618 697176 584960 697232
rect 582557 697174 584960 697176
rect 582557 697171 582623 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 582649 670714 582715 670717
rect 583520 670714 584960 670804
rect 582649 670712 584960 670714
rect 582649 670656 582654 670712
rect 582710 670656 584960 670712
rect 582649 670654 584960 670656
rect 582649 670651 582715 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 582741 617538 582807 617541
rect 583520 617538 584960 617628
rect 582741 617536 584960 617538
rect 582741 617480 582746 617536
rect 582802 617480 584960 617536
rect 582741 617478 584960 617480
rect 582741 617475 582807 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect -960 579942 6930 580002
rect -960 579852 480 579942
rect 6870 579730 6930 579942
rect 121494 579730 121500 579732
rect 6870 579670 121500 579730
rect 121494 579668 121500 579670
rect 121564 579668 121570 579732
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 583520 564362 584960 564452
rect 583342 564302 584960 564362
rect 583342 564226 583402 564302
rect 583520 564226 584960 564302
rect 583342 564212 584960 564226
rect 583342 564166 583770 564212
rect 583710 563818 583770 564166
rect 583845 563818 583911 563821
rect 583710 563816 583911 563818
rect 583710 563760 583850 563816
rect 583906 563760 583911 563816
rect 583710 563758 583911 563760
rect 583845 563755 583911 563758
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 580257 524514 580323 524517
rect 583520 524514 584960 524604
rect 580257 524512 584960 524514
rect 580257 524456 580262 524512
rect 580318 524456 584960 524512
rect 580257 524454 584960 524456
rect 580257 524451 580323 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 579654 511260 579660 511324
rect 579724 511322 579730 511324
rect 583520 511322 584960 511412
rect 579724 511262 584960 511322
rect 579724 511260 579730 511262
rect 583520 511172 584960 511262
rect 305729 510642 305795 510645
rect 579654 510642 579660 510644
rect 305729 510640 579660 510642
rect 305729 510584 305734 510640
rect 305790 510584 579660 510640
rect 305729 510582 579660 510584
rect 305729 510579 305795 510582
rect 579654 510580 579660 510582
rect 579724 510580 579730 510644
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3233 462634 3299 462637
rect -960 462632 3299 462634
rect -960 462576 3238 462632
rect 3294 462576 3299 462632
rect -960 462574 3299 462576
rect -960 462484 480 462574
rect 3233 462571 3299 462574
rect 578877 458146 578943 458149
rect 583520 458146 584960 458236
rect 578877 458144 584960 458146
rect 578877 458088 578882 458144
rect 578938 458088 584960 458144
rect 578877 458086 584960 458088
rect 578877 458083 578943 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3417 423602 3483 423605
rect -960 423600 3483 423602
rect -960 423544 3422 423600
rect 3478 423544 3483 423600
rect -960 423542 3483 423544
rect -960 423452 480 423542
rect 3417 423539 3483 423542
rect 579613 418298 579679 418301
rect 583520 418298 584960 418388
rect 579613 418296 584960 418298
rect 579613 418240 579618 418296
rect 579674 418240 584960 418296
rect 579613 418238 584960 418240
rect 579613 418235 579679 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3141 410546 3207 410549
rect -960 410544 3207 410546
rect -960 410488 3146 410544
rect 3202 410488 3207 410544
rect -960 410486 3207 410488
rect -960 410396 480 410486
rect 3141 410483 3207 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3417 397490 3483 397493
rect -960 397488 3483 397490
rect -960 397432 3422 397488
rect 3478 397432 3483 397488
rect -960 397430 3483 397432
rect -960 397340 480 397430
rect 3417 397427 3483 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3417 371378 3483 371381
rect -960 371376 3483 371378
rect -960 371320 3422 371376
rect 3478 371320 3483 371376
rect -960 371318 3483 371320
rect -960 371228 480 371318
rect 3417 371315 3483 371318
rect 152457 365802 152523 365805
rect 295926 365802 295932 365804
rect 152457 365800 295932 365802
rect 152457 365744 152462 365800
rect 152518 365744 295932 365800
rect 152457 365742 295932 365744
rect 152457 365739 152523 365742
rect 295926 365740 295932 365742
rect 295996 365740 296002 365804
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect 213913 364442 213979 364445
rect 570086 364442 570092 364444
rect 213913 364440 570092 364442
rect 213913 364384 213918 364440
rect 213974 364384 570092 364440
rect 213913 364382 570092 364384
rect 213913 364379 213979 364382
rect 570086 364380 570092 364382
rect 570156 364380 570162 364444
rect 69054 363020 69060 363084
rect 69124 363082 69130 363084
rect 243629 363082 243695 363085
rect 69124 363080 243695 363082
rect 69124 363024 243634 363080
rect 243690 363024 243695 363080
rect 69124 363022 243695 363024
rect 69124 363020 69130 363022
rect 243629 363019 243695 363022
rect 258901 358866 258967 358869
rect 294086 358866 294092 358868
rect 258901 358864 294092 358866
rect 258901 358808 258906 358864
rect 258962 358808 294092 358864
rect 258901 358806 294092 358808
rect 258901 358803 258967 358806
rect 294086 358804 294092 358806
rect 294156 358804 294162 358868
rect -960 358458 480 358548
rect 3417 358458 3483 358461
rect -960 358456 3483 358458
rect -960 358400 3422 358456
rect 3478 358400 3483 358456
rect -960 358398 3483 358400
rect -960 358308 480 358398
rect 3417 358395 3483 358398
rect 179781 357778 179847 357781
rect 211797 357778 211863 357781
rect 179781 357776 211863 357778
rect 179781 357720 179786 357776
rect 179842 357720 211802 357776
rect 211858 357720 211863 357776
rect 179781 357718 211863 357720
rect 179781 357715 179847 357718
rect 211797 357715 211863 357718
rect 269021 357778 269087 357781
rect 324957 357778 325023 357781
rect 269021 357776 325023 357778
rect 269021 357720 269026 357776
rect 269082 357720 324962 357776
rect 325018 357720 325023 357776
rect 269021 357718 325023 357720
rect 269021 357715 269087 357718
rect 324957 357715 325023 357718
rect 193213 357642 193279 357645
rect 193857 357642 193923 357645
rect 296161 357642 296227 357645
rect 193213 357640 296227 357642
rect 193213 357584 193218 357640
rect 193274 357584 193862 357640
rect 193918 357584 296166 357640
rect 296222 357584 296227 357640
rect 193213 357582 296227 357584
rect 193213 357579 193279 357582
rect 193857 357579 193923 357582
rect 296161 357579 296227 357582
rect 130469 357506 130535 357509
rect 206277 357506 206343 357509
rect 130469 357504 206343 357506
rect 130469 357448 130474 357504
rect 130530 357448 206282 357504
rect 206338 357448 206343 357504
rect 130469 357446 206343 357448
rect 130469 357443 130535 357446
rect 206277 357443 206343 357446
rect 242157 357506 242223 357509
rect 355317 357506 355383 357509
rect 242157 357504 355383 357506
rect 242157 357448 242162 357504
rect 242218 357448 355322 357504
rect 355378 357448 355383 357504
rect 242157 357446 355383 357448
rect 242157 357443 242223 357446
rect 355317 357443 355383 357446
rect 282085 356282 282151 356285
rect 292430 356282 292436 356284
rect 282085 356280 292436 356282
rect 282085 356224 282090 356280
rect 282146 356224 292436 356280
rect 282085 356222 292436 356224
rect 282085 356219 282151 356222
rect 292430 356220 292436 356222
rect 292500 356220 292506 356284
rect 274541 356146 274607 356149
rect 335854 356146 335860 356148
rect 274541 356144 335860 356146
rect 274541 356088 274546 356144
rect 274602 356088 335860 356144
rect 274541 356086 335860 356088
rect 274541 356083 274607 356086
rect 335854 356084 335860 356086
rect 335924 356084 335930 356148
rect 201493 355330 201559 355333
rect 552289 355330 552355 355333
rect 201493 355328 552355 355330
rect 201493 355272 201498 355328
rect 201554 355272 552294 355328
rect 552350 355272 552355 355328
rect 201493 355270 552355 355272
rect 201493 355267 201559 355270
rect 552289 355267 552355 355270
rect 167494 354860 167500 354924
rect 167564 354922 167570 354924
rect 209957 354922 210023 354925
rect 167564 354920 210023 354922
rect 167564 354864 209962 354920
rect 210018 354864 210023 354920
rect 167564 354862 210023 354864
rect 167564 354860 167570 354862
rect 209957 354859 210023 354862
rect 256785 354922 256851 354925
rect 293166 354922 293172 354924
rect 256785 354920 293172 354922
rect 256785 354864 256790 354920
rect 256846 354864 293172 354920
rect 256785 354862 293172 354864
rect 256785 354859 256851 354862
rect 293166 354860 293172 354862
rect 293236 354860 293242 354924
rect 171726 354724 171732 354788
rect 171796 354786 171802 354788
rect 247033 354786 247099 354789
rect 248137 354786 248203 354789
rect 568573 354786 568639 354789
rect 171796 354784 568639 354786
rect 171796 354728 247038 354784
rect 247094 354728 248142 354784
rect 248198 354728 568578 354784
rect 568634 354728 568639 354784
rect 171796 354726 568639 354728
rect 171796 354724 171802 354726
rect 247033 354723 247099 354726
rect 248137 354723 248203 354726
rect 568573 354723 568639 354726
rect 291745 354650 291811 354653
rect 292205 354650 292271 354653
rect 291745 354648 291946 354650
rect 291745 354592 291750 354648
rect 291806 354592 291946 354648
rect 291745 354590 291946 354592
rect 291745 354587 291811 354590
rect 291886 354514 291946 354590
rect 292205 354648 296730 354650
rect 292205 354592 292210 354648
rect 292266 354592 296730 354648
rect 292205 354590 296730 354592
rect 292205 354587 292271 354590
rect 296670 354514 296730 354590
rect 580257 354514 580323 354517
rect 291886 354454 292866 354514
rect 296670 354512 580323 354514
rect 296670 354456 580262 354512
rect 580318 354456 580323 354512
rect 296670 354454 580323 354456
rect 176653 354378 176719 354381
rect 292806 354378 292866 354454
rect 580257 354451 580323 354454
rect 296069 354378 296135 354381
rect 176653 354376 180044 354378
rect 176653 354320 176658 354376
rect 176714 354320 180044 354376
rect 292806 354376 296135 354378
rect 292806 354348 296074 354376
rect 176653 354318 180044 354320
rect 292836 354320 296074 354348
rect 296130 354320 296135 354376
rect 292836 354318 296135 354320
rect 176653 354315 176719 354318
rect 296069 354315 296135 354318
rect 292614 352956 292620 353020
rect 292684 353018 292690 353020
rect 292684 352958 296730 353018
rect 292684 352956 292690 352958
rect 296670 352610 296730 352958
rect 316033 352610 316099 352613
rect 296670 352608 316099 352610
rect 296670 352552 316038 352608
rect 316094 352552 316099 352608
rect 296670 352550 316099 352552
rect 316033 352547 316099 352550
rect 295374 352338 295380 352340
rect 292836 352278 295380 352338
rect 295374 352276 295380 352278
rect 295444 352276 295450 352340
rect 179462 352210 180044 352270
rect 176561 352202 176627 352205
rect 179462 352202 179522 352210
rect 176561 352200 179522 352202
rect 176561 352144 176566 352200
rect 176622 352144 179522 352200
rect 176561 352142 179522 352144
rect 176561 352139 176627 352142
rect 580349 351930 580415 351933
rect 583520 351930 584960 352020
rect 580349 351928 584960 351930
rect 580349 351872 580354 351928
rect 580410 351872 584960 351928
rect 580349 351870 584960 351872
rect 580349 351867 580415 351870
rect 583520 351780 584960 351870
rect 179462 350170 180044 350230
rect 177062 350100 177068 350164
rect 177132 350162 177138 350164
rect 179462 350162 179522 350170
rect 177132 350102 179522 350162
rect 177132 350100 177138 350102
rect 295333 349618 295399 349621
rect 292836 349616 295399 349618
rect 292836 349560 295338 349616
rect 295394 349560 295399 349616
rect 292836 349558 295399 349560
rect 295333 349555 295399 349558
rect 179505 348190 179571 348193
rect 179505 348188 180044 348190
rect 179505 348132 179510 348188
rect 179566 348132 180044 348188
rect 179505 348130 180044 348132
rect 179505 348127 179571 348130
rect 293902 347578 293908 347580
rect 292836 347518 293908 347578
rect 293902 347516 293908 347518
rect 293972 347516 293978 347580
rect 295977 345538 296043 345541
rect 292836 345536 296043 345538
rect -960 345402 480 345492
rect 292836 345480 295982 345536
rect 296038 345480 296043 345536
rect 292836 345478 296043 345480
rect 295977 345475 296043 345478
rect 179462 345410 180044 345470
rect 3509 345402 3575 345405
rect -960 345400 3575 345402
rect -960 345344 3514 345400
rect 3570 345344 3575 345400
rect -960 345342 3575 345344
rect -960 345252 480 345342
rect 3509 345339 3575 345342
rect 176653 345402 176719 345405
rect 179462 345402 179522 345410
rect 176653 345400 179522 345402
rect 176653 345344 176658 345400
rect 176714 345344 179522 345400
rect 176653 345342 179522 345344
rect 176653 345339 176719 345342
rect 295742 343498 295748 343500
rect 292836 343438 295748 343498
rect 295742 343436 295748 343438
rect 295812 343436 295818 343500
rect 179462 343370 180044 343430
rect 176837 343362 176903 343365
rect 179462 343362 179522 343370
rect 176837 343360 179522 343362
rect 176837 343304 176842 343360
rect 176898 343304 179522 343360
rect 176837 343302 179522 343304
rect 176837 343299 176903 343302
rect 295742 341396 295748 341460
rect 295812 341458 295818 341460
rect 377397 341458 377463 341461
rect 295812 341456 377463 341458
rect 295812 341400 377402 341456
rect 377458 341400 377463 341456
rect 295812 341398 377463 341400
rect 295812 341396 295818 341398
rect 377397 341395 377463 341398
rect 179505 341390 179571 341393
rect 179505 341388 180044 341390
rect 179505 341332 179510 341388
rect 179566 341332 180044 341388
rect 179505 341330 180044 341332
rect 179505 341327 179571 341330
rect 295333 340778 295399 340781
rect 292836 340776 295399 340778
rect 292836 340720 295338 340776
rect 295394 340720 295399 340776
rect 292836 340718 295399 340720
rect 295333 340715 295399 340718
rect 179462 339290 180044 339350
rect 173750 339220 173756 339284
rect 173820 339282 173826 339284
rect 179462 339282 179522 339290
rect 173820 339222 179522 339282
rect 173820 339220 173826 339222
rect 293125 338738 293191 338741
rect 293861 338738 293927 338741
rect 292836 338736 293927 338738
rect 292836 338680 293130 338736
rect 293186 338680 293866 338736
rect 293922 338680 293927 338736
rect 292836 338678 293927 338680
rect 293125 338675 293191 338678
rect 293861 338675 293927 338678
rect 583520 338452 584960 338692
rect 295333 336698 295399 336701
rect 292836 336696 295399 336698
rect 292836 336640 295338 336696
rect 295394 336640 295399 336696
rect 292836 336638 295399 336640
rect 295333 336635 295399 336638
rect 179462 336570 180044 336630
rect 179137 336562 179203 336565
rect 179462 336562 179522 336570
rect 179137 336560 179522 336562
rect 179137 336504 179142 336560
rect 179198 336504 179522 336560
rect 179137 336502 179522 336504
rect 179137 336499 179203 336502
rect 293953 334658 294019 334661
rect 292836 334656 294019 334658
rect 292836 334600 293958 334656
rect 294014 334600 294019 334656
rect 292836 334598 294019 334600
rect 293953 334595 294019 334598
rect 179830 334530 180044 334590
rect 176837 334522 176903 334525
rect 179270 334522 179276 334524
rect 176837 334520 179276 334522
rect 176837 334464 176842 334520
rect 176898 334464 179276 334520
rect 176837 334462 179276 334464
rect 176837 334459 176903 334462
rect 179270 334460 179276 334462
rect 179340 334522 179346 334524
rect 179830 334522 179890 334530
rect 179340 334462 179890 334522
rect 179340 334460 179346 334462
rect 176653 332618 176719 332621
rect 176653 332616 179890 332618
rect 176653 332560 176658 332616
rect 176714 332560 179890 332616
rect 176653 332558 179890 332560
rect 176653 332555 176719 332558
rect 179830 332550 179890 332558
rect 179830 332490 180044 332550
rect -960 332196 480 332436
rect 295333 331938 295399 331941
rect 292836 331936 295399 331938
rect 292836 331880 295338 331936
rect 295394 331880 295399 331936
rect 292836 331878 295399 331880
rect 295333 331875 295399 331878
rect 179462 330450 180044 330510
rect 175038 330380 175044 330444
rect 175108 330442 175114 330444
rect 179462 330442 179522 330450
rect 175108 330382 179522 330442
rect 175108 330380 175114 330382
rect 294045 329898 294111 329901
rect 294321 329898 294387 329901
rect 292836 329896 294387 329898
rect 292836 329840 294050 329896
rect 294106 329840 294326 329896
rect 294382 329840 294387 329896
rect 292836 329838 294387 329840
rect 294045 329835 294111 329838
rect 294321 329835 294387 329838
rect 293033 328402 293099 328405
rect 292806 328400 293099 328402
rect 292806 328344 293038 328400
rect 293094 328344 293099 328400
rect 292806 328342 293099 328344
rect 292806 327828 292866 328342
rect 293033 328339 293099 328342
rect 179462 327730 180044 327790
rect 176653 327722 176719 327725
rect 179462 327722 179522 327730
rect 176653 327720 179522 327722
rect 176653 327664 176658 327720
rect 176714 327664 179522 327720
rect 176653 327662 179522 327664
rect 176653 327659 176719 327662
rect 176653 325818 176719 325821
rect 294137 325818 294203 325821
rect 176653 325816 179522 325818
rect 176653 325760 176658 325816
rect 176714 325760 179522 325816
rect 176653 325758 179522 325760
rect 292836 325816 294203 325818
rect 292836 325760 294142 325816
rect 294198 325760 294203 325816
rect 292836 325758 294203 325760
rect 176653 325755 176719 325758
rect 179462 325750 179522 325758
rect 294137 325755 294203 325758
rect 179462 325690 180044 325750
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 179462 323650 180044 323710
rect 176326 323580 176332 323644
rect 176396 323642 176402 323644
rect 179462 323642 179522 323650
rect 176396 323582 179522 323642
rect 176396 323580 176402 323582
rect 294229 323098 294295 323101
rect 292836 323096 294295 323098
rect 292836 323040 294234 323096
rect 294290 323040 294295 323096
rect 292836 323038 294295 323040
rect 294229 323035 294295 323038
rect 179462 321610 180044 321670
rect 177941 321602 178007 321605
rect 179462 321602 179522 321610
rect 177941 321600 179522 321602
rect 177941 321544 177946 321600
rect 178002 321544 179522 321600
rect 177941 321542 179522 321544
rect 177941 321539 178007 321542
rect 295333 321058 295399 321061
rect 292836 321056 295399 321058
rect 292836 321000 295338 321056
rect 295394 321000 295399 321056
rect 292836 320998 295399 321000
rect 295333 320995 295399 320998
rect -960 319290 480 319380
rect 3417 319290 3483 319293
rect -960 319288 3483 319290
rect -960 319232 3422 319288
rect 3478 319232 3483 319288
rect -960 319230 3483 319232
rect -960 319140 480 319230
rect 3417 319227 3483 319230
rect 295333 319018 295399 319021
rect 292836 319016 295399 319018
rect 292836 318960 295338 319016
rect 295394 318960 295399 319016
rect 292836 318958 295399 318960
rect 295333 318955 295399 318958
rect 179462 318890 180044 318950
rect 177849 318882 177915 318885
rect 179462 318882 179522 318890
rect 177849 318880 179522 318882
rect 177849 318824 177854 318880
rect 177910 318824 179522 318880
rect 177849 318822 179522 318824
rect 177849 318819 177915 318822
rect 295333 316978 295399 316981
rect 292836 316976 295399 316978
rect 292836 316920 295338 316976
rect 295394 316920 295399 316976
rect 292836 316918 295399 316920
rect 295333 316915 295399 316918
rect 179462 316850 180044 316910
rect 176510 316780 176516 316844
rect 176580 316842 176586 316844
rect 179462 316842 179522 316850
rect 176580 316782 179522 316842
rect 176580 316780 176586 316782
rect 179462 314810 180044 314870
rect 176653 314802 176719 314805
rect 179462 314802 179522 314810
rect 176653 314800 179522 314802
rect 176653 314744 176658 314800
rect 176714 314744 179522 314800
rect 176653 314742 179522 314744
rect 176653 314739 176719 314742
rect 295333 314258 295399 314261
rect 292836 314256 295399 314258
rect 292836 314200 295338 314256
rect 295394 314200 295399 314256
rect 292836 314198 295399 314200
rect 295333 314195 295399 314198
rect 179462 312770 180044 312830
rect 176653 312762 176719 312765
rect 179462 312762 179522 312770
rect 176653 312760 179522 312762
rect 176653 312704 176658 312760
rect 176714 312704 179522 312760
rect 176653 312702 179522 312704
rect 176653 312699 176719 312702
rect 160553 311946 160619 311949
rect 292622 311948 292682 312188
rect 580257 312082 580323 312085
rect 583520 312082 584960 312172
rect 580257 312080 584960 312082
rect 580257 312024 580262 312080
rect 580318 312024 584960 312080
rect 580257 312022 584960 312024
rect 580257 312019 580323 312022
rect 161238 311946 161244 311948
rect 160553 311944 161244 311946
rect 160553 311888 160558 311944
rect 160614 311888 161244 311944
rect 160553 311886 161244 311888
rect 160553 311883 160619 311886
rect 161238 311884 161244 311886
rect 161308 311884 161314 311948
rect 292614 311884 292620 311948
rect 292684 311946 292690 311948
rect 295333 311946 295399 311949
rect 292684 311944 295399 311946
rect 292684 311888 295338 311944
rect 295394 311888 295399 311944
rect 583520 311932 584960 312022
rect 292684 311886 295399 311888
rect 292684 311884 292690 311886
rect 295333 311883 295399 311886
rect 388478 311068 388484 311132
rect 388548 311130 388554 311132
rect 462313 311130 462379 311133
rect 388548 311128 462379 311130
rect 388548 311072 462318 311128
rect 462374 311072 462379 311128
rect 388548 311070 462379 311072
rect 388548 311068 388554 311070
rect 462313 311067 462379 311070
rect 295333 310178 295399 310181
rect 292836 310176 295399 310178
rect 292836 310120 295338 310176
rect 295394 310120 295399 310176
rect 292836 310118 295399 310120
rect 295333 310115 295399 310118
rect 179462 310050 180044 310110
rect 176469 310042 176535 310045
rect 179462 310042 179522 310050
rect 176469 310040 179522 310042
rect 176469 309984 176474 310040
rect 176530 309984 179522 310040
rect 176469 309982 179522 309984
rect 176469 309979 176535 309982
rect 295333 308138 295399 308141
rect 292836 308136 295399 308138
rect 292836 308080 295338 308136
rect 295394 308080 295399 308136
rect 292836 308078 295399 308080
rect 295333 308075 295399 308078
rect 179505 308070 179571 308073
rect 179505 308068 180044 308070
rect 179505 308012 179510 308068
rect 179566 308012 180044 308068
rect 179505 308010 180044 308012
rect 179505 308007 179571 308010
rect -960 306234 480 306324
rect 3233 306234 3299 306237
rect -960 306232 3299 306234
rect -960 306176 3238 306232
rect 3294 306176 3299 306232
rect -960 306174 3299 306176
rect -960 306084 480 306174
rect 3233 306171 3299 306174
rect 179462 305970 180044 306030
rect 176653 305962 176719 305965
rect 179462 305962 179522 305970
rect 176653 305960 179522 305962
rect 176653 305904 176658 305960
rect 176714 305904 179522 305960
rect 176653 305902 179522 305904
rect 176653 305899 176719 305902
rect 295333 305418 295399 305421
rect 292836 305416 295399 305418
rect 292836 305360 295338 305416
rect 295394 305360 295399 305416
rect 292836 305358 295399 305360
rect 295333 305355 295399 305358
rect 179462 303930 180044 303990
rect 179229 303922 179295 303925
rect 179462 303922 179522 303930
rect 179229 303920 179522 303922
rect 179229 303864 179234 303920
rect 179290 303864 179522 303920
rect 179229 303862 179522 303864
rect 179229 303859 179295 303862
rect 295333 303378 295399 303381
rect 292836 303376 295399 303378
rect 292836 303320 295338 303376
rect 295394 303320 295399 303376
rect 292836 303318 295399 303320
rect 295333 303315 295399 303318
rect 387006 301412 387012 301476
rect 387076 301474 387082 301476
rect 391197 301474 391263 301477
rect 387076 301472 391263 301474
rect 387076 301416 391202 301472
rect 391258 301416 391263 301472
rect 387076 301414 391263 301416
rect 387076 301412 387082 301414
rect 391197 301411 391263 301414
rect 293217 301338 293283 301341
rect 292836 301336 293283 301338
rect 292836 301280 293222 301336
rect 293278 301280 293283 301336
rect 292836 301278 293283 301280
rect 293217 301275 293283 301278
rect 179462 301210 180044 301270
rect 176653 301202 176719 301205
rect 179462 301202 179522 301210
rect 176653 301200 179522 301202
rect 176653 301144 176658 301200
rect 176714 301144 179522 301200
rect 176653 301142 179522 301144
rect 176653 301139 176719 301142
rect 149697 299436 149763 299437
rect 149646 299434 149652 299436
rect 149606 299374 149652 299434
rect 149716 299432 149763 299436
rect 149758 299376 149763 299432
rect 149646 299372 149652 299374
rect 149716 299372 149763 299376
rect 149697 299371 149763 299372
rect 293953 299298 294019 299301
rect 292836 299296 294019 299298
rect 292836 299240 293958 299296
rect 294014 299240 294019 299296
rect 292836 299238 294019 299240
rect 293953 299235 294019 299238
rect 179462 299170 180044 299230
rect 176653 299162 176719 299165
rect 179462 299162 179522 299170
rect 176653 299160 179522 299162
rect 176653 299104 176658 299160
rect 176714 299104 179522 299160
rect 176653 299102 179522 299104
rect 176653 299099 176719 299102
rect 293166 298692 293172 298756
rect 293236 298754 293242 298756
rect 579613 298754 579679 298757
rect 583520 298754 584960 298844
rect 293236 298752 584960 298754
rect 293236 298696 579618 298752
rect 579674 298696 584960 298752
rect 293236 298694 584960 298696
rect 293236 298692 293242 298694
rect 579613 298691 579679 298694
rect 583520 298604 584960 298694
rect 97717 298346 97783 298349
rect 167678 298346 167684 298348
rect 97717 298344 167684 298346
rect 97717 298288 97722 298344
rect 97778 298288 167684 298344
rect 97717 298286 167684 298288
rect 97717 298283 97783 298286
rect 167678 298284 167684 298286
rect 167748 298284 167754 298348
rect 64597 298210 64663 298213
rect 149646 298210 149652 298212
rect 64597 298208 149652 298210
rect 64597 298152 64602 298208
rect 64658 298152 149652 298208
rect 64597 298150 149652 298152
rect 64597 298147 64663 298150
rect 149646 298148 149652 298150
rect 149716 298148 149722 298212
rect 66110 297332 66116 297396
rect 66180 297394 66186 297396
rect 169753 297394 169819 297397
rect 66180 297392 169819 297394
rect 66180 297336 169758 297392
rect 169814 297336 169819 297392
rect 66180 297334 169819 297336
rect 66180 297332 66186 297334
rect 169753 297331 169819 297334
rect 176653 297258 176719 297261
rect 176653 297256 179522 297258
rect 176653 297200 176658 297256
rect 176714 297200 179522 297256
rect 176653 297198 179522 297200
rect 176653 297195 176719 297198
rect 179462 297190 179522 297198
rect 179462 297130 180044 297190
rect 94589 296986 94655 296989
rect 166206 296986 166212 296988
rect 94589 296984 166212 296986
rect 94589 296928 94594 296984
rect 94650 296928 166212 296984
rect 94589 296926 166212 296928
rect 94589 296923 94655 296926
rect 166206 296924 166212 296926
rect 166276 296924 166282 296988
rect 158437 296852 158503 296853
rect 158437 296848 158484 296852
rect 158548 296850 158554 296852
rect 158437 296792 158442 296848
rect 158437 296788 158484 296792
rect 158548 296790 158594 296850
rect 158548 296788 158554 296790
rect 158437 296787 158503 296788
rect 295333 296578 295399 296581
rect 292836 296576 295399 296578
rect 292836 296520 295338 296576
rect 295394 296520 295399 296576
rect 292836 296518 295399 296520
rect 295333 296515 295399 296518
rect 95141 296034 95207 296037
rect 129641 296034 129707 296037
rect 95141 296032 129707 296034
rect 95141 295976 95146 296032
rect 95202 295976 129646 296032
rect 129702 295976 129707 296032
rect 95141 295974 129707 295976
rect 95141 295971 95207 295974
rect 129641 295971 129707 295974
rect 111241 295354 111307 295357
rect 127617 295354 127683 295357
rect 111241 295352 127683 295354
rect 111241 295296 111246 295352
rect 111302 295296 127622 295352
rect 127678 295296 127683 295352
rect 111241 295294 127683 295296
rect 111241 295291 111307 295294
rect 127617 295291 127683 295294
rect 179462 295090 180044 295150
rect 176653 295082 176719 295085
rect 179462 295082 179522 295090
rect 176653 295080 179522 295082
rect 176653 295024 176658 295080
rect 176714 295024 179522 295080
rect 176653 295022 179522 295024
rect 176653 295019 176719 295022
rect 73889 294538 73955 294541
rect 98729 294538 98795 294541
rect 295333 294538 295399 294541
rect 73889 294536 98795 294538
rect 73889 294480 73894 294536
rect 73950 294480 98734 294536
rect 98790 294480 98795 294536
rect 73889 294478 98795 294480
rect 292836 294536 295399 294538
rect 292836 294480 295338 294536
rect 295394 294480 295399 294536
rect 292836 294478 295399 294480
rect 73889 294475 73955 294478
rect 98729 294475 98795 294478
rect 295333 294475 295399 294478
rect 574686 294476 574692 294540
rect 574756 294538 574762 294540
rect 579613 294538 579679 294541
rect 574756 294536 579679 294538
rect 574756 294480 579618 294536
rect 579674 294480 579679 294536
rect 574756 294478 579679 294480
rect 574756 294476 574762 294478
rect 579613 294475 579679 294478
rect 103513 294266 103579 294269
rect 120901 294266 120967 294269
rect 103513 294264 120967 294266
rect 103513 294208 103518 294264
rect 103574 294208 120906 294264
rect 120962 294208 120967 294264
rect 103513 294206 120967 294208
rect 103513 294203 103579 294206
rect 120901 294203 120967 294206
rect 95785 294130 95851 294133
rect 117221 294130 117287 294133
rect 95785 294128 117287 294130
rect 95785 294072 95790 294128
rect 95846 294072 117226 294128
rect 117282 294072 117287 294128
rect 95785 294070 117287 294072
rect 95785 294067 95851 294070
rect 117221 294067 117287 294070
rect 117681 294130 117747 294133
rect 170254 294130 170260 294132
rect 117681 294128 170260 294130
rect 117681 294072 117686 294128
rect 117742 294072 170260 294128
rect 117681 294070 170260 294072
rect 117681 294067 117747 294070
rect 170254 294068 170260 294070
rect 170324 294068 170330 294132
rect 106733 293994 106799 293997
rect 170489 293994 170555 293997
rect 106733 293992 170555 293994
rect 106733 293936 106738 293992
rect 106794 293936 170494 293992
rect 170550 293936 170555 293992
rect 106733 293934 170555 293936
rect 106733 293931 106799 293934
rect 170489 293931 170555 293934
rect -960 293178 480 293268
rect 3417 293178 3483 293181
rect -960 293176 3483 293178
rect -960 293120 3422 293176
rect 3478 293120 3483 293176
rect -960 293118 3483 293120
rect -960 293028 480 293118
rect 3417 293115 3483 293118
rect 66897 293042 66963 293045
rect 126094 293042 126100 293044
rect 66897 293040 126100 293042
rect 66897 292984 66902 293040
rect 66958 292984 126100 293040
rect 66897 292982 126100 292984
rect 66897 292979 66963 292982
rect 126094 292980 126100 292982
rect 126164 292980 126170 293044
rect 108021 292906 108087 292909
rect 146886 292906 146892 292908
rect 108021 292904 146892 292906
rect 108021 292848 108026 292904
rect 108082 292848 146892 292904
rect 108021 292846 146892 292848
rect 108021 292843 108087 292846
rect 146886 292844 146892 292846
rect 146956 292844 146962 292908
rect 77753 292770 77819 292773
rect 120809 292770 120875 292773
rect 77753 292768 120875 292770
rect 77753 292712 77758 292768
rect 77814 292712 120814 292768
rect 120870 292712 120875 292768
rect 77753 292710 120875 292712
rect 77753 292707 77819 292710
rect 120809 292707 120875 292710
rect 64638 292572 64644 292636
rect 64708 292634 64714 292636
rect 70669 292634 70735 292637
rect 64708 292632 70735 292634
rect 64708 292576 70674 292632
rect 70730 292576 70735 292632
rect 64708 292574 70735 292576
rect 64708 292572 64714 292574
rect 70669 292571 70735 292574
rect 296621 292498 296687 292501
rect 292836 292496 296687 292498
rect 292836 292440 296626 292496
rect 296682 292440 296687 292496
rect 292836 292438 296687 292440
rect 296621 292435 296687 292438
rect 179462 292370 180044 292430
rect 71681 292362 71747 292365
rect 70718 292360 71747 292362
rect 70718 292304 71686 292360
rect 71742 292304 71747 292360
rect 70718 292302 71747 292304
rect 70718 291788 70778 292302
rect 71681 292299 71747 292302
rect 176377 292362 176443 292365
rect 179462 292362 179522 292370
rect 176377 292360 179522 292362
rect 176377 292304 176382 292360
rect 176438 292304 179522 292360
rect 176377 292302 179522 292304
rect 176377 292299 176443 292302
rect 114185 291954 114251 291957
rect 145649 291954 145715 291957
rect 114185 291952 145715 291954
rect 114185 291896 114190 291952
rect 114246 291896 145654 291952
rect 145710 291896 145715 291952
rect 114185 291894 145715 291896
rect 114185 291891 114251 291894
rect 145649 291891 145715 291894
rect 121453 291818 121519 291821
rect 119876 291816 121519 291818
rect 119876 291760 121458 291816
rect 121514 291760 121519 291816
rect 119876 291758 121519 291760
rect 121453 291755 121519 291758
rect 68737 291138 68803 291141
rect 121453 291138 121519 291141
rect 68737 291136 70196 291138
rect 68737 291080 68742 291136
rect 68798 291080 70196 291136
rect 68737 291078 70196 291080
rect 119876 291136 121519 291138
rect 119876 291080 121458 291136
rect 121514 291080 121519 291136
rect 119876 291078 121519 291080
rect 68737 291075 68803 291078
rect 121453 291075 121519 291078
rect 67633 290458 67699 290461
rect 121545 290458 121611 290461
rect 296069 290458 296135 290461
rect 67633 290456 70196 290458
rect 67633 290400 67638 290456
rect 67694 290400 70196 290456
rect 67633 290398 70196 290400
rect 119876 290456 121611 290458
rect 119876 290400 121550 290456
rect 121606 290400 121611 290456
rect 119876 290398 121611 290400
rect 292836 290456 296135 290458
rect 292836 290400 296074 290456
rect 296130 290400 296135 290456
rect 292836 290398 296135 290400
rect 67633 290395 67699 290398
rect 121545 290395 121611 290398
rect 296069 290395 296135 290398
rect 179462 290330 180044 290390
rect 176653 290322 176719 290325
rect 179462 290322 179522 290330
rect 176653 290320 179522 290322
rect 176653 290264 176658 290320
rect 176714 290264 179522 290320
rect 176653 290262 179522 290264
rect 176653 290259 176719 290262
rect 67725 289778 67791 289781
rect 121453 289778 121519 289781
rect 67725 289776 70196 289778
rect 67725 289720 67730 289776
rect 67786 289720 70196 289776
rect 67725 289718 70196 289720
rect 119876 289776 121519 289778
rect 119876 289720 121458 289776
rect 121514 289720 121519 289776
rect 119876 289718 121519 289720
rect 67725 289715 67791 289718
rect 121453 289715 121519 289718
rect 67633 289098 67699 289101
rect 122005 289098 122071 289101
rect 67633 289096 70196 289098
rect 67633 289040 67638 289096
rect 67694 289040 70196 289096
rect 67633 289038 70196 289040
rect 119876 289096 122071 289098
rect 119876 289040 122010 289096
rect 122066 289040 122071 289096
rect 119876 289038 122071 289040
rect 67633 289035 67699 289038
rect 122005 289035 122071 289038
rect 68829 288418 68895 288421
rect 121545 288418 121611 288421
rect 68829 288416 70196 288418
rect 68829 288360 68834 288416
rect 68890 288360 70196 288416
rect 68829 288358 70196 288360
rect 119876 288416 121611 288418
rect 119876 288360 121550 288416
rect 121606 288360 121611 288416
rect 119876 288358 121611 288360
rect 68829 288355 68895 288358
rect 121545 288355 121611 288358
rect 178677 288418 178743 288421
rect 178677 288416 179522 288418
rect 178677 288360 178682 288416
rect 178738 288360 179522 288416
rect 178677 288358 179522 288360
rect 178677 288355 178743 288358
rect 179462 288350 179522 288358
rect 179462 288290 180044 288350
rect 67633 287738 67699 287741
rect 121453 287738 121519 287741
rect 293125 287738 293191 287741
rect 67633 287736 70196 287738
rect 67633 287680 67638 287736
rect 67694 287680 70196 287736
rect 67633 287678 70196 287680
rect 119876 287736 121519 287738
rect 119876 287680 121458 287736
rect 121514 287680 121519 287736
rect 119876 287678 121519 287680
rect 292836 287736 293191 287738
rect 292836 287680 293130 287736
rect 293186 287680 293191 287736
rect 292836 287678 293191 287680
rect 67633 287675 67699 287678
rect 121453 287675 121519 287678
rect 293125 287675 293191 287678
rect 67725 287058 67791 287061
rect 121637 287058 121703 287061
rect 67725 287056 70196 287058
rect 67725 287000 67730 287056
rect 67786 287000 70196 287056
rect 67725 286998 70196 287000
rect 119876 287056 121703 287058
rect 119876 287000 121642 287056
rect 121698 287000 121703 287056
rect 119876 286998 121703 287000
rect 67725 286995 67791 286998
rect 121637 286995 121703 286998
rect 66897 286378 66963 286381
rect 121453 286378 121519 286381
rect 66897 286376 70196 286378
rect 66897 286320 66902 286376
rect 66958 286320 70196 286376
rect 66897 286318 70196 286320
rect 119876 286376 121519 286378
rect 119876 286320 121458 286376
rect 121514 286320 121519 286376
rect 119876 286318 121519 286320
rect 66897 286315 66963 286318
rect 121453 286315 121519 286318
rect 179462 286250 180044 286310
rect 176653 286242 176719 286245
rect 179462 286242 179522 286250
rect 176653 286240 179522 286242
rect 176653 286184 176658 286240
rect 176714 286184 179522 286240
rect 176653 286182 179522 286184
rect 176653 286179 176719 286182
rect 67633 285698 67699 285701
rect 122097 285698 122163 285701
rect 295333 285698 295399 285701
rect 67633 285696 70196 285698
rect 67633 285640 67638 285696
rect 67694 285640 70196 285696
rect 67633 285638 70196 285640
rect 119876 285696 122163 285698
rect 119876 285640 122102 285696
rect 122158 285640 122163 285696
rect 119876 285638 122163 285640
rect 292836 285696 295399 285698
rect 292836 285640 295338 285696
rect 295394 285640 295399 285696
rect 292836 285638 295399 285640
rect 67633 285635 67699 285638
rect 122097 285635 122163 285638
rect 295333 285635 295399 285638
rect 347681 285698 347747 285701
rect 568614 285698 568620 285700
rect 347681 285696 568620 285698
rect 347681 285640 347686 285696
rect 347742 285640 568620 285696
rect 347681 285638 568620 285640
rect 347681 285635 347747 285638
rect 568614 285636 568620 285638
rect 568684 285636 568690 285700
rect 583520 285276 584960 285516
rect 68553 285018 68619 285021
rect 121545 285018 121611 285021
rect 68553 285016 70196 285018
rect 68553 284960 68558 285016
rect 68614 284960 70196 285016
rect 68553 284958 70196 284960
rect 119876 285016 121611 285018
rect 119876 284960 121550 285016
rect 121606 284960 121611 285016
rect 119876 284958 121611 284960
rect 68553 284955 68619 284958
rect 121545 284955 121611 284958
rect 363689 284882 363755 284885
rect 565813 284882 565879 284885
rect 571558 284882 571564 284884
rect 363689 284880 571564 284882
rect 363689 284824 363694 284880
rect 363750 284824 565818 284880
rect 565874 284824 571564 284880
rect 363689 284822 571564 284824
rect 363689 284819 363755 284822
rect 565813 284819 565879 284822
rect 571558 284820 571564 284822
rect 571628 284820 571634 284884
rect 67633 284338 67699 284341
rect 121453 284338 121519 284341
rect 67633 284336 70196 284338
rect 67633 284280 67638 284336
rect 67694 284280 70196 284336
rect 67633 284278 70196 284280
rect 119876 284336 121519 284338
rect 119876 284280 121458 284336
rect 121514 284280 121519 284336
rect 119876 284278 121519 284280
rect 67633 284275 67699 284278
rect 121453 284275 121519 284278
rect 67725 283658 67791 283661
rect 295333 283658 295399 283661
rect 67725 283656 70196 283658
rect 67725 283600 67730 283656
rect 67786 283600 70196 283656
rect 292836 283656 295399 283658
rect 67725 283598 70196 283600
rect 67725 283595 67791 283598
rect 119846 283250 119906 283628
rect 292836 283600 295338 283656
rect 295394 283600 295399 283656
rect 292836 283598 295399 283600
rect 295333 283595 295399 283598
rect 179462 283530 180044 283590
rect 176653 283522 176719 283525
rect 179462 283522 179522 283530
rect 176653 283520 179522 283522
rect 176653 283464 176658 283520
rect 176714 283464 179522 283520
rect 176653 283462 179522 283464
rect 176653 283459 176719 283462
rect 178534 283250 178540 283252
rect 119846 283190 178540 283250
rect 178534 283188 178540 283190
rect 178604 283188 178610 283252
rect 67817 282978 67883 282981
rect 121453 282978 121519 282981
rect 67817 282976 70196 282978
rect 67817 282920 67822 282976
rect 67878 282920 70196 282976
rect 67817 282918 70196 282920
rect 119876 282976 121519 282978
rect 119876 282920 121458 282976
rect 121514 282920 121519 282976
rect 119876 282918 121519 282920
rect 67817 282915 67883 282918
rect 121453 282915 121519 282918
rect 120809 282298 120875 282301
rect 119876 282296 120875 282298
rect 119876 282240 120814 282296
rect 120870 282240 120875 282296
rect 119876 282238 120875 282240
rect 120809 282235 120875 282238
rect 67633 281618 67699 281621
rect 121453 281618 121519 281621
rect 67633 281616 70196 281618
rect 67633 281560 67638 281616
rect 67694 281560 70196 281616
rect 67633 281558 70196 281560
rect 119876 281616 121519 281618
rect 119876 281560 121458 281616
rect 121514 281560 121519 281616
rect 119876 281558 121519 281560
rect 67633 281555 67699 281558
rect 121453 281555 121519 281558
rect 176653 281618 176719 281621
rect 295333 281618 295399 281621
rect 176653 281616 179522 281618
rect 176653 281560 176658 281616
rect 176714 281560 179522 281616
rect 176653 281558 179522 281560
rect 292836 281616 295399 281618
rect 292836 281560 295338 281616
rect 295394 281560 295399 281616
rect 292836 281558 295399 281560
rect 176653 281555 176719 281558
rect 179462 281550 179522 281558
rect 295333 281555 295399 281558
rect 360929 281618 360995 281621
rect 582557 281618 582623 281621
rect 360929 281616 582623 281618
rect 360929 281560 360934 281616
rect 360990 281560 582562 281616
rect 582618 281560 582623 281616
rect 360929 281558 582623 281560
rect 360929 281555 360995 281558
rect 582557 281555 582623 281558
rect 179462 281490 180044 281550
rect 582649 281482 582715 281485
rect 583201 281482 583267 281485
rect 582649 281480 583267 281482
rect 582649 281424 582654 281480
rect 582710 281424 583206 281480
rect 583262 281424 583267 281480
rect 582649 281422 583267 281424
rect 582649 281419 582715 281422
rect 583201 281419 583267 281422
rect 68277 280938 68343 280941
rect 122373 280938 122439 280941
rect 68277 280936 70196 280938
rect 68277 280880 68282 280936
rect 68338 280880 70196 280936
rect 68277 280878 70196 280880
rect 119876 280936 122439 280938
rect 119876 280880 122378 280936
rect 122434 280880 122439 280936
rect 119876 280878 122439 280880
rect 68277 280875 68343 280878
rect 122373 280875 122439 280878
rect 390686 280468 390692 280532
rect 390756 280530 390762 280532
rect 580993 280530 581059 280533
rect 390756 280528 581059 280530
rect 390756 280472 580998 280528
rect 581054 280472 581059 280528
rect 390756 280470 581059 280472
rect 390756 280468 390762 280470
rect 580993 280467 581059 280470
rect 377581 280394 377647 280397
rect 576853 280394 576919 280397
rect 377581 280392 576919 280394
rect 377581 280336 377586 280392
rect 377642 280336 576858 280392
rect 576914 280336 576919 280392
rect 377581 280334 576919 280336
rect 377581 280331 377647 280334
rect 576853 280331 576919 280334
rect 67633 280258 67699 280261
rect 121453 280258 121519 280261
rect 67633 280256 70196 280258
rect -960 279972 480 280212
rect 67633 280200 67638 280256
rect 67694 280200 70196 280256
rect 67633 280198 70196 280200
rect 119876 280256 121519 280258
rect 119876 280200 121458 280256
rect 121514 280200 121519 280256
rect 119876 280198 121519 280200
rect 67633 280195 67699 280198
rect 121453 280195 121519 280198
rect 359549 280258 359615 280261
rect 583201 280258 583267 280261
rect 359549 280256 583267 280258
rect 359549 280200 359554 280256
rect 359610 280200 583206 280256
rect 583262 280200 583267 280256
rect 359549 280198 583267 280200
rect 359549 280195 359615 280198
rect 583201 280195 583267 280198
rect 67633 279578 67699 279581
rect 121545 279578 121611 279581
rect 67633 279576 70196 279578
rect 67633 279520 67638 279576
rect 67694 279520 70196 279576
rect 67633 279518 70196 279520
rect 119876 279576 121611 279578
rect 119876 279520 121550 279576
rect 121606 279520 121611 279576
rect 119876 279518 121611 279520
rect 67633 279515 67699 279518
rect 121545 279515 121611 279518
rect 176653 279578 176719 279581
rect 176653 279576 179522 279578
rect 176653 279520 176658 279576
rect 176714 279520 179522 279576
rect 176653 279518 179522 279520
rect 176653 279515 176719 279518
rect 179462 279510 179522 279518
rect 179462 279450 180044 279510
rect 385033 279170 385099 279173
rect 476297 279170 476363 279173
rect 385033 279168 476363 279170
rect 385033 279112 385038 279168
rect 385094 279112 476302 279168
rect 476358 279112 476363 279168
rect 385033 279110 476363 279112
rect 385033 279107 385099 279110
rect 476297 279107 476363 279110
rect 365161 279034 365227 279037
rect 540053 279034 540119 279037
rect 365161 279032 540119 279034
rect 365161 278976 365166 279032
rect 365222 278976 540058 279032
rect 540114 278976 540119 279032
rect 365161 278974 540119 278976
rect 365161 278971 365227 278974
rect 540053 278971 540119 278974
rect 67541 278898 67607 278901
rect 121453 278898 121519 278901
rect 295333 278898 295399 278901
rect 67541 278896 70196 278898
rect 67541 278840 67546 278896
rect 67602 278840 70196 278896
rect 67541 278838 70196 278840
rect 119876 278896 121519 278898
rect 119876 278840 121458 278896
rect 121514 278840 121519 278896
rect 119876 278838 121519 278840
rect 292836 278896 295399 278898
rect 292836 278840 295338 278896
rect 295394 278840 295399 278896
rect 292836 278838 295399 278840
rect 67541 278835 67607 278838
rect 121453 278835 121519 278838
rect 295333 278835 295399 278838
rect 380341 278898 380407 278901
rect 579613 278898 579679 278901
rect 380341 278896 579679 278898
rect 380341 278840 380346 278896
rect 380402 278840 579618 278896
rect 579674 278840 579679 278896
rect 380341 278838 579679 278840
rect 380341 278835 380407 278838
rect 579613 278835 579679 278838
rect 568573 278762 568639 278765
rect 569534 278762 569540 278764
rect 568573 278760 569540 278762
rect 568573 278704 568578 278760
rect 568634 278704 569540 278760
rect 568573 278702 569540 278704
rect 568573 278699 568639 278702
rect 569534 278700 569540 278702
rect 569604 278700 569610 278764
rect 68093 278218 68159 278221
rect 121545 278218 121611 278221
rect 68093 278216 70196 278218
rect 68093 278160 68098 278216
rect 68154 278160 70196 278216
rect 68093 278158 70196 278160
rect 119876 278216 121611 278218
rect 119876 278160 121550 278216
rect 121606 278160 121611 278216
rect 119876 278158 121611 278160
rect 68093 278155 68159 278158
rect 121545 278155 121611 278158
rect 388529 277810 388595 277813
rect 460197 277810 460263 277813
rect 388529 277808 460263 277810
rect 388529 277752 388534 277808
rect 388590 277752 460202 277808
rect 460258 277752 460263 277808
rect 388529 277750 460263 277752
rect 388529 277747 388595 277750
rect 460197 277747 460263 277750
rect 384297 277674 384363 277677
rect 479517 277674 479583 277677
rect 384297 277672 479583 277674
rect 384297 277616 384302 277672
rect 384358 277616 479522 277672
rect 479578 277616 479583 277672
rect 384297 277614 479583 277616
rect 384297 277611 384363 277614
rect 479517 277611 479583 277614
rect 67633 277538 67699 277541
rect 121453 277538 121519 277541
rect 67633 277536 70196 277538
rect 67633 277480 67638 277536
rect 67694 277480 70196 277536
rect 67633 277478 70196 277480
rect 119876 277536 121519 277538
rect 119876 277480 121458 277536
rect 121514 277480 121519 277536
rect 119876 277478 121519 277480
rect 67633 277475 67699 277478
rect 121453 277475 121519 277478
rect 176653 277538 176719 277541
rect 384481 277538 384547 277541
rect 558729 277538 558795 277541
rect 176653 277536 179522 277538
rect 176653 277480 176658 277536
rect 176714 277480 179522 277536
rect 176653 277478 179522 277480
rect 176653 277475 176719 277478
rect 179462 277470 179522 277478
rect 384481 277536 558795 277538
rect 384481 277480 384486 277536
rect 384542 277480 558734 277536
rect 558790 277480 558795 277536
rect 384481 277478 558795 277480
rect 384481 277475 384547 277478
rect 558729 277475 558795 277478
rect 179462 277410 180044 277470
rect 67725 276858 67791 276861
rect 121545 276858 121611 276861
rect 295333 276858 295399 276861
rect 67725 276856 70196 276858
rect 67725 276800 67730 276856
rect 67786 276800 70196 276856
rect 67725 276798 70196 276800
rect 119876 276856 121611 276858
rect 119876 276800 121550 276856
rect 121606 276800 121611 276856
rect 119876 276798 121611 276800
rect 292836 276856 295399 276858
rect 292836 276800 295338 276856
rect 295394 276800 295399 276856
rect 292836 276798 295399 276800
rect 67725 276795 67791 276798
rect 121545 276795 121611 276798
rect 295333 276795 295399 276798
rect 385534 276252 385540 276316
rect 385604 276314 385610 276316
rect 444741 276314 444807 276317
rect 385604 276312 444807 276314
rect 385604 276256 444746 276312
rect 444802 276256 444807 276312
rect 385604 276254 444807 276256
rect 385604 276252 385610 276254
rect 444741 276251 444807 276254
rect 67633 276178 67699 276181
rect 121453 276178 121519 276181
rect 67633 276176 70196 276178
rect 67633 276120 67638 276176
rect 67694 276120 70196 276176
rect 67633 276118 70196 276120
rect 119876 276176 121519 276178
rect 119876 276120 121458 276176
rect 121514 276120 121519 276176
rect 119876 276118 121519 276120
rect 67633 276115 67699 276118
rect 121453 276115 121519 276118
rect 389766 276116 389772 276180
rect 389836 276178 389842 276180
rect 579705 276178 579771 276181
rect 389836 276176 579771 276178
rect 389836 276120 579710 276176
rect 579766 276120 579771 276176
rect 389836 276118 579771 276120
rect 389836 276116 389842 276118
rect 579705 276115 579771 276118
rect 293166 275980 293172 276044
rect 293236 276042 293242 276044
rect 510797 276042 510863 276045
rect 293236 276040 510863 276042
rect 293236 275984 510802 276040
rect 510858 275984 510863 276040
rect 293236 275982 510863 275984
rect 293236 275980 293242 275982
rect 510797 275979 510863 275982
rect 390461 275636 390527 275637
rect 390461 275632 390508 275636
rect 390572 275634 390578 275636
rect 390461 275576 390466 275632
rect 390461 275572 390508 275576
rect 390572 275574 390618 275634
rect 390572 275572 390578 275574
rect 502006 275572 502012 275636
rect 502076 275634 502082 275636
rect 504357 275634 504423 275637
rect 502076 275632 504423 275634
rect 502076 275576 504362 275632
rect 504418 275576 504423 275632
rect 502076 275574 504423 275576
rect 502076 275572 502082 275574
rect 390461 275571 390527 275572
rect 504357 275571 504423 275574
rect 67633 275498 67699 275501
rect 121545 275498 121611 275501
rect 67633 275496 70196 275498
rect 67633 275440 67638 275496
rect 67694 275440 70196 275496
rect 67633 275438 70196 275440
rect 119876 275496 121611 275498
rect 119876 275440 121550 275496
rect 121606 275440 121611 275496
rect 119876 275438 121611 275440
rect 67633 275435 67699 275438
rect 121545 275435 121611 275438
rect 380249 274954 380315 274957
rect 568573 274954 568639 274957
rect 380249 274952 568639 274954
rect 380249 274896 380254 274952
rect 380310 274896 568578 274952
rect 568634 274896 568639 274952
rect 380249 274894 568639 274896
rect 380249 274891 380315 274894
rect 568573 274891 568639 274894
rect 67449 274818 67515 274821
rect 121453 274818 121519 274821
rect 67449 274816 70196 274818
rect 67449 274760 67454 274816
rect 67510 274760 70196 274816
rect 67449 274758 70196 274760
rect 119876 274816 121519 274818
rect 119876 274760 121458 274816
rect 121514 274760 121519 274816
rect 119876 274758 121519 274760
rect 67449 274755 67515 274758
rect 121453 274755 121519 274758
rect 177481 274818 177547 274821
rect 295333 274818 295399 274821
rect 177481 274816 179890 274818
rect 177481 274760 177486 274816
rect 177542 274760 179890 274816
rect 177481 274758 179890 274760
rect 292836 274816 295399 274818
rect 292836 274760 295338 274816
rect 295394 274760 295399 274816
rect 292836 274758 295399 274760
rect 177481 274755 177547 274758
rect 179830 274750 179890 274758
rect 295333 274755 295399 274758
rect 333237 274818 333303 274821
rect 572713 274818 572779 274821
rect 333237 274816 572779 274818
rect 333237 274760 333242 274816
rect 333298 274760 572718 274816
rect 572774 274760 572779 274816
rect 333237 274758 572779 274760
rect 333237 274755 333303 274758
rect 572713 274755 572779 274758
rect 179830 274690 180044 274750
rect 383101 274682 383167 274685
rect 502006 274682 502012 274684
rect 383101 274680 502012 274682
rect 383101 274624 383106 274680
rect 383162 274624 502012 274680
rect 383101 274622 502012 274624
rect 383101 274619 383167 274622
rect 502006 274620 502012 274622
rect 502076 274620 502082 274684
rect 568614 274484 568620 274548
rect 568684 274546 568690 274548
rect 568684 274486 569418 274546
rect 568684 274484 568690 274486
rect 390502 274274 390508 274276
rect 373950 274214 390508 274274
rect 67725 274138 67791 274141
rect 121453 274138 121519 274141
rect 67725 274136 70196 274138
rect 67725 274080 67730 274136
rect 67786 274080 70196 274136
rect 67725 274078 70196 274080
rect 119876 274136 121519 274138
rect 119876 274080 121458 274136
rect 121514 274080 121519 274136
rect 119876 274078 121519 274080
rect 67725 274075 67791 274078
rect 121453 274075 121519 274078
rect 340137 273866 340203 273869
rect 373950 273866 374010 274214
rect 390502 274212 390508 274214
rect 390572 274212 390578 274276
rect 569358 274244 569418 274486
rect 340137 273864 374010 273866
rect 340137 273808 340142 273864
rect 340198 273808 374010 273864
rect 340137 273806 374010 273808
rect 340137 273803 340203 273806
rect 67633 273458 67699 273461
rect 121453 273458 121519 273461
rect 67633 273456 70196 273458
rect 67633 273400 67638 273456
rect 67694 273400 70196 273456
rect 67633 273398 70196 273400
rect 119876 273456 121519 273458
rect 119876 273400 121458 273456
rect 121514 273400 121519 273456
rect 119876 273398 121519 273400
rect 67633 273395 67699 273398
rect 121453 273395 121519 273398
rect 386873 273458 386939 273461
rect 386873 273456 390172 273458
rect 386873 273400 386878 273456
rect 386934 273400 390172 273456
rect 386873 273398 390172 273400
rect 386873 273395 386939 273398
rect 67633 272778 67699 272781
rect 121494 272778 121500 272780
rect 67633 272776 70196 272778
rect 67633 272720 67638 272776
rect 67694 272720 70196 272776
rect 67633 272718 70196 272720
rect 119876 272718 121500 272778
rect 67633 272715 67699 272718
rect 121494 272716 121500 272718
rect 121564 272778 121570 272780
rect 122281 272778 122347 272781
rect 295333 272778 295399 272781
rect 121564 272776 122347 272778
rect 121564 272720 122286 272776
rect 122342 272720 122347 272776
rect 121564 272718 122347 272720
rect 292836 272776 295399 272778
rect 292836 272720 295338 272776
rect 295394 272720 295399 272776
rect 292836 272718 295399 272720
rect 121564 272716 121570 272718
rect 122281 272715 122347 272718
rect 295333 272715 295399 272718
rect 179462 272650 180044 272710
rect 176653 272642 176719 272645
rect 179462 272642 179522 272650
rect 176653 272640 179522 272642
rect 176653 272584 176658 272640
rect 176714 272584 179522 272640
rect 176653 272582 179522 272584
rect 176653 272579 176719 272582
rect 358077 272506 358143 272509
rect 390502 272506 390508 272508
rect 358077 272504 390508 272506
rect 358077 272448 358082 272504
rect 358138 272448 390508 272504
rect 358077 272446 390508 272448
rect 358077 272443 358143 272446
rect 390502 272444 390508 272446
rect 390572 272444 390578 272508
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 68369 272098 68435 272101
rect 121453 272098 121519 272101
rect 68369 272096 70196 272098
rect 68369 272040 68374 272096
rect 68430 272040 70196 272096
rect 68369 272038 70196 272040
rect 119876 272096 121519 272098
rect 119876 272040 121458 272096
rect 121514 272040 121519 272096
rect 583520 272084 584960 272174
rect 119876 272038 121519 272040
rect 68369 272035 68435 272038
rect 121453 272035 121519 272038
rect 67633 271418 67699 271421
rect 121453 271418 121519 271421
rect 67633 271416 70196 271418
rect 67633 271360 67638 271416
rect 67694 271360 70196 271416
rect 67633 271358 70196 271360
rect 119876 271416 121519 271418
rect 119876 271360 121458 271416
rect 121514 271360 121519 271416
rect 119876 271358 121519 271360
rect 67633 271355 67699 271358
rect 121453 271355 121519 271358
rect 571609 270874 571675 270877
rect 569940 270872 571675 270874
rect 569940 270816 571614 270872
rect 571670 270816 571675 270872
rect 569940 270814 571675 270816
rect 571609 270811 571675 270814
rect 67725 270738 67791 270741
rect 67725 270736 70196 270738
rect 67725 270680 67730 270736
rect 67786 270680 70196 270736
rect 67725 270678 70196 270680
rect 67725 270675 67791 270678
rect 179462 270610 180044 270670
rect 177757 270602 177823 270605
rect 179462 270602 179522 270610
rect 177757 270600 179522 270602
rect 177757 270544 177762 270600
rect 177818 270544 179522 270600
rect 177757 270542 179522 270544
rect 177757 270539 177823 270542
rect 67633 270058 67699 270061
rect 121545 270058 121611 270061
rect 295333 270058 295399 270061
rect 67633 270056 70196 270058
rect 67633 270000 67638 270056
rect 67694 270000 70196 270056
rect 67633 269998 70196 270000
rect 119876 270056 121611 270058
rect 119876 270000 121550 270056
rect 121606 270000 121611 270056
rect 119876 269998 121611 270000
rect 292836 270056 295399 270058
rect 292836 270000 295338 270056
rect 295394 270000 295399 270056
rect 292836 269998 295399 270000
rect 67633 269995 67699 269998
rect 121545 269995 121611 269998
rect 295333 269995 295399 269998
rect 387149 270058 387215 270061
rect 387701 270058 387767 270061
rect 387149 270056 390172 270058
rect 387149 270000 387154 270056
rect 387210 270000 387706 270056
rect 387762 270000 390172 270056
rect 387149 269998 390172 270000
rect 387149 269995 387215 269998
rect 387701 269995 387767 269998
rect 67357 269378 67423 269381
rect 121453 269378 121519 269381
rect 67357 269376 70196 269378
rect 67357 269320 67362 269376
rect 67418 269320 70196 269376
rect 67357 269318 70196 269320
rect 119876 269376 121519 269378
rect 119876 269320 121458 269376
rect 121514 269320 121519 269376
rect 119876 269318 121519 269320
rect 67357 269315 67423 269318
rect 121453 269315 121519 269318
rect 68185 268698 68251 268701
rect 120717 268698 120783 268701
rect 68185 268696 70196 268698
rect 68185 268640 68190 268696
rect 68246 268640 70196 268696
rect 68185 268638 70196 268640
rect 119876 268696 120783 268698
rect 119876 268640 120722 268696
rect 120778 268640 120783 268696
rect 119876 268638 120783 268640
rect 68185 268635 68251 268638
rect 120717 268635 120783 268638
rect 179462 268570 180044 268630
rect 176653 268562 176719 268565
rect 179462 268562 179522 268570
rect 176653 268560 179522 268562
rect 176653 268504 176658 268560
rect 176714 268504 179522 268560
rect 176653 268502 179522 268504
rect 176653 268499 176719 268502
rect 293033 268154 293099 268157
rect 292806 268152 293099 268154
rect 292806 268096 293038 268152
rect 293094 268096 293099 268152
rect 292806 268094 293099 268096
rect 67633 268018 67699 268021
rect 67633 268016 70196 268018
rect 67633 267960 67638 268016
rect 67694 267960 70196 268016
rect 67633 267958 70196 267960
rect 119876 267958 122850 268018
rect 292806 267988 292866 268094
rect 293033 268091 293099 268094
rect 67633 267955 67699 267958
rect 122790 267882 122850 267958
rect 171910 267882 171916 267884
rect 122790 267822 171916 267882
rect 171910 267820 171916 267822
rect 171980 267820 171986 267884
rect 571517 267474 571583 267477
rect 569940 267472 571583 267474
rect 569940 267416 571522 267472
rect 571578 267416 571583 267472
rect 569940 267414 571583 267416
rect 571517 267411 571583 267414
rect 68921 267338 68987 267341
rect 122097 267338 122163 267341
rect 68921 267336 70196 267338
rect -960 267202 480 267292
rect 68921 267280 68926 267336
rect 68982 267280 70196 267336
rect 68921 267278 70196 267280
rect 119876 267336 122163 267338
rect 119876 267280 122102 267336
rect 122158 267280 122163 267336
rect 119876 267278 122163 267280
rect 68921 267275 68987 267278
rect 122097 267275 122163 267278
rect 3049 267202 3115 267205
rect -960 267200 3115 267202
rect -960 267144 3054 267200
rect 3110 267144 3115 267200
rect -960 267142 3115 267144
rect -960 267052 480 267142
rect 3049 267139 3115 267142
rect 67633 266658 67699 266661
rect 121453 266658 121519 266661
rect 67633 266656 70196 266658
rect 67633 266600 67638 266656
rect 67694 266600 70196 266656
rect 67633 266598 70196 266600
rect 119876 266656 121519 266658
rect 119876 266600 121458 266656
rect 121514 266600 121519 266656
rect 119876 266598 121519 266600
rect 67633 266595 67699 266598
rect 121453 266595 121519 266598
rect 387057 266658 387123 266661
rect 387057 266656 390172 266658
rect 387057 266600 387062 266656
rect 387118 266600 390172 266656
rect 387057 266598 390172 266600
rect 387057 266595 387123 266598
rect 161974 266324 161980 266388
rect 162044 266386 162050 266388
rect 165613 266386 165679 266389
rect 162044 266384 165679 266386
rect 162044 266328 165618 266384
rect 165674 266328 165679 266384
rect 162044 266326 165679 266328
rect 162044 266324 162050 266326
rect 165613 266323 165679 266326
rect 67725 265978 67791 265981
rect 121453 265978 121519 265981
rect 67725 265976 70196 265978
rect 67725 265920 67730 265976
rect 67786 265920 70196 265976
rect 67725 265918 70196 265920
rect 119876 265976 121519 265978
rect 119876 265920 121458 265976
rect 121514 265920 121519 265976
rect 119876 265918 121519 265920
rect 67725 265915 67791 265918
rect 121453 265915 121519 265918
rect 176653 265978 176719 265981
rect 295333 265978 295399 265981
rect 176653 265976 179522 265978
rect 176653 265920 176658 265976
rect 176714 265920 179522 265976
rect 176653 265918 179522 265920
rect 292836 265976 295399 265978
rect 292836 265920 295338 265976
rect 295394 265920 295399 265976
rect 292836 265918 295399 265920
rect 176653 265915 176719 265918
rect 179462 265910 179522 265918
rect 295333 265915 295399 265918
rect 179462 265850 180044 265910
rect 67633 265298 67699 265301
rect 67633 265296 70196 265298
rect 67633 265240 67638 265296
rect 67694 265240 70196 265296
rect 67633 265238 70196 265240
rect 119876 265238 122850 265298
rect 67633 265235 67699 265238
rect 122790 265162 122850 265238
rect 169150 265162 169156 265164
rect 122790 265102 169156 265162
rect 169150 265100 169156 265102
rect 169220 265100 169226 265164
rect 67633 264618 67699 264621
rect 121545 264618 121611 264621
rect 569953 264618 570019 264621
rect 67633 264616 70196 264618
rect 67633 264560 67638 264616
rect 67694 264560 70196 264616
rect 67633 264558 70196 264560
rect 119876 264616 121611 264618
rect 119876 264560 121550 264616
rect 121606 264560 121611 264616
rect 119876 264558 121611 264560
rect 67633 264555 67699 264558
rect 121545 264555 121611 264558
rect 569910 264616 570019 264618
rect 569910 264560 569958 264616
rect 570014 264560 570019 264616
rect 569910 264555 570019 264560
rect 569910 264044 569970 264555
rect 67633 263938 67699 263941
rect 121453 263938 121519 263941
rect 294045 263938 294111 263941
rect 67633 263936 70196 263938
rect 67633 263880 67638 263936
rect 67694 263880 70196 263936
rect 67633 263878 70196 263880
rect 119876 263936 121519 263938
rect 119876 263880 121458 263936
rect 121514 263880 121519 263936
rect 119876 263878 121519 263880
rect 292836 263936 294111 263938
rect 292836 263880 294050 263936
rect 294106 263880 294111 263936
rect 292836 263878 294111 263880
rect 67633 263875 67699 263878
rect 121453 263875 121519 263878
rect 294045 263875 294111 263878
rect 179462 263810 180044 263870
rect 179321 263802 179387 263805
rect 179462 263802 179522 263810
rect 179321 263800 179522 263802
rect 179321 263744 179326 263800
rect 179382 263744 179522 263800
rect 179321 263742 179522 263744
rect 179321 263739 179387 263742
rect 59169 263668 59235 263669
rect 59118 263666 59124 263668
rect 59078 263606 59124 263666
rect 59188 263664 59235 263668
rect 59230 263608 59235 263664
rect 59118 263604 59124 263606
rect 59188 263604 59235 263608
rect 59169 263603 59235 263604
rect 67725 263258 67791 263261
rect 121453 263258 121519 263261
rect 67725 263256 70196 263258
rect 67725 263200 67730 263256
rect 67786 263200 70196 263256
rect 67725 263198 70196 263200
rect 119876 263256 121519 263258
rect 119876 263200 121458 263256
rect 121514 263200 121519 263256
rect 119876 263198 121519 263200
rect 67725 263195 67791 263198
rect 121453 263195 121519 263198
rect 386873 263258 386939 263261
rect 386873 263256 390172 263258
rect 386873 263200 386878 263256
rect 386934 263200 390172 263256
rect 386873 263198 390172 263200
rect 386873 263195 386939 263198
rect 67633 262578 67699 262581
rect 121453 262578 121519 262581
rect 67633 262576 70196 262578
rect 67633 262520 67638 262576
rect 67694 262520 70196 262576
rect 67633 262518 70196 262520
rect 119876 262576 121519 262578
rect 119876 262520 121458 262576
rect 121514 262520 121519 262576
rect 119876 262518 121519 262520
rect 67633 262515 67699 262518
rect 121453 262515 121519 262518
rect 67725 261898 67791 261901
rect 121545 261898 121611 261901
rect 67725 261896 70196 261898
rect 67725 261840 67730 261896
rect 67786 261840 70196 261896
rect 67725 261838 70196 261840
rect 119876 261896 121611 261898
rect 119876 261840 121550 261896
rect 121606 261840 121611 261896
rect 119876 261838 121611 261840
rect 67725 261835 67791 261838
rect 121545 261835 121611 261838
rect 179462 261770 180044 261830
rect 176653 261762 176719 261765
rect 179462 261762 179522 261770
rect 176653 261760 179522 261762
rect 176653 261704 176658 261760
rect 176714 261704 179522 261760
rect 176653 261702 179522 261704
rect 176653 261699 176719 261702
rect 68185 261218 68251 261221
rect 121453 261218 121519 261221
rect 295333 261218 295399 261221
rect 68185 261216 70196 261218
rect 68185 261160 68190 261216
rect 68246 261160 70196 261216
rect 68185 261158 70196 261160
rect 119876 261216 121519 261218
rect 119876 261160 121458 261216
rect 121514 261160 121519 261216
rect 119876 261158 121519 261160
rect 292836 261216 295399 261218
rect 292836 261160 295338 261216
rect 295394 261160 295399 261216
rect 292836 261158 295399 261160
rect 68185 261155 68251 261158
rect 121453 261155 121519 261158
rect 295333 261155 295399 261158
rect 572621 260674 572687 260677
rect 569940 260672 572687 260674
rect 569940 260616 572626 260672
rect 572682 260616 572687 260672
rect 569940 260614 572687 260616
rect 572621 260611 572687 260614
rect 67633 260538 67699 260541
rect 121545 260538 121611 260541
rect 67633 260536 70196 260538
rect 67633 260480 67638 260536
rect 67694 260480 70196 260536
rect 67633 260478 70196 260480
rect 119876 260536 121611 260538
rect 119876 260480 121550 260536
rect 121606 260480 121611 260536
rect 119876 260478 121611 260480
rect 67633 260475 67699 260478
rect 121545 260475 121611 260478
rect 386873 259994 386939 259997
rect 386873 259992 390172 259994
rect 386873 259936 386878 259992
rect 386934 259936 390172 259992
rect 386873 259934 390172 259936
rect 386873 259931 386939 259934
rect 67633 259858 67699 259861
rect 121453 259858 121519 259861
rect 67633 259856 70196 259858
rect 67633 259800 67638 259856
rect 67694 259800 70196 259856
rect 67633 259798 70196 259800
rect 119876 259856 121519 259858
rect 119876 259800 121458 259856
rect 121514 259800 121519 259856
rect 119876 259798 121519 259800
rect 67633 259795 67699 259798
rect 121453 259795 121519 259798
rect 179462 259730 180044 259790
rect 176653 259722 176719 259725
rect 179462 259722 179522 259730
rect 176653 259720 179522 259722
rect 176653 259664 176658 259720
rect 176714 259664 179522 259720
rect 176653 259662 179522 259664
rect 176653 259659 176719 259662
rect 67725 259178 67791 259181
rect 121545 259178 121611 259181
rect 295333 259178 295399 259181
rect 67725 259176 70196 259178
rect 67725 259120 67730 259176
rect 67786 259120 70196 259176
rect 67725 259118 70196 259120
rect 119876 259176 121611 259178
rect 119876 259120 121550 259176
rect 121606 259120 121611 259176
rect 119876 259118 121611 259120
rect 292836 259176 295399 259178
rect 292836 259120 295338 259176
rect 295394 259120 295399 259176
rect 292836 259118 295399 259120
rect 67725 259115 67791 259118
rect 121545 259115 121611 259118
rect 295333 259115 295399 259118
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect 67633 258498 67699 258501
rect 121453 258498 121519 258501
rect 67633 258496 70196 258498
rect 67633 258440 67638 258496
rect 67694 258440 70196 258496
rect 67633 258438 70196 258440
rect 119876 258496 121519 258498
rect 119876 258440 121458 258496
rect 121514 258440 121519 258496
rect 119876 258438 121519 258440
rect 67633 258435 67699 258438
rect 121453 258435 121519 258438
rect 67633 257818 67699 257821
rect 121545 257818 121611 257821
rect 67633 257816 70196 257818
rect 67633 257760 67638 257816
rect 67694 257760 70196 257816
rect 67633 257758 70196 257760
rect 119876 257816 121611 257818
rect 119876 257760 121550 257816
rect 121606 257760 121611 257816
rect 119876 257758 121611 257760
rect 67633 257755 67699 257758
rect 121545 257755 121611 257758
rect 569309 257682 569375 257685
rect 569309 257680 569418 257682
rect 569309 257624 569314 257680
rect 569370 257624 569418 257680
rect 569309 257619 569418 257624
rect 156505 257276 156571 257277
rect 120022 257212 120028 257276
rect 120092 257274 120098 257276
rect 156454 257274 156460 257276
rect 120092 257214 156460 257274
rect 156524 257272 156571 257276
rect 156566 257216 156571 257272
rect 569358 257244 569418 257619
rect 120092 257212 120098 257214
rect 156454 257212 156460 257214
rect 156524 257212 156571 257216
rect 156505 257211 156571 257212
rect 67633 257138 67699 257141
rect 121453 257138 121519 257141
rect 67633 257136 70196 257138
rect 67633 257080 67638 257136
rect 67694 257080 70196 257136
rect 67633 257078 70196 257080
rect 119876 257136 121519 257138
rect 119876 257080 121458 257136
rect 121514 257080 121519 257136
rect 119876 257078 121519 257080
rect 67633 257075 67699 257078
rect 121453 257075 121519 257078
rect 179045 257138 179111 257141
rect 295977 257138 296043 257141
rect 179045 257136 179890 257138
rect 179045 257080 179050 257136
rect 179106 257080 179890 257136
rect 179045 257078 179890 257080
rect 292836 257136 296043 257138
rect 292836 257080 295982 257136
rect 296038 257080 296043 257136
rect 292836 257078 296043 257080
rect 179045 257075 179111 257078
rect 179830 257070 179890 257078
rect 295977 257075 296043 257078
rect 179830 257010 180044 257070
rect 69197 256458 69263 256461
rect 121545 256458 121611 256461
rect 69197 256456 70196 256458
rect 69197 256400 69202 256456
rect 69258 256400 70196 256456
rect 69197 256398 70196 256400
rect 119876 256456 121611 256458
rect 119876 256400 121550 256456
rect 121606 256400 121611 256456
rect 119876 256398 121611 256400
rect 69197 256395 69263 256398
rect 121545 256395 121611 256398
rect 386873 256458 386939 256461
rect 386873 256456 390172 256458
rect 386873 256400 386878 256456
rect 386934 256400 390172 256456
rect 386873 256398 390172 256400
rect 386873 256395 386939 256398
rect 67633 255778 67699 255781
rect 121453 255778 121519 255781
rect 67633 255776 70196 255778
rect 67633 255720 67638 255776
rect 67694 255720 70196 255776
rect 67633 255718 70196 255720
rect 119876 255776 121519 255778
rect 119876 255720 121458 255776
rect 121514 255720 121519 255776
rect 119876 255718 121519 255720
rect 67633 255715 67699 255718
rect 121453 255715 121519 255718
rect 124806 255098 124812 255100
rect 70166 254554 70226 255068
rect 119876 255038 124812 255098
rect 124806 255036 124812 255038
rect 124876 255036 124882 255100
rect 295609 255098 295675 255101
rect 292836 255096 295675 255098
rect 292836 255040 295614 255096
rect 295670 255040 295675 255096
rect 292836 255038 295675 255040
rect 295609 255035 295675 255038
rect 179416 254970 180044 255030
rect 176653 254962 176719 254965
rect 179416 254962 179476 254970
rect 176653 254960 179476 254962
rect 176653 254904 176658 254960
rect 176714 254904 179476 254960
rect 176653 254902 179476 254904
rect 176653 254899 176719 254902
rect 64830 254494 70226 254554
rect -960 254146 480 254236
rect 2773 254146 2839 254149
rect -960 254144 2839 254146
rect -960 254088 2778 254144
rect 2834 254088 2839 254144
rect -960 254086 2839 254088
rect -960 253996 480 254086
rect 2773 254083 2839 254086
rect 61878 254084 61884 254148
rect 61948 254146 61954 254148
rect 64830 254146 64890 254494
rect 67725 254418 67791 254421
rect 121453 254418 121519 254421
rect 67725 254416 70196 254418
rect 67725 254360 67730 254416
rect 67786 254360 70196 254416
rect 67725 254358 70196 254360
rect 119876 254416 121519 254418
rect 119876 254360 121458 254416
rect 121514 254360 121519 254416
rect 119876 254358 121519 254360
rect 67725 254355 67791 254358
rect 121453 254355 121519 254358
rect 120574 254220 120580 254284
rect 120644 254282 120650 254284
rect 157333 254282 157399 254285
rect 120644 254280 157399 254282
rect 120644 254224 157338 254280
rect 157394 254224 157399 254280
rect 120644 254222 157399 254224
rect 120644 254220 120650 254222
rect 157333 254219 157399 254222
rect 61948 254086 64890 254146
rect 61948 254084 61954 254086
rect 571425 253874 571491 253877
rect 569940 253872 571491 253874
rect 569940 253816 571430 253872
rect 571486 253816 571491 253872
rect 569940 253814 571491 253816
rect 571425 253811 571491 253814
rect 67633 253738 67699 253741
rect 121545 253738 121611 253741
rect 67633 253736 70196 253738
rect 67633 253680 67638 253736
rect 67694 253680 70196 253736
rect 67633 253678 70196 253680
rect 119876 253736 121611 253738
rect 119876 253680 121550 253736
rect 121606 253680 121611 253736
rect 119876 253678 121611 253680
rect 67633 253675 67699 253678
rect 121545 253675 121611 253678
rect 69013 253058 69079 253061
rect 121453 253058 121519 253061
rect 69013 253056 70196 253058
rect 69013 253000 69018 253056
rect 69074 253000 70196 253056
rect 69013 252998 70196 253000
rect 119876 253056 121519 253058
rect 119876 253000 121458 253056
rect 121514 253000 121519 253056
rect 119876 252998 121519 253000
rect 69013 252995 69079 252998
rect 121453 252995 121519 252998
rect 386873 253058 386939 253061
rect 386873 253056 390172 253058
rect 386873 253000 386878 253056
rect 386934 253000 390172 253056
rect 386873 252998 390172 253000
rect 386873 252995 386939 252998
rect 179416 252930 180044 252990
rect 176469 252922 176535 252925
rect 179416 252922 179476 252930
rect 176469 252920 179476 252922
rect 176469 252864 176474 252920
rect 176530 252864 179476 252920
rect 176469 252862 179476 252864
rect 176469 252859 176535 252862
rect 68921 252378 68987 252381
rect 121545 252378 121611 252381
rect 68921 252376 70196 252378
rect 68921 252320 68926 252376
rect 68982 252320 70196 252376
rect 68921 252318 70196 252320
rect 119876 252376 121611 252378
rect 119876 252320 121550 252376
rect 121606 252320 121611 252376
rect 119876 252318 121611 252320
rect 68921 252315 68987 252318
rect 121545 252315 121611 252318
rect 292806 252106 292866 252348
rect 296529 252106 296595 252109
rect 297173 252106 297239 252109
rect 292806 252104 297239 252106
rect 292806 252048 296534 252104
rect 296590 252048 297178 252104
rect 297234 252048 297239 252104
rect 292806 252046 297239 252048
rect 296529 252043 296595 252046
rect 297173 252043 297239 252046
rect 67265 251698 67331 251701
rect 121453 251698 121519 251701
rect 67265 251696 70196 251698
rect 67265 251640 67270 251696
rect 67326 251640 70196 251696
rect 67265 251638 70196 251640
rect 119876 251696 121519 251698
rect 119876 251640 121458 251696
rect 121514 251640 121519 251696
rect 119876 251638 121519 251640
rect 67265 251635 67331 251638
rect 121453 251635 121519 251638
rect 572621 251154 572687 251157
rect 569940 251152 572687 251154
rect 569940 251096 572626 251152
rect 572682 251096 572687 251152
rect 569940 251094 572687 251096
rect 572621 251091 572687 251094
rect 67725 251018 67791 251021
rect 120165 251018 120231 251021
rect 120717 251018 120783 251021
rect 67725 251016 70196 251018
rect 67725 250960 67730 251016
rect 67786 250960 70196 251016
rect 67725 250958 70196 250960
rect 119876 251016 120783 251018
rect 119876 250960 120170 251016
rect 120226 250960 120722 251016
rect 120778 250960 120783 251016
rect 119876 250958 120783 250960
rect 67725 250955 67791 250958
rect 120165 250955 120231 250958
rect 120717 250955 120783 250958
rect 179416 250890 180044 250950
rect 177665 250882 177731 250885
rect 179416 250882 179476 250890
rect 177665 250880 179476 250882
rect 177665 250824 177670 250880
rect 177726 250824 179476 250880
rect 177665 250822 179476 250824
rect 177665 250819 177731 250822
rect 67633 250338 67699 250341
rect 121453 250338 121519 250341
rect 296621 250338 296687 250341
rect 67633 250336 70196 250338
rect 67633 250280 67638 250336
rect 67694 250280 70196 250336
rect 67633 250278 70196 250280
rect 119876 250336 121519 250338
rect 119876 250280 121458 250336
rect 121514 250280 121519 250336
rect 119876 250278 121519 250280
rect 292836 250336 296687 250338
rect 292836 250280 296626 250336
rect 296682 250280 296687 250336
rect 292836 250278 296687 250280
rect 67633 250275 67699 250278
rect 121453 250275 121519 250278
rect 296621 250275 296687 250278
rect 67633 249658 67699 249661
rect 387517 249658 387583 249661
rect 67633 249656 70196 249658
rect 67633 249600 67638 249656
rect 67694 249600 70196 249656
rect 387517 249656 390172 249658
rect 67633 249598 70196 249600
rect 67633 249595 67699 249598
rect 119846 249114 119906 249628
rect 387517 249600 387522 249656
rect 387578 249600 390172 249656
rect 387517 249598 390172 249600
rect 387517 249595 387583 249598
rect 119846 249054 122850 249114
rect 67633 248978 67699 248981
rect 121453 248978 121519 248981
rect 67633 248976 70196 248978
rect 67633 248920 67638 248976
rect 67694 248920 70196 248976
rect 67633 248918 70196 248920
rect 119876 248976 121519 248978
rect 119876 248920 121458 248976
rect 121514 248920 121519 248976
rect 119876 248918 121519 248920
rect 67633 248915 67699 248918
rect 121453 248915 121519 248918
rect 122790 248434 122850 249054
rect 142654 248434 142660 248436
rect 122790 248374 142660 248434
rect 142654 248372 142660 248374
rect 142724 248372 142730 248436
rect 296529 248434 296595 248437
rect 296662 248434 296668 248436
rect 296529 248432 296668 248434
rect 296529 248376 296534 248432
rect 296590 248376 296668 248432
rect 296529 248374 296668 248376
rect 296529 248371 296595 248374
rect 296662 248372 296668 248374
rect 296732 248372 296738 248436
rect 67725 248298 67791 248301
rect 121453 248298 121519 248301
rect 295517 248298 295583 248301
rect 67725 248296 70196 248298
rect 67725 248240 67730 248296
rect 67786 248240 70196 248296
rect 67725 248238 70196 248240
rect 119876 248296 121519 248298
rect 119876 248240 121458 248296
rect 121514 248240 121519 248296
rect 119876 248238 121519 248240
rect 292836 248296 295583 248298
rect 292836 248240 295522 248296
rect 295578 248240 295583 248296
rect 292836 248238 295583 248240
rect 67725 248235 67791 248238
rect 121453 248235 121519 248238
rect 295517 248235 295583 248238
rect 179462 248170 180044 248230
rect 179462 248165 179522 248170
rect 179413 248160 179522 248165
rect 179413 248104 179418 248160
rect 179474 248104 179522 248160
rect 179413 248102 179522 248104
rect 179413 248099 179479 248102
rect 572621 247754 572687 247757
rect 569940 247752 572687 247754
rect 569940 247696 572626 247752
rect 572682 247696 572687 247752
rect 569940 247694 572687 247696
rect 572621 247691 572687 247694
rect 67633 247618 67699 247621
rect 67633 247616 70196 247618
rect 67633 247560 67638 247616
rect 67694 247560 70196 247616
rect 67633 247558 70196 247560
rect 67633 247555 67699 247558
rect 119846 247074 119906 247588
rect 171726 247074 171732 247076
rect 119846 247014 171732 247074
rect 171726 247012 171732 247014
rect 171796 247012 171802 247076
rect 121545 246938 121611 246941
rect 119876 246936 121611 246938
rect 70166 246394 70226 246908
rect 119876 246880 121550 246936
rect 121606 246880 121611 246936
rect 119876 246878 121611 246880
rect 121545 246875 121611 246878
rect 64830 246334 70226 246394
rect 386873 246394 386939 246397
rect 386873 246392 390172 246394
rect 386873 246336 386878 246392
rect 386934 246336 390172 246392
rect 386873 246334 390172 246336
rect 63350 245788 63356 245852
rect 63420 245850 63426 245852
rect 64830 245850 64890 246334
rect 386873 246331 386939 246334
rect 67398 246196 67404 246260
rect 67468 246258 67474 246260
rect 121453 246258 121519 246261
rect 295517 246258 295583 246261
rect 67468 246198 70196 246258
rect 119876 246256 121519 246258
rect 119876 246200 121458 246256
rect 121514 246200 121519 246256
rect 119876 246198 121519 246200
rect 292836 246256 295583 246258
rect 292836 246200 295522 246256
rect 295578 246200 295583 246256
rect 292836 246198 295583 246200
rect 67468 246196 67474 246198
rect 121453 246195 121519 246198
rect 295517 246195 295583 246198
rect 179830 246130 180044 246190
rect 176653 246122 176719 246125
rect 179045 246122 179111 246125
rect 179830 246122 179890 246130
rect 176653 246120 179890 246122
rect 176653 246064 176658 246120
rect 176714 246064 179050 246120
rect 179106 246064 179890 246120
rect 176653 246062 179890 246064
rect 176653 246059 176719 246062
rect 179045 246059 179111 246062
rect 63420 245790 64890 245850
rect 63420 245788 63426 245790
rect 68093 245578 68159 245581
rect 69289 245578 69355 245581
rect 121545 245578 121611 245581
rect 68093 245576 70196 245578
rect 68093 245520 68098 245576
rect 68154 245520 69294 245576
rect 69350 245520 70196 245576
rect 68093 245518 70196 245520
rect 119876 245576 121611 245578
rect 119876 245520 121550 245576
rect 121606 245520 121611 245576
rect 119876 245518 121611 245520
rect 68093 245515 68159 245518
rect 69289 245515 69355 245518
rect 121545 245515 121611 245518
rect 582741 245578 582807 245581
rect 583520 245578 584960 245668
rect 582741 245576 584960 245578
rect 582741 245520 582746 245576
rect 582802 245520 584960 245576
rect 582741 245518 584960 245520
rect 582741 245515 582807 245518
rect 583520 245428 584960 245518
rect 68001 244898 68067 244901
rect 121453 244898 121519 244901
rect 68001 244896 70196 244898
rect 68001 244840 68006 244896
rect 68062 244840 70196 244896
rect 68001 244838 70196 244840
rect 119876 244896 121519 244898
rect 119876 244840 121458 244896
rect 121514 244840 121519 244896
rect 119876 244838 121519 244840
rect 68001 244835 68067 244838
rect 121453 244835 121519 244838
rect 160093 244898 160159 244901
rect 161289 244898 161355 244901
rect 167494 244898 167500 244900
rect 160093 244896 167500 244898
rect 160093 244840 160098 244896
rect 160154 244840 161294 244896
rect 161350 244840 167500 244896
rect 160093 244838 167500 244840
rect 160093 244835 160159 244838
rect 161289 244835 161355 244838
rect 167494 244836 167500 244838
rect 167564 244836 167570 244900
rect 571374 244354 571380 244356
rect 569940 244294 571380 244354
rect 571374 244292 571380 244294
rect 571444 244292 571450 244356
rect 67541 244218 67607 244221
rect 121545 244218 121611 244221
rect 67541 244216 70196 244218
rect 67541 244160 67546 244216
rect 67602 244160 70196 244216
rect 67541 244158 70196 244160
rect 119876 244216 121611 244218
rect 119876 244160 121550 244216
rect 121606 244160 121611 244216
rect 119876 244158 121611 244160
rect 67541 244155 67607 244158
rect 121545 244155 121611 244158
rect 179781 244150 179847 244153
rect 179781 244148 180044 244150
rect 179781 244092 179786 244148
rect 179842 244092 180044 244148
rect 179781 244090 180044 244092
rect 179781 244087 179847 244090
rect 121453 243538 121519 243541
rect 295793 243538 295859 243541
rect 119876 243536 121519 243538
rect 46197 242994 46263 242997
rect 69054 242994 69060 242996
rect 46197 242992 69060 242994
rect 46197 242936 46202 242992
rect 46258 242936 69060 242992
rect 46197 242934 69060 242936
rect 46197 242931 46263 242934
rect 69054 242932 69060 242934
rect 69124 242994 69130 242996
rect 70166 242994 70226 243508
rect 119876 243480 121458 243536
rect 121514 243480 121519 243536
rect 292652 243536 295859 243538
rect 292652 243508 295798 243536
rect 119876 243478 121519 243480
rect 121453 243475 121519 243478
rect 292622 243480 295798 243508
rect 295854 243480 295859 243536
rect 292622 243478 295859 243480
rect 69124 242934 70226 242994
rect 179505 242994 179571 242997
rect 292622 242996 292682 243478
rect 295793 243475 295859 243478
rect 386597 243538 386663 243541
rect 386597 243536 390172 243538
rect 386597 243480 386602 243536
rect 386658 243480 390172 243536
rect 386597 243478 390172 243480
rect 386597 243475 386663 243478
rect 179822 242994 179828 242996
rect 179505 242992 179828 242994
rect 179505 242936 179510 242992
rect 179566 242936 179828 242992
rect 179505 242934 179828 242936
rect 69124 242932 69130 242934
rect 179505 242931 179571 242934
rect 179822 242932 179828 242934
rect 179892 242932 179898 242996
rect 292614 242932 292620 242996
rect 292684 242932 292690 242996
rect 121453 242858 121519 242861
rect 119876 242856 121519 242858
rect 70166 242314 70226 242828
rect 119876 242800 121458 242856
rect 121514 242800 121519 242856
rect 119876 242798 121519 242800
rect 121453 242795 121519 242798
rect 120022 242524 120028 242588
rect 120092 242586 120098 242588
rect 124121 242586 124187 242589
rect 120092 242584 124187 242586
rect 120092 242528 124126 242584
rect 124182 242528 124187 242584
rect 120092 242526 124187 242528
rect 120092 242524 120098 242526
rect 124121 242523 124187 242526
rect 64830 242254 70226 242314
rect 63166 241708 63172 241772
rect 63236 241770 63242 241772
rect 64830 241770 64890 242254
rect 67633 242178 67699 242181
rect 121637 242178 121703 242181
rect 67633 242176 70196 242178
rect 67633 242120 67638 242176
rect 67694 242120 70196 242176
rect 67633 242118 70196 242120
rect 119876 242176 121703 242178
rect 119876 242120 121642 242176
rect 121698 242120 121703 242176
rect 119876 242118 121703 242120
rect 67633 242115 67699 242118
rect 121637 242115 121703 242118
rect 126094 242116 126100 242180
rect 126164 242178 126170 242180
rect 168373 242178 168439 242181
rect 126164 242176 168439 242178
rect 126164 242120 168378 242176
rect 168434 242120 168439 242176
rect 126164 242118 168439 242120
rect 126164 242116 126170 242118
rect 168373 242115 168439 242118
rect 179462 242050 180044 242110
rect 177573 242042 177639 242045
rect 179462 242042 179522 242050
rect 177573 242040 179522 242042
rect 177573 241984 177578 242040
rect 177634 241984 179522 242040
rect 177573 241982 179522 241984
rect 177573 241979 177639 241982
rect 63236 241710 64890 241770
rect 63236 241708 63242 241710
rect 66110 241436 66116 241500
rect 66180 241498 66186 241500
rect 120073 241498 120139 241501
rect 293309 241498 293375 241501
rect 66180 241438 70196 241498
rect 119876 241496 120139 241498
rect 119876 241440 120078 241496
rect 120134 241440 120139 241496
rect 119876 241438 120139 241440
rect 292836 241496 293375 241498
rect 292836 241440 293314 241496
rect 293370 241440 293375 241496
rect 292836 241438 293375 241440
rect 66180 241436 66186 241438
rect 120073 241435 120139 241438
rect 293309 241435 293375 241438
rect 368473 241498 368539 241501
rect 369301 241498 369367 241501
rect 368473 241496 369367 241498
rect 368473 241440 368478 241496
rect 368534 241440 369306 241496
rect 369362 241440 369367 241496
rect 368473 241438 369367 241440
rect 368473 241435 368539 241438
rect 369301 241435 369367 241438
rect 165061 241226 165127 241229
rect 368473 241226 368539 241229
rect 165061 241224 368539 241226
rect -960 241090 480 241180
rect 165061 241168 165066 241224
rect 165122 241168 368478 241224
rect 368534 241168 368539 241224
rect 165061 241166 368539 241168
rect 165061 241163 165127 241166
rect 368473 241163 368539 241166
rect 3417 241090 3483 241093
rect -960 241088 3483 241090
rect -960 241032 3422 241088
rect 3478 241032 3483 241088
rect -960 241030 3483 241032
rect -960 240940 480 241030
rect 3417 241027 3483 241030
rect 572621 240954 572687 240957
rect 569940 240952 572687 240954
rect 569940 240896 572626 240952
rect 572682 240896 572687 240952
rect 569940 240894 572687 240896
rect 572621 240891 572687 240894
rect 121453 240818 121519 240821
rect 119876 240816 121519 240818
rect 70534 240276 70594 240788
rect 119876 240760 121458 240816
rect 121514 240760 121519 240816
rect 119876 240758 121519 240760
rect 121453 240755 121519 240758
rect 123569 240818 123635 240821
rect 299473 240818 299539 240821
rect 123569 240816 200130 240818
rect 123569 240760 123574 240816
rect 123630 240760 200130 240816
rect 123569 240758 200130 240760
rect 123569 240755 123635 240758
rect 200070 240682 200130 240758
rect 277350 240816 299539 240818
rect 277350 240760 299478 240816
rect 299534 240760 299539 240816
rect 277350 240758 299539 240760
rect 204253 240682 204319 240685
rect 200070 240680 204319 240682
rect 200070 240624 204258 240680
rect 204314 240624 204319 240680
rect 200070 240622 204319 240624
rect 204253 240619 204319 240622
rect 276289 240682 276355 240685
rect 277350 240682 277410 240758
rect 299473 240755 299539 240758
rect 276289 240680 277410 240682
rect 276289 240624 276294 240680
rect 276350 240624 277410 240680
rect 276289 240622 277410 240624
rect 276289 240619 276355 240622
rect 70526 240212 70532 240276
rect 70596 240212 70602 240276
rect 386873 240274 386939 240277
rect 386873 240272 390172 240274
rect 386873 240216 386878 240272
rect 386934 240216 390172 240272
rect 386873 240214 390172 240216
rect 386873 240211 386939 240214
rect 61837 240140 61903 240141
rect 61837 240136 61884 240140
rect 61948 240138 61954 240140
rect 121545 240138 121611 240141
rect 61837 240080 61842 240136
rect 61837 240076 61884 240080
rect 61948 240078 61994 240138
rect 119876 240136 121611 240138
rect 119876 240080 121550 240136
rect 121606 240080 121611 240136
rect 119876 240078 121611 240080
rect 61948 240076 61954 240078
rect 61837 240075 61903 240076
rect 121545 240075 121611 240078
rect 288934 240076 288940 240140
rect 289004 240138 289010 240140
rect 294086 240138 294092 240140
rect 289004 240078 294092 240138
rect 289004 240076 289010 240078
rect 294086 240076 294092 240078
rect 294156 240076 294162 240140
rect 57605 239866 57671 239869
rect 313273 239866 313339 239869
rect 57605 239864 313339 239866
rect 57605 239808 57610 239864
rect 57666 239808 313278 239864
rect 313334 239808 313339 239864
rect 57605 239806 313339 239808
rect 57605 239803 57671 239806
rect 313273 239803 313339 239806
rect 117037 239730 117103 239733
rect 120574 239730 120580 239732
rect 117037 239728 120580 239730
rect 117037 239672 117042 239728
rect 117098 239672 120580 239728
rect 117037 239670 120580 239672
rect 117037 239667 117103 239670
rect 120574 239668 120580 239670
rect 120644 239668 120650 239732
rect 35157 239458 35223 239461
rect 35801 239458 35867 239461
rect 161974 239458 161980 239460
rect 35157 239456 161980 239458
rect 35157 239400 35162 239456
rect 35218 239400 35806 239456
rect 35862 239400 161980 239456
rect 35157 239398 161980 239400
rect 35157 239395 35223 239398
rect 35801 239395 35867 239398
rect 161974 239396 161980 239398
rect 162044 239396 162050 239460
rect 178534 239396 178540 239460
rect 178604 239458 178610 239460
rect 215201 239458 215267 239461
rect 178604 239456 215267 239458
rect 178604 239400 215206 239456
rect 215262 239400 215267 239456
rect 178604 239398 215267 239400
rect 178604 239396 178610 239398
rect 215201 239395 215267 239398
rect 287697 238914 287763 238917
rect 287697 238912 288082 238914
rect 287697 238856 287702 238912
rect 287758 238856 288082 238912
rect 287697 238854 288082 238856
rect 287697 238851 287763 238854
rect 149646 238716 149652 238780
rect 149716 238778 149722 238780
rect 287881 238778 287947 238781
rect 149716 238776 287947 238778
rect 149716 238720 287886 238776
rect 287942 238720 287947 238776
rect 149716 238718 287947 238720
rect 288022 238778 288082 238854
rect 291101 238778 291167 238781
rect 389766 238778 389772 238780
rect 288022 238776 389772 238778
rect 288022 238720 291106 238776
rect 291162 238720 389772 238776
rect 288022 238718 389772 238720
rect 149716 238716 149722 238718
rect 287881 238715 287947 238718
rect 291101 238715 291167 238718
rect 389766 238716 389772 238718
rect 389836 238716 389842 238780
rect 118969 238642 119035 238645
rect 119838 238642 119844 238644
rect 118969 238640 119844 238642
rect 118969 238584 118974 238640
rect 119030 238584 119844 238640
rect 118969 238582 119844 238584
rect 118969 238579 119035 238582
rect 119838 238580 119844 238582
rect 119908 238580 119914 238644
rect 240501 238642 240567 238645
rect 371969 238642 372035 238645
rect 240501 238640 372035 238642
rect 240501 238584 240506 238640
rect 240562 238584 371974 238640
rect 372030 238584 372035 238640
rect 240501 238582 372035 238584
rect 240501 238579 240567 238582
rect 371969 238579 372035 238582
rect 115105 238506 115171 238509
rect 236269 238506 236335 238509
rect 115105 238504 236335 238506
rect 115105 238448 115110 238504
rect 115166 238448 236274 238504
rect 236330 238448 236335 238504
rect 115105 238446 236335 238448
rect 115105 238443 115171 238446
rect 236269 238443 236335 238446
rect 254669 238506 254735 238509
rect 293166 238506 293172 238508
rect 254669 238504 293172 238506
rect 254669 238448 254674 238504
rect 254730 238448 293172 238504
rect 254669 238446 293172 238448
rect 254669 238443 254735 238446
rect 293166 238444 293172 238446
rect 293236 238444 293242 238508
rect 106733 238370 106799 238373
rect 119654 238370 119660 238372
rect 106733 238368 119660 238370
rect 106733 238312 106738 238368
rect 106794 238312 119660 238368
rect 106733 238310 119660 238312
rect 106733 238307 106799 238310
rect 119654 238308 119660 238310
rect 119724 238308 119730 238372
rect 98361 238234 98427 238237
rect 233877 238234 233943 238237
rect 98361 238232 233943 238234
rect 98361 238176 98366 238232
rect 98422 238176 233882 238232
rect 233938 238176 233943 238232
rect 98361 238174 233943 238176
rect 98361 238171 98427 238174
rect 233877 238171 233943 238174
rect 207381 237418 207447 237421
rect 208158 237418 208164 237420
rect 207381 237416 208164 237418
rect 207381 237360 207386 237416
rect 207442 237360 208164 237416
rect 207381 237358 208164 237360
rect 207381 237355 207447 237358
rect 208158 237356 208164 237358
rect 208228 237356 208234 237420
rect 569910 237285 569970 237388
rect 157241 237282 157307 237285
rect 380341 237282 380407 237285
rect 157241 237280 380407 237282
rect 157241 237224 157246 237280
rect 157302 237224 380346 237280
rect 380402 237224 380407 237280
rect 157241 237222 380407 237224
rect 569910 237280 570019 237285
rect 569910 237224 569958 237280
rect 570014 237224 570019 237280
rect 569910 237222 570019 237224
rect 157241 237219 157307 237222
rect 380341 237219 380407 237222
rect 569953 237219 570019 237222
rect 117221 237146 117287 237149
rect 192201 237146 192267 237149
rect 370589 237146 370655 237149
rect 117221 237144 370655 237146
rect 117221 237088 117226 237144
rect 117282 237088 192206 237144
rect 192262 237088 370594 237144
rect 370650 237088 370655 237144
rect 117221 237086 370655 237088
rect 117221 237083 117287 237086
rect 192201 237083 192267 237086
rect 370589 237083 370655 237086
rect 386781 236738 386847 236741
rect 386781 236736 390172 236738
rect 386781 236680 386786 236736
rect 386842 236680 390172 236736
rect 386781 236678 390172 236680
rect 386781 236675 386847 236678
rect 167678 235860 167684 235924
rect 167748 235922 167754 235924
rect 383101 235922 383167 235925
rect 167748 235920 383167 235922
rect 167748 235864 383106 235920
rect 383162 235864 383167 235920
rect 167748 235862 383167 235864
rect 167748 235860 167754 235862
rect 383101 235859 383167 235862
rect 146886 235180 146892 235244
rect 146956 235242 146962 235244
rect 202137 235242 202203 235245
rect 146956 235240 202203 235242
rect 146956 235184 202142 235240
rect 202198 235184 202203 235240
rect 146956 235182 202203 235184
rect 146956 235180 146962 235182
rect 202137 235179 202203 235182
rect 382273 234698 382339 234701
rect 383101 234698 383167 234701
rect 382273 234696 383167 234698
rect 382273 234640 382278 234696
rect 382334 234640 383106 234696
rect 383162 234640 383167 234696
rect 382273 234638 383167 234640
rect 382273 234635 382339 234638
rect 383101 234635 383167 234638
rect 161238 234500 161244 234564
rect 161308 234562 161314 234564
rect 359549 234562 359615 234565
rect 161308 234560 359615 234562
rect 161308 234504 359554 234560
rect 359610 234504 359615 234560
rect 161308 234502 359615 234504
rect 161308 234500 161314 234502
rect 359549 234499 359615 234502
rect 180885 234426 180951 234429
rect 296478 234426 296484 234428
rect 180885 234424 296484 234426
rect 180885 234368 180890 234424
rect 180946 234368 296484 234424
rect 180885 234366 296484 234368
rect 180885 234363 180951 234366
rect 296478 234364 296484 234366
rect 296548 234364 296554 234428
rect 572621 234154 572687 234157
rect 569940 234152 572687 234154
rect 569940 234096 572626 234152
rect 572682 234096 572687 234152
rect 569940 234094 572687 234096
rect 572621 234091 572687 234094
rect 386505 233474 386571 233477
rect 386505 233472 390172 233474
rect 386505 233416 386510 233472
rect 386566 233416 390172 233472
rect 386505 233414 390172 233416
rect 386505 233411 386571 233414
rect 166206 233140 166212 233204
rect 166276 233202 166282 233204
rect 306465 233202 306531 233205
rect 166276 233200 306531 233202
rect 166276 233144 306470 233200
rect 306526 233144 306531 233200
rect 166276 233142 306531 233144
rect 166276 233140 166282 233142
rect 306465 233139 306531 233142
rect 158478 232596 158484 232660
rect 158548 232658 158554 232660
rect 206277 232658 206343 232661
rect 158548 232656 206343 232658
rect 158548 232600 206282 232656
rect 206338 232600 206343 232656
rect 158548 232598 206343 232600
rect 158548 232596 158554 232598
rect 206277 232595 206343 232598
rect 122097 232522 122163 232525
rect 322054 232522 322060 232524
rect 122097 232520 322060 232522
rect 122097 232464 122102 232520
rect 122158 232464 322060 232520
rect 122097 232462 322060 232464
rect 122097 232459 122163 232462
rect 322054 232460 322060 232462
rect 322124 232460 322130 232524
rect 583385 232386 583451 232389
rect 583520 232386 584960 232476
rect 583385 232384 584960 232386
rect 583385 232328 583390 232384
rect 583446 232328 584960 232384
rect 583385 232326 584960 232328
rect 583385 232323 583451 232326
rect 583520 232236 584960 232326
rect 159449 231842 159515 231845
rect 300945 231842 301011 231845
rect 159449 231840 301011 231842
rect 159449 231784 159454 231840
rect 159510 231784 300950 231840
rect 301006 231784 301011 231840
rect 159449 231782 301011 231784
rect 159449 231779 159515 231782
rect 300945 231779 301011 231782
rect 572621 230754 572687 230757
rect 569940 230752 572687 230754
rect 569940 230696 572626 230752
rect 572682 230696 572687 230752
rect 569940 230694 572687 230696
rect 572621 230691 572687 230694
rect 75821 230482 75887 230485
rect 292614 230482 292620 230484
rect 75821 230480 292620 230482
rect 75821 230424 75826 230480
rect 75882 230424 292620 230480
rect 75821 230422 292620 230424
rect 75821 230419 75887 230422
rect 292614 230420 292620 230422
rect 292684 230420 292690 230484
rect 387149 230074 387215 230077
rect 387149 230072 390172 230074
rect 387149 230016 387154 230072
rect 387210 230016 390172 230072
rect 387149 230014 390172 230016
rect 387149 230011 387215 230014
rect 59118 229740 59124 229804
rect 59188 229802 59194 229804
rect 162301 229802 162367 229805
rect 59188 229800 162367 229802
rect 59188 229744 162306 229800
rect 162362 229744 162367 229800
rect 59188 229742 162367 229744
rect 59188 229740 59194 229742
rect 162301 229739 162367 229742
rect 63166 228924 63172 228988
rect 63236 228986 63242 228988
rect 265617 228986 265683 228989
rect 63236 228984 265683 228986
rect 63236 228928 265622 228984
rect 265678 228928 265683 228984
rect 63236 228926 265683 228928
rect 63236 228924 63242 228926
rect 265617 228923 265683 228926
rect 161974 228788 161980 228852
rect 162044 228850 162050 228852
rect 356789 228850 356855 228853
rect 162044 228848 356855 228850
rect 162044 228792 356794 228848
rect 356850 228792 356855 228848
rect 162044 228790 356855 228792
rect 162044 228788 162050 228790
rect 356789 228787 356855 228790
rect -960 227884 480 228124
rect 265617 227764 265683 227765
rect 265566 227700 265572 227764
rect 265636 227762 265683 227764
rect 265636 227760 265728 227762
rect 265678 227704 265728 227760
rect 265636 227702 265728 227704
rect 265636 227700 265683 227702
rect 265617 227699 265683 227700
rect 145649 227626 145715 227629
rect 347681 227626 347747 227629
rect 145649 227624 347747 227626
rect 145649 227568 145654 227624
rect 145710 227568 347686 227624
rect 347742 227568 347747 227624
rect 145649 227566 347747 227568
rect 145649 227563 145715 227566
rect 347681 227563 347747 227566
rect 572621 227354 572687 227357
rect 569940 227352 572687 227354
rect 569940 227296 572626 227352
rect 572682 227296 572687 227352
rect 569940 227294 572687 227296
rect 572621 227291 572687 227294
rect 386413 226674 386479 226677
rect 386413 226672 390172 226674
rect 386413 226616 386418 226672
rect 386474 226616 390172 226672
rect 386413 226614 390172 226616
rect 386413 226611 386479 226614
rect 147213 226266 147279 226269
rect 291694 226266 291700 226268
rect 147213 226264 291700 226266
rect 147213 226208 147218 226264
rect 147274 226208 291700 226264
rect 147213 226206 291700 226208
rect 147213 226203 147279 226206
rect 291694 226204 291700 226206
rect 291764 226204 291770 226268
rect 70894 224844 70900 224908
rect 70964 224906 70970 224908
rect 373993 224906 374059 224909
rect 374729 224906 374795 224909
rect 70964 224904 374795 224906
rect 70964 224848 373998 224904
rect 374054 224848 374734 224904
rect 374790 224848 374795 224904
rect 70964 224846 374795 224848
rect 70964 224844 70970 224846
rect 373993 224843 374059 224846
rect 374729 224843 374795 224846
rect 63350 224708 63356 224772
rect 63420 224770 63426 224772
rect 301037 224770 301103 224773
rect 63420 224768 301103 224770
rect 63420 224712 301042 224768
rect 301098 224712 301103 224768
rect 63420 224710 301103 224712
rect 63420 224708 63426 224710
rect 301037 224707 301103 224710
rect 179045 224634 179111 224637
rect 387006 224634 387012 224636
rect 179045 224632 387012 224634
rect 179045 224576 179050 224632
rect 179106 224576 387012 224632
rect 179045 224574 387012 224576
rect 179045 224571 179111 224574
rect 387006 224572 387012 224574
rect 387076 224572 387082 224636
rect 570137 223954 570203 223957
rect 569940 223952 570203 223954
rect 569940 223896 570142 223952
rect 570198 223896 570203 223952
rect 569940 223894 570203 223896
rect 570137 223891 570203 223894
rect 386965 223274 387031 223277
rect 387149 223274 387215 223277
rect 386965 223272 390172 223274
rect 386965 223216 386970 223272
rect 387026 223216 387154 223272
rect 387210 223216 390172 223272
rect 386965 223214 390172 223216
rect 386965 223211 387031 223214
rect 387149 223211 387215 223214
rect 64638 222804 64644 222868
rect 64708 222866 64714 222868
rect 353293 222866 353359 222869
rect 64708 222864 353359 222866
rect 64708 222808 353298 222864
rect 353354 222808 353359 222864
rect 64708 222806 353359 222808
rect 64708 222804 64714 222806
rect 353293 222803 353359 222806
rect 387057 222186 387123 222189
rect 388294 222186 388300 222188
rect 387057 222184 388300 222186
rect 387057 222128 387062 222184
rect 387118 222128 388300 222184
rect 387057 222126 388300 222128
rect 387057 222123 387123 222126
rect 388294 222124 388300 222126
rect 388364 222124 388370 222188
rect 569309 220826 569375 220829
rect 569309 220824 569418 220826
rect 569309 220768 569314 220824
rect 569370 220768 569418 220824
rect 569309 220763 569418 220768
rect 569358 220524 569418 220763
rect 386873 219874 386939 219877
rect 386873 219872 390172 219874
rect 386873 219816 386878 219872
rect 386934 219816 390172 219872
rect 386873 219814 390172 219816
rect 386873 219811 386939 219814
rect 580073 219058 580139 219061
rect 583520 219058 584960 219148
rect 580073 219056 584960 219058
rect 580073 219000 580078 219056
rect 580134 219000 584960 219056
rect 580073 218998 584960 219000
rect 580073 218995 580139 218998
rect 583520 218908 584960 218998
rect 61929 218650 61995 218653
rect 255262 218650 255268 218652
rect 61929 218648 255268 218650
rect 61929 218592 61934 218648
rect 61990 218592 255268 218648
rect 61929 218590 255268 218592
rect 61929 218587 61995 218590
rect 255262 218588 255268 218590
rect 255332 218588 255338 218652
rect 570229 217154 570295 217157
rect 569940 217152 570295 217154
rect 569940 217096 570234 217152
rect 570290 217096 570295 217152
rect 569940 217094 570295 217096
rect 570229 217091 570295 217094
rect 142654 216548 142660 216612
rect 142724 216610 142730 216612
rect 310605 216610 310671 216613
rect 142724 216608 310671 216610
rect 142724 216552 310610 216608
rect 310666 216552 310671 216608
rect 142724 216550 310671 216552
rect 142724 216548 142730 216550
rect 310605 216547 310671 216550
rect 387517 216474 387583 216477
rect 388989 216474 389055 216477
rect 387517 216472 390172 216474
rect 387517 216416 387522 216472
rect 387578 216416 388994 216472
rect 389050 216416 390172 216472
rect 387517 216414 390172 216416
rect 387517 216411 387583 216414
rect 388989 216411 389055 216414
rect 310605 215386 310671 215389
rect 311249 215386 311315 215389
rect 310605 215384 311315 215386
rect 310605 215328 310610 215384
rect 310666 215328 311254 215384
rect 311310 215328 311315 215384
rect 310605 215326 311315 215328
rect 310605 215323 310671 215326
rect 311249 215323 311315 215326
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 161289 213890 161355 213893
rect 388437 213892 388503 213893
rect 388437 213890 388484 213892
rect 161289 213888 388484 213890
rect 161289 213832 161294 213888
rect 161350 213832 388442 213888
rect 161289 213830 388484 213832
rect 161289 213827 161355 213830
rect 388437 213828 388484 213830
rect 388548 213828 388554 213892
rect 388437 213827 388503 213828
rect 572621 213618 572687 213621
rect 569940 213616 572687 213618
rect 569940 213560 572626 213616
rect 572682 213560 572687 213616
rect 569940 213558 572687 213560
rect 572621 213555 572687 213558
rect 386873 212938 386939 212941
rect 386873 212936 390172 212938
rect 386873 212880 386878 212936
rect 386934 212880 390172 212936
rect 386873 212878 390172 212880
rect 386873 212875 386939 212878
rect 171910 211788 171916 211852
rect 171980 211850 171986 211852
rect 338113 211850 338179 211853
rect 171980 211848 338179 211850
rect 171980 211792 338118 211848
rect 338174 211792 338179 211848
rect 171980 211790 338179 211792
rect 171980 211788 171986 211790
rect 338113 211787 338179 211790
rect 572621 210354 572687 210357
rect 569940 210352 572687 210354
rect 569940 210296 572626 210352
rect 572682 210296 572687 210352
rect 569940 210294 572687 210296
rect 572621 210291 572687 210294
rect 386873 209538 386939 209541
rect 386873 209536 390172 209538
rect 386873 209480 386878 209536
rect 386934 209480 390172 209536
rect 386873 209478 390172 209480
rect 386873 209475 386939 209478
rect 67398 207572 67404 207636
rect 67468 207634 67474 207636
rect 342437 207634 342503 207637
rect 67468 207632 342503 207634
rect 67468 207576 342442 207632
rect 342498 207576 342503 207632
rect 67468 207574 342503 207576
rect 67468 207572 67474 207574
rect 342437 207571 342503 207574
rect 572437 206954 572503 206957
rect 569940 206952 572503 206954
rect 569940 206896 572442 206952
rect 572498 206896 572503 206952
rect 569940 206894 572503 206896
rect 572437 206891 572503 206894
rect 386873 206138 386939 206141
rect 386873 206136 390172 206138
rect 386873 206080 386878 206136
rect 386934 206080 390172 206136
rect 386873 206078 390172 206080
rect 386873 206075 386939 206078
rect 580901 205730 580967 205733
rect 583109 205730 583175 205733
rect 583520 205730 584960 205820
rect 580901 205728 584960 205730
rect 580901 205672 580906 205728
rect 580962 205672 583114 205728
rect 583170 205672 584960 205728
rect 580901 205670 584960 205672
rect 580901 205667 580967 205670
rect 583109 205667 583175 205670
rect 583520 205580 584960 205670
rect 131757 204914 131823 204917
rect 263542 204914 263548 204916
rect 131757 204912 263548 204914
rect 131757 204856 131762 204912
rect 131818 204856 263548 204912
rect 131757 204854 263548 204856
rect 131757 204851 131823 204854
rect 263542 204852 263548 204854
rect 263612 204852 263618 204916
rect 54937 203554 55003 203557
rect 256734 203554 256740 203556
rect 54937 203552 256740 203554
rect 54937 203496 54942 203552
rect 54998 203496 256740 203552
rect 54937 203494 256740 203496
rect 54937 203491 55003 203494
rect 256734 203492 256740 203494
rect 256804 203492 256810 203556
rect 571517 203554 571583 203557
rect 569940 203552 571583 203554
rect 569940 203496 571522 203552
rect 571578 203496 571583 203552
rect 569940 203494 571583 203496
rect 571517 203491 571583 203494
rect 386873 202738 386939 202741
rect 386873 202736 390172 202738
rect 386873 202680 386878 202736
rect 386934 202680 390172 202736
rect 386873 202678 390172 202680
rect 386873 202675 386939 202678
rect -960 201922 480 202012
rect 3417 201922 3483 201925
rect -960 201920 3483 201922
rect -960 201864 3422 201920
rect 3478 201864 3483 201920
rect -960 201862 3483 201864
rect -960 201772 480 201862
rect 3417 201859 3483 201862
rect 156454 200772 156460 200836
rect 156524 200834 156530 200836
rect 373349 200834 373415 200837
rect 571558 200834 571564 200836
rect 156524 200832 373415 200834
rect 156524 200776 373354 200832
rect 373410 200776 373415 200832
rect 156524 200774 373415 200776
rect 569940 200774 571564 200834
rect 156524 200772 156530 200774
rect 373349 200771 373415 200774
rect 571558 200772 571564 200774
rect 571628 200772 571634 200836
rect 124806 200636 124812 200700
rect 124876 200698 124882 200700
rect 349245 200698 349311 200701
rect 124876 200696 349311 200698
rect 124876 200640 349250 200696
rect 349306 200640 349311 200696
rect 124876 200638 349311 200640
rect 124876 200636 124882 200638
rect 349245 200635 349311 200638
rect 387057 199338 387123 199341
rect 387057 199336 390172 199338
rect 387057 199280 387062 199336
rect 387118 199280 390172 199336
rect 387057 199278 390172 199280
rect 387057 199275 387123 199278
rect 572621 197434 572687 197437
rect 569940 197432 572687 197434
rect 569940 197376 572626 197432
rect 572682 197376 572687 197432
rect 569940 197374 572687 197376
rect 572621 197371 572687 197374
rect 386873 196074 386939 196077
rect 386873 196072 390172 196074
rect 386873 196016 386878 196072
rect 386934 196016 390172 196072
rect 386873 196014 390172 196016
rect 386873 196011 386939 196014
rect 59261 195258 59327 195261
rect 269062 195258 269068 195260
rect 59261 195256 269068 195258
rect 59261 195200 59266 195256
rect 59322 195200 269068 195256
rect 59261 195198 269068 195200
rect 59261 195195 59327 195198
rect 269062 195196 269068 195198
rect 269132 195196 269138 195260
rect 319437 195258 319503 195261
rect 337326 195258 337332 195260
rect 319437 195256 337332 195258
rect 319437 195200 319442 195256
rect 319498 195200 337332 195256
rect 319437 195198 337332 195200
rect 319437 195195 319503 195198
rect 337326 195196 337332 195198
rect 337396 195196 337402 195260
rect 275134 193836 275140 193900
rect 275204 193898 275210 193900
rect 303613 193898 303679 193901
rect 571558 193898 571564 193900
rect 275204 193896 303679 193898
rect 275204 193840 303618 193896
rect 303674 193840 303679 193896
rect 275204 193838 303679 193840
rect 569940 193838 571564 193898
rect 275204 193836 275210 193838
rect 303613 193835 303679 193838
rect 571558 193836 571564 193838
rect 571628 193836 571634 193900
rect 386413 193354 386479 193357
rect 386413 193352 390172 193354
rect 386413 193296 386418 193352
rect 386474 193296 390172 193352
rect 386413 193294 390172 193296
rect 386413 193291 386479 193294
rect 583845 193082 583911 193085
rect 583526 193080 583911 193082
rect 583526 193024 583850 193080
rect 583906 193024 583911 193080
rect 583526 193022 583911 193024
rect 583526 192674 583586 193022
rect 583845 193019 583911 193022
rect 583342 192628 583586 192674
rect 583342 192614 584960 192628
rect 580349 192538 580415 192541
rect 583342 192538 583402 192614
rect 583520 192538 584960 192614
rect 580349 192536 584960 192538
rect 580349 192480 580354 192536
rect 580410 192480 584960 192536
rect 580349 192478 584960 192480
rect 580349 192475 580415 192478
rect 583520 192388 584960 192478
rect 197997 191178 198063 191181
rect 266302 191178 266308 191180
rect 197997 191176 266308 191178
rect 197997 191120 198002 191176
rect 198058 191120 266308 191176
rect 197997 191118 266308 191120
rect 197997 191115 198063 191118
rect 266302 191116 266308 191118
rect 266372 191116 266378 191180
rect 133137 191042 133203 191045
rect 256918 191042 256924 191044
rect 133137 191040 256924 191042
rect 133137 190984 133142 191040
rect 133198 190984 256924 191040
rect 133137 190982 256924 190984
rect 133137 190979 133203 190982
rect 256918 190980 256924 190982
rect 256988 190980 256994 191044
rect 571701 190634 571767 190637
rect 569940 190632 571767 190634
rect 569940 190576 571706 190632
rect 571762 190576 571767 190632
rect 569940 190574 571767 190576
rect 571701 190571 571767 190574
rect 229093 189818 229159 189821
rect 264094 189818 264100 189820
rect 229093 189816 264100 189818
rect 229093 189760 229098 189816
rect 229154 189760 264100 189816
rect 229093 189758 264100 189760
rect 229093 189755 229159 189758
rect 264094 189756 264100 189758
rect 264164 189756 264170 189820
rect 386873 189818 386939 189821
rect 386873 189816 390172 189818
rect 386873 189760 386878 189816
rect 386934 189760 390172 189816
rect 386873 189758 390172 189760
rect 386873 189755 386939 189758
rect 164969 189682 165035 189685
rect 254526 189682 254532 189684
rect 164969 189680 254532 189682
rect 164969 189624 164974 189680
rect 165030 189624 254532 189680
rect 164969 189622 254532 189624
rect 164969 189619 165035 189622
rect 254526 189620 254532 189622
rect 254596 189620 254602 189684
rect 324262 189076 324268 189140
rect 324332 189138 324338 189140
rect 324405 189138 324471 189141
rect 324332 189136 324471 189138
rect 324332 189080 324410 189136
rect 324466 189080 324471 189136
rect 324332 189078 324471 189080
rect 324332 189076 324338 189078
rect 324405 189075 324471 189078
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 67449 188458 67515 188461
rect 252502 188458 252508 188460
rect 67449 188456 252508 188458
rect 67449 188400 67454 188456
rect 67510 188400 252508 188456
rect 67449 188398 252508 188400
rect 67449 188395 67515 188398
rect 252502 188396 252508 188398
rect 252572 188396 252578 188460
rect 59169 188322 59235 188325
rect 259494 188322 259500 188324
rect 59169 188320 259500 188322
rect 59169 188264 59174 188320
rect 59230 188264 259500 188320
rect 59169 188262 259500 188264
rect 59169 188259 59235 188262
rect 259494 188260 259500 188262
rect 259564 188260 259570 188324
rect 186957 187234 187023 187237
rect 326654 187234 326660 187236
rect 186957 187232 326660 187234
rect 186957 187176 186962 187232
rect 187018 187176 326660 187232
rect 186957 187174 326660 187176
rect 186957 187171 187023 187174
rect 326654 187172 326660 187174
rect 326724 187172 326730 187236
rect 572621 187234 572687 187237
rect 569940 187232 572687 187234
rect 569940 187176 572626 187232
rect 572682 187176 572687 187232
rect 569940 187174 572687 187176
rect 572621 187171 572687 187174
rect 50981 187098 51047 187101
rect 265014 187098 265020 187100
rect 50981 187096 265020 187098
rect 50981 187040 50986 187096
rect 51042 187040 265020 187096
rect 50981 187038 265020 187040
rect 50981 187035 51047 187038
rect 265014 187036 265020 187038
rect 265084 187036 265090 187100
rect 73153 186962 73219 186965
rect 320214 186962 320220 186964
rect 73153 186960 320220 186962
rect 73153 186904 73158 186960
rect 73214 186904 320220 186960
rect 73153 186902 320220 186904
rect 73153 186899 73219 186902
rect 320214 186900 320220 186902
rect 320284 186900 320290 186964
rect 386781 186554 386847 186557
rect 386781 186552 390172 186554
rect 386781 186496 386786 186552
rect 386842 186496 390172 186552
rect 386781 186494 390172 186496
rect 386781 186491 386847 186494
rect 323669 185058 323735 185061
rect 328494 185058 328500 185060
rect 323669 185056 328500 185058
rect 323669 185000 323674 185056
rect 323730 185000 328500 185056
rect 323669 184998 328500 185000
rect 323669 184995 323735 184998
rect 328494 184996 328500 184998
rect 328564 184996 328570 185060
rect 167729 184378 167795 184381
rect 354765 184378 354831 184381
rect 167729 184376 354831 184378
rect 167729 184320 167734 184376
rect 167790 184320 354770 184376
rect 354826 184320 354831 184376
rect 167729 184318 354831 184320
rect 167729 184315 167795 184318
rect 354765 184315 354831 184318
rect 127617 184242 127683 184245
rect 331806 184242 331812 184244
rect 127617 184240 331812 184242
rect 127617 184184 127622 184240
rect 127678 184184 331812 184240
rect 127617 184182 331812 184184
rect 127617 184179 127683 184182
rect 331806 184180 331812 184182
rect 331876 184180 331882 184244
rect 571425 183834 571491 183837
rect 569940 183832 571491 183834
rect 569940 183776 571430 183832
rect 571486 183776 571491 183832
rect 569940 183774 571491 183776
rect 571425 183771 571491 183774
rect 41321 183018 41387 183021
rect 171174 183018 171180 183020
rect 41321 183016 171180 183018
rect 41321 182960 41326 183016
rect 41382 182960 171180 183016
rect 41321 182958 171180 182960
rect 41321 182955 41387 182958
rect 171174 182956 171180 182958
rect 171244 182956 171250 183020
rect 229737 183018 229803 183021
rect 261150 183018 261156 183020
rect 229737 183016 261156 183018
rect 229737 182960 229742 183016
rect 229798 182960 261156 183016
rect 229737 182958 261156 182960
rect 229737 182955 229803 182958
rect 261150 182956 261156 182958
rect 261220 182956 261226 183020
rect 386413 183018 386479 183021
rect 386413 183016 390172 183018
rect 386413 182960 386418 183016
rect 386474 182960 390172 183016
rect 386413 182958 390172 182960
rect 386413 182955 386479 182958
rect 123477 182882 123543 182885
rect 327574 182882 327580 182884
rect 123477 182880 327580 182882
rect 123477 182824 123482 182880
rect 123538 182824 327580 182880
rect 123477 182822 327580 182824
rect 123477 182819 123543 182822
rect 327574 182820 327580 182822
rect 327644 182820 327650 182884
rect 125041 181658 125107 181661
rect 167494 181658 167500 181660
rect 125041 181656 167500 181658
rect 125041 181600 125046 181656
rect 125102 181600 167500 181656
rect 125041 181598 167500 181600
rect 125041 181595 125107 181598
rect 167494 181596 167500 181598
rect 167564 181596 167570 181660
rect 238017 181658 238083 181661
rect 260782 181658 260788 181660
rect 238017 181656 260788 181658
rect 238017 181600 238022 181656
rect 238078 181600 260788 181656
rect 238017 181598 260788 181600
rect 238017 181595 238083 181598
rect 260782 181596 260788 181598
rect 260852 181596 260858 181660
rect 64781 181522 64847 181525
rect 251214 181522 251220 181524
rect 64781 181520 251220 181522
rect 64781 181464 64786 181520
rect 64842 181464 251220 181520
rect 64781 181462 251220 181464
rect 64781 181459 64847 181462
rect 251214 181460 251220 181462
rect 251284 181460 251290 181524
rect 74533 181386 74599 181389
rect 262254 181386 262260 181388
rect 74533 181384 262260 181386
rect 74533 181328 74538 181384
rect 74594 181328 262260 181384
rect 74533 181326 262260 181328
rect 74533 181323 74599 181326
rect 262254 181324 262260 181326
rect 262324 181324 262330 181388
rect 570137 180298 570203 180301
rect 569940 180296 570203 180298
rect 569940 180240 570142 180296
rect 570198 180240 570203 180296
rect 569940 180238 570203 180240
rect 570137 180235 570203 180238
rect 164141 180026 164207 180029
rect 211797 180026 211863 180029
rect 164141 180024 211863 180026
rect 164141 179968 164146 180024
rect 164202 179968 211802 180024
rect 211858 179968 211863 180024
rect 164141 179966 211863 179968
rect 164141 179963 164207 179966
rect 211797 179963 211863 179966
rect 310421 180026 310487 180029
rect 332542 180026 332548 180028
rect 310421 180024 332548 180026
rect 310421 179968 310426 180024
rect 310482 179968 332548 180024
rect 310421 179966 332548 179968
rect 310421 179963 310487 179966
rect 332542 179964 332548 179966
rect 332612 179964 332618 180028
rect 386873 179618 386939 179621
rect 386873 179616 390172 179618
rect 386873 179560 386878 179616
rect 386934 179560 390172 179616
rect 386873 179558 390172 179560
rect 386873 179555 386939 179558
rect 110413 179482 110479 179485
rect 383009 179482 383075 179485
rect 110413 179480 383075 179482
rect 110413 179424 110418 179480
rect 110474 179424 383014 179480
rect 383070 179424 383075 179480
rect 110413 179422 383075 179424
rect 110413 179419 110479 179422
rect 383009 179419 383075 179422
rect 246389 179210 246455 179213
rect 249006 179210 249012 179212
rect 246389 179208 249012 179210
rect 246389 179152 246394 179208
rect 246450 179152 249012 179208
rect 246389 179150 249012 179152
rect 246389 179147 246455 179150
rect 249006 179148 249012 179150
rect 249076 179148 249082 179212
rect 580441 179210 580507 179213
rect 583520 179210 584960 179300
rect 580441 179208 584960 179210
rect 580441 179152 580446 179208
rect 580502 179152 584960 179208
rect 580441 179150 584960 179152
rect 580441 179147 580507 179150
rect 583520 179060 584960 179150
rect 166257 178802 166323 178805
rect 359549 178802 359615 178805
rect 166257 178800 359615 178802
rect 166257 178744 166262 178800
rect 166318 178744 359554 178800
rect 359610 178744 359615 178800
rect 166257 178742 359615 178744
rect 166257 178739 166323 178742
rect 359549 178739 359615 178742
rect 98637 178666 98703 178669
rect 326429 178666 326495 178669
rect 98637 178664 326495 178666
rect 98637 178608 98642 178664
rect 98698 178608 326434 178664
rect 326490 178608 326495 178664
rect 98637 178606 326495 178608
rect 98637 178603 98703 178606
rect 326429 178603 326495 178606
rect 166390 178122 166396 178124
rect 97030 178062 166396 178122
rect 97030 177988 97090 178062
rect 166390 178060 166396 178062
rect 166460 178060 166466 178124
rect 273846 178060 273852 178124
rect 273916 178122 273922 178124
rect 316033 178122 316099 178125
rect 317321 178122 317387 178125
rect 273916 178120 317387 178122
rect 273916 178064 316038 178120
rect 316094 178064 317326 178120
rect 317382 178064 317387 178120
rect 273916 178062 317387 178064
rect 273916 178060 273922 178062
rect 316033 178059 316099 178062
rect 317321 178059 317387 178062
rect 97022 177924 97028 177988
rect 97092 177924 97098 177988
rect 100702 177652 100708 177716
rect 100772 177714 100778 177716
rect 102041 177714 102107 177717
rect 100772 177712 102107 177714
rect 100772 177656 102046 177712
rect 102102 177656 102107 177712
rect 100772 177654 102107 177656
rect 100772 177652 100778 177654
rect 102041 177651 102107 177654
rect 99414 177516 99420 177580
rect 99484 177578 99490 177580
rect 100661 177578 100727 177581
rect 99484 177576 100727 177578
rect 99484 177520 100666 177576
rect 100722 177520 100727 177576
rect 99484 177518 100727 177520
rect 99484 177516 99490 177518
rect 100661 177515 100727 177518
rect 103278 177516 103284 177580
rect 103348 177578 103354 177580
rect 103421 177578 103487 177581
rect 110689 177580 110755 177581
rect 110638 177578 110644 177580
rect 103348 177576 103487 177578
rect 103348 177520 103426 177576
rect 103482 177520 103487 177576
rect 103348 177518 103487 177520
rect 110598 177518 110644 177578
rect 110708 177576 110755 177580
rect 110750 177520 110755 177576
rect 103348 177516 103354 177518
rect 103421 177515 103487 177518
rect 110638 177516 110644 177518
rect 110708 177516 110755 177520
rect 112110 177516 112116 177580
rect 112180 177578 112186 177580
rect 112989 177578 113055 177581
rect 115841 177580 115907 177581
rect 115790 177578 115796 177580
rect 112180 177576 113055 177578
rect 112180 177520 112994 177576
rect 113050 177520 113055 177576
rect 112180 177518 113055 177520
rect 115750 177518 115796 177578
rect 115860 177576 115907 177580
rect 115902 177520 115907 177576
rect 112180 177516 112186 177518
rect 110689 177515 110755 177516
rect 112989 177515 113055 177518
rect 115790 177516 115796 177518
rect 115860 177516 115907 177520
rect 119654 177516 119660 177580
rect 119724 177578 119730 177580
rect 119981 177578 120047 177581
rect 119724 177576 120047 177578
rect 119724 177520 119986 177576
rect 120042 177520 120047 177576
rect 119724 177518 120047 177520
rect 119724 177516 119730 177518
rect 115841 177515 115907 177516
rect 119981 177515 120047 177518
rect 120758 177516 120764 177580
rect 120828 177578 120834 177580
rect 121085 177578 121151 177581
rect 120828 177576 121151 177578
rect 120828 177520 121090 177576
rect 121146 177520 121151 177576
rect 120828 177518 121151 177520
rect 120828 177516 120834 177518
rect 121085 177515 121151 177518
rect 125726 177516 125732 177580
rect 125796 177578 125802 177580
rect 126881 177578 126947 177581
rect 125796 177576 126947 177578
rect 125796 177520 126886 177576
rect 126942 177520 126947 177576
rect 125796 177518 126947 177520
rect 125796 177516 125802 177518
rect 126881 177515 126947 177518
rect 127014 177516 127020 177580
rect 127084 177578 127090 177580
rect 128077 177578 128143 177581
rect 130745 177580 130811 177581
rect 130694 177578 130700 177580
rect 127084 177576 128143 177578
rect 127084 177520 128082 177576
rect 128138 177520 128143 177576
rect 127084 177518 128143 177520
rect 130654 177518 130700 177578
rect 130764 177576 130811 177580
rect 130806 177520 130811 177576
rect 127084 177516 127090 177518
rect 128077 177515 128143 177518
rect 130694 177516 130700 177518
rect 130764 177516 130811 177520
rect 130745 177515 130811 177516
rect 233877 177578 233943 177581
rect 249190 177578 249196 177580
rect 233877 177576 249196 177578
rect 233877 177520 233882 177576
rect 233938 177520 249196 177576
rect 233877 177518 249196 177520
rect 233877 177515 233943 177518
rect 249190 177516 249196 177518
rect 249260 177516 249266 177580
rect 244273 177442 244339 177445
rect 259678 177442 259684 177444
rect 244273 177440 259684 177442
rect 244273 177384 244278 177440
rect 244334 177384 259684 177440
rect 244273 177382 259684 177384
rect 244273 177379 244339 177382
rect 259678 177380 259684 177382
rect 259748 177380 259754 177444
rect 157977 177306 158043 177309
rect 254209 177306 254275 177309
rect 157977 177304 254275 177306
rect 157977 177248 157982 177304
rect 158038 177248 254214 177304
rect 254270 177248 254275 177304
rect 157977 177246 254275 177248
rect 157977 177243 158043 177246
rect 254209 177243 254275 177246
rect 313917 177306 313983 177309
rect 327022 177306 327028 177308
rect 313917 177304 327028 177306
rect 313917 177248 313922 177304
rect 313978 177248 327028 177304
rect 313917 177246 327028 177248
rect 313917 177243 313983 177246
rect 327022 177244 327028 177246
rect 327092 177244 327098 177308
rect 109534 176972 109540 177036
rect 109604 177034 109610 177036
rect 110229 177034 110295 177037
rect 109604 177032 110295 177034
rect 109604 176976 110234 177032
rect 110290 176976 110295 177032
rect 109604 176974 110295 176976
rect 109604 176972 109610 176974
rect 110229 176971 110295 176974
rect 113214 176972 113220 177036
rect 113284 177034 113290 177036
rect 114369 177034 114435 177037
rect 132033 177036 132099 177037
rect 131982 177034 131988 177036
rect 113284 177032 114435 177034
rect 113284 176976 114374 177032
rect 114430 176976 114435 177032
rect 113284 176974 114435 176976
rect 131942 176974 131988 177034
rect 132052 177032 132099 177036
rect 572069 177034 572135 177037
rect 132094 176976 132099 177032
rect 113284 176972 113290 176974
rect 114369 176971 114435 176974
rect 131982 176972 131988 176974
rect 132052 176972 132099 176976
rect 569940 177032 572135 177034
rect 569940 176976 572074 177032
rect 572130 176976 572135 177032
rect 569940 176974 572135 176976
rect 132033 176971 132099 176972
rect 572069 176971 572135 176974
rect 101990 176836 101996 176900
rect 102060 176898 102066 176900
rect 166993 176898 167059 176901
rect 102060 176896 167059 176898
rect 102060 176840 166998 176896
rect 167054 176840 167059 176896
rect 102060 176838 167059 176840
rect 102060 176836 102066 176838
rect 166993 176835 167059 176838
rect 104617 176764 104683 176765
rect 107009 176764 107075 176765
rect 108113 176764 108179 176765
rect 118417 176764 118483 176765
rect 104566 176762 104572 176764
rect 104526 176702 104572 176762
rect 104636 176760 104683 176764
rect 106958 176762 106964 176764
rect 104678 176704 104683 176760
rect 104566 176700 104572 176702
rect 104636 176700 104683 176704
rect 106918 176702 106964 176762
rect 107028 176760 107075 176764
rect 108062 176762 108068 176764
rect 107070 176704 107075 176760
rect 106958 176700 106964 176702
rect 107028 176700 107075 176704
rect 108022 176702 108068 176762
rect 108132 176760 108179 176764
rect 118366 176762 118372 176764
rect 108174 176704 108179 176760
rect 108062 176700 108068 176702
rect 108132 176700 108179 176704
rect 118326 176702 118372 176762
rect 118436 176760 118483 176764
rect 118478 176704 118483 176760
rect 118366 176700 118372 176702
rect 118436 176700 118483 176704
rect 121862 176700 121868 176764
rect 121932 176762 121938 176764
rect 122741 176762 122807 176765
rect 123017 176764 123083 176765
rect 121932 176760 122807 176762
rect 121932 176704 122746 176760
rect 122802 176704 122807 176760
rect 121932 176702 122807 176704
rect 121932 176700 121938 176702
rect 104617 176699 104683 176700
rect 107009 176699 107075 176700
rect 108113 176699 108179 176700
rect 118417 176699 118483 176700
rect 122741 176699 122807 176702
rect 122966 176700 122972 176764
rect 123036 176762 123083 176764
rect 128169 176762 128235 176765
rect 129457 176764 129523 176765
rect 133137 176764 133203 176765
rect 135713 176764 135779 176765
rect 148225 176764 148291 176765
rect 129406 176762 129412 176764
rect 123036 176760 123128 176762
rect 123078 176704 123128 176760
rect 123036 176702 123128 176704
rect 128126 176760 128235 176762
rect 128126 176704 128174 176760
rect 128230 176704 128235 176760
rect 123036 176700 123083 176702
rect 123017 176699 123083 176700
rect 128126 176699 128235 176704
rect 129366 176702 129412 176762
rect 129476 176760 129523 176764
rect 133086 176762 133092 176764
rect 129518 176704 129523 176760
rect 129406 176700 129412 176702
rect 129476 176700 129523 176704
rect 133046 176702 133092 176762
rect 133156 176760 133203 176764
rect 135662 176762 135668 176764
rect 133198 176704 133203 176760
rect 133086 176700 133092 176702
rect 133156 176700 133203 176704
rect 135622 176702 135668 176762
rect 135732 176760 135779 176764
rect 148174 176762 148180 176764
rect 135774 176704 135779 176760
rect 135662 176700 135668 176702
rect 135732 176700 135779 176704
rect 148134 176702 148180 176762
rect 148244 176760 148291 176764
rect 148286 176704 148291 176760
rect 148174 176700 148180 176702
rect 148244 176700 148291 176704
rect 158846 176700 158852 176764
rect 158916 176762 158922 176764
rect 158989 176762 159055 176765
rect 158916 176760 159055 176762
rect 158916 176704 158994 176760
rect 159050 176704 159055 176760
rect 158916 176702 159055 176704
rect 158916 176700 158922 176702
rect 129457 176699 129523 176700
rect 133137 176699 133203 176700
rect 135713 176699 135779 176700
rect 148225 176699 148291 176700
rect 158989 176699 159055 176702
rect 320173 176762 320239 176765
rect 321318 176762 321324 176764
rect 320173 176760 321324 176762
rect 320173 176704 320178 176760
rect 320234 176704 321324 176760
rect 320173 176702 321324 176704
rect 320173 176699 320239 176702
rect 321318 176700 321324 176702
rect 321388 176700 321394 176764
rect 128126 176492 128186 176699
rect 128118 176428 128124 176492
rect 128188 176428 128194 176492
rect 255313 176490 255379 176493
rect 255446 176490 255452 176492
rect 255313 176488 255452 176490
rect 255313 176432 255318 176488
rect 255374 176432 255452 176488
rect 255313 176430 255452 176432
rect 255313 176427 255379 176430
rect 255446 176428 255452 176430
rect 255516 176428 255522 176492
rect 387006 176292 387012 176356
rect 387076 176354 387082 176356
rect 387076 176294 390172 176354
rect 387076 176292 387082 176294
rect 247677 176082 247743 176085
rect 252686 176082 252692 176084
rect 247677 176080 252692 176082
rect -960 175796 480 176036
rect 247677 176024 247682 176080
rect 247738 176024 252692 176080
rect 247677 176022 252692 176024
rect 247677 176019 247743 176022
rect 252686 176020 252692 176022
rect 252756 176020 252762 176084
rect 318149 176082 318215 176085
rect 328678 176082 328684 176084
rect 318149 176080 328684 176082
rect 318149 176024 318154 176080
rect 318210 176024 328684 176080
rect 318149 176022 328684 176024
rect 318149 176019 318215 176022
rect 328678 176020 328684 176022
rect 328748 176020 328754 176084
rect 232497 175946 232563 175949
rect 257838 175946 257844 175948
rect 232497 175944 257844 175946
rect 232497 175888 232502 175944
rect 232558 175888 257844 175944
rect 232497 175886 257844 175888
rect 232497 175883 232563 175886
rect 257838 175884 257844 175886
rect 257908 175884 257914 175948
rect 271086 175884 271092 175948
rect 271156 175946 271162 175948
rect 306373 175946 306439 175949
rect 315481 175946 315547 175949
rect 342294 175946 342300 175948
rect 271156 175944 310162 175946
rect 271156 175888 306378 175944
rect 306434 175888 310162 175944
rect 271156 175886 310162 175888
rect 271156 175884 271162 175886
rect 306373 175883 306439 175886
rect 248045 175810 248111 175813
rect 248045 175808 248338 175810
rect 248045 175752 248050 175808
rect 248106 175752 248338 175808
rect 248045 175750 248338 175752
rect 248045 175747 248111 175750
rect 116945 175676 117011 175677
rect 124489 175676 124555 175677
rect 134425 175676 134491 175677
rect 116894 175674 116900 175676
rect 116854 175614 116900 175674
rect 116964 175672 117011 175676
rect 124438 175674 124444 175676
rect 117006 175616 117011 175672
rect 116894 175612 116900 175614
rect 116964 175612 117011 175616
rect 124398 175614 124444 175674
rect 124508 175672 124555 175676
rect 134374 175674 134380 175676
rect 124550 175616 124555 175672
rect 124438 175612 124444 175614
rect 124508 175612 124555 175616
rect 134334 175614 134380 175674
rect 134444 175672 134491 175676
rect 134486 175616 134491 175672
rect 134374 175612 134380 175614
rect 134444 175612 134491 175616
rect 116945 175611 117011 175612
rect 124489 175611 124555 175612
rect 134425 175611 134491 175612
rect 213913 175674 213979 175677
rect 213913 175672 217212 175674
rect 213913 175616 213918 175672
rect 213974 175616 217212 175672
rect 248278 175644 248338 175750
rect 310102 175644 310162 175886
rect 315481 175944 342300 175946
rect 315481 175888 315486 175944
rect 315542 175888 342300 175944
rect 315481 175886 342300 175888
rect 315481 175883 315547 175886
rect 342294 175884 342300 175886
rect 342364 175884 342370 175948
rect 387558 175884 387564 175948
rect 387628 175946 387634 175948
rect 387793 175946 387859 175949
rect 387628 175944 387859 175946
rect 387628 175888 387798 175944
rect 387854 175888 387859 175944
rect 387628 175886 387859 175888
rect 387628 175884 387634 175886
rect 387793 175883 387859 175886
rect 213913 175614 217212 175616
rect 213913 175611 213979 175614
rect 114318 175476 114324 175540
rect 114388 175538 114394 175540
rect 166206 175538 166212 175540
rect 114388 175478 166212 175538
rect 114388 175476 114394 175478
rect 166206 175476 166212 175478
rect 166276 175476 166282 175540
rect 324313 175538 324379 175541
rect 321908 175536 324379 175538
rect 321908 175480 324318 175536
rect 324374 175480 324379 175536
rect 321908 175478 324379 175480
rect 324313 175475 324379 175478
rect 98361 175404 98427 175405
rect 98310 175402 98316 175404
rect 98270 175342 98316 175402
rect 98380 175400 98427 175404
rect 98422 175344 98427 175400
rect 98310 175340 98316 175342
rect 98380 175340 98427 175344
rect 105670 175340 105676 175404
rect 105740 175402 105746 175404
rect 167678 175402 167684 175404
rect 105740 175342 167684 175402
rect 105740 175340 105746 175342
rect 167678 175340 167684 175342
rect 167748 175340 167754 175404
rect 98361 175339 98427 175340
rect 249149 175266 249215 175269
rect 248860 175264 249215 175266
rect 248860 175208 249154 175264
rect 249210 175208 249215 175264
rect 248860 175206 249215 175208
rect 249149 175203 249215 175206
rect 306966 175204 306972 175268
rect 307036 175266 307042 175268
rect 307036 175206 310132 175266
rect 307036 175204 307042 175206
rect 213913 174994 213979 174997
rect 213913 174992 217212 174994
rect 213913 174936 213918 174992
rect 213974 174936 217212 174992
rect 213913 174934 217212 174936
rect 213913 174931 213979 174934
rect 306741 174858 306807 174861
rect 306741 174856 310132 174858
rect 306741 174800 306746 174856
rect 306802 174800 310132 174856
rect 306741 174798 310132 174800
rect 306741 174795 306807 174798
rect 249374 174722 249380 174724
rect 248860 174662 249380 174722
rect 249374 174660 249380 174662
rect 249444 174660 249450 174724
rect 325049 174722 325115 174725
rect 321908 174720 325115 174722
rect 321908 174664 325054 174720
rect 325110 174664 325115 174720
rect 321908 174662 325115 174664
rect 325049 174659 325115 174662
rect 307661 174450 307727 174453
rect 307661 174448 310132 174450
rect 307661 174392 307666 174448
rect 307722 174392 310132 174448
rect 307661 174390 310132 174392
rect 307661 174387 307727 174390
rect 214005 174314 214071 174317
rect 254526 174314 254532 174316
rect 214005 174312 217212 174314
rect 214005 174256 214010 174312
rect 214066 174256 217212 174312
rect 214005 174254 217212 174256
rect 248860 174254 254532 174314
rect 214005 174251 214071 174254
rect 254526 174252 254532 174254
rect 254596 174252 254602 174316
rect 307293 174042 307359 174045
rect 324313 174042 324379 174045
rect 307293 174040 310132 174042
rect 307293 173984 307298 174040
rect 307354 173984 310132 174040
rect 307293 173982 310132 173984
rect 321908 174040 324379 174042
rect 321908 173984 324318 174040
rect 324374 173984 324379 174040
rect 321908 173982 324379 173984
rect 307293 173979 307359 173982
rect 324313 173979 324379 173982
rect 326654 173906 326660 173908
rect 325650 173846 326660 173906
rect 249190 173770 249196 173772
rect 248860 173710 249196 173770
rect 249190 173708 249196 173710
rect 249260 173708 249266 173772
rect 325650 173770 325710 173846
rect 326654 173844 326660 173846
rect 326724 173906 326730 173908
rect 382917 173906 382983 173909
rect 326724 173904 382983 173906
rect 326724 173848 382922 173904
rect 382978 173848 382983 173904
rect 326724 173846 382983 173848
rect 326724 173844 326730 173846
rect 382917 173843 382983 173846
rect 569534 173844 569540 173908
rect 569604 173844 569610 173908
rect 321878 173710 325710 173770
rect 213913 173634 213979 173637
rect 307569 173634 307635 173637
rect 213913 173632 217212 173634
rect 213913 173576 213918 173632
rect 213974 173576 217212 173632
rect 213913 173574 217212 173576
rect 307569 173632 310132 173634
rect 307569 173576 307574 173632
rect 307630 173576 310132 173632
rect 307569 173574 310132 173576
rect 213913 173571 213979 173574
rect 307569 173571 307635 173574
rect 249333 173362 249399 173365
rect 248860 173360 249399 173362
rect 248860 173304 249338 173360
rect 249394 173304 249399 173360
rect 248860 173302 249399 173304
rect 249333 173299 249399 173302
rect 307293 173226 307359 173229
rect 307293 173224 310132 173226
rect 307293 173168 307298 173224
rect 307354 173168 310132 173224
rect 321878 173196 321938 173710
rect 569542 173604 569602 173844
rect 307293 173166 310132 173168
rect 307293 173163 307359 173166
rect 214005 172954 214071 172957
rect 387149 172954 387215 172957
rect 214005 172952 217212 172954
rect 214005 172896 214010 172952
rect 214066 172896 217212 172952
rect 214005 172894 217212 172896
rect 387149 172952 390172 172954
rect 387149 172896 387154 172952
rect 387210 172896 390172 172952
rect 387149 172894 390172 172896
rect 214005 172891 214071 172894
rect 387149 172891 387215 172894
rect 249425 172818 249491 172821
rect 248860 172816 249491 172818
rect 248860 172760 249430 172816
rect 249486 172760 249491 172816
rect 248860 172758 249491 172760
rect 249425 172755 249491 172758
rect 307661 172682 307727 172685
rect 307661 172680 310132 172682
rect 307661 172624 307666 172680
rect 307722 172624 310132 172680
rect 307661 172622 310132 172624
rect 307661 172619 307727 172622
rect 251817 172410 251883 172413
rect 248860 172408 251883 172410
rect 248860 172352 251822 172408
rect 251878 172352 251883 172408
rect 248860 172350 251883 172352
rect 251817 172347 251883 172350
rect 214189 172274 214255 172277
rect 306925 172274 306991 172277
rect 214189 172272 217212 172274
rect 214189 172216 214194 172272
rect 214250 172216 217212 172272
rect 214189 172214 217212 172216
rect 306925 172272 310132 172274
rect 306925 172216 306930 172272
rect 306986 172216 310132 172272
rect 306925 172214 310132 172216
rect 214189 172211 214255 172214
rect 306925 172211 306991 172214
rect 321326 172140 321386 172380
rect 321318 172076 321324 172140
rect 321388 172138 321394 172140
rect 324865 172138 324931 172141
rect 321388 172136 324931 172138
rect 321388 172080 324870 172136
rect 324926 172080 324931 172136
rect 321388 172078 324931 172080
rect 321388 172076 321394 172078
rect 324865 172075 324931 172078
rect 249241 171866 249307 171869
rect 248860 171864 249307 171866
rect 248860 171808 249246 171864
rect 249302 171808 249307 171864
rect 248860 171806 249307 171808
rect 249241 171803 249307 171806
rect 306557 171866 306623 171869
rect 306557 171864 310132 171866
rect 306557 171808 306562 171864
rect 306618 171808 310132 171864
rect 306557 171806 310132 171808
rect 306557 171803 306623 171806
rect 170254 171668 170260 171732
rect 170324 171730 170330 171732
rect 206369 171730 206435 171733
rect 324313 171730 324379 171733
rect 170324 171728 206435 171730
rect 170324 171672 206374 171728
rect 206430 171672 206435 171728
rect 170324 171670 206435 171672
rect 321908 171728 324379 171730
rect 321908 171672 324318 171728
rect 324374 171672 324379 171728
rect 321908 171670 324379 171672
rect 170324 171668 170330 171670
rect 206369 171667 206435 171670
rect 324313 171667 324379 171670
rect 167637 171594 167703 171597
rect 164694 171592 167703 171594
rect 164694 171536 167642 171592
rect 167698 171536 167703 171592
rect 164694 171534 167703 171536
rect -960 162890 480 162980
rect 3693 162890 3759 162893
rect -960 162888 3759 162890
rect -960 162832 3698 162888
rect 3754 162832 3759 162888
rect -960 162830 3759 162832
rect -960 162740 480 162830
rect 3693 162827 3759 162830
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect -960 136778 480 136868
rect 3233 136778 3299 136781
rect -960 136776 3299 136778
rect -960 136720 3238 136776
rect 3294 136720 3299 136776
rect -960 136718 3299 136720
rect -960 136628 480 136718
rect 3233 136715 3299 136718
rect 167637 171531 167703 171534
rect 214097 171594 214163 171597
rect 214097 171592 217212 171594
rect 214097 171536 214102 171592
rect 214158 171536 217212 171592
rect 214097 171534 217212 171536
rect 214097 171531 214163 171534
rect 252553 171458 252619 171461
rect 248860 171456 252619 171458
rect 248860 171400 252558 171456
rect 252614 171400 252619 171456
rect 248860 171398 252619 171400
rect 252553 171395 252619 171398
rect 307661 171458 307727 171461
rect 307661 171456 310132 171458
rect 307661 171400 307666 171456
rect 307722 171400 310132 171456
rect 307661 171398 310132 171400
rect 307661 171395 307727 171398
rect 214741 171050 214807 171053
rect 307385 171050 307451 171053
rect 214741 171048 217212 171050
rect 214741 170992 214746 171048
rect 214802 170992 217212 171048
rect 214741 170990 217212 170992
rect 307385 171048 310132 171050
rect 307385 170992 307390 171048
rect 307446 170992 310132 171048
rect 307385 170990 310132 170992
rect 214741 170987 214807 170990
rect 307385 170987 307451 170990
rect 251725 170914 251791 170917
rect 324313 170914 324379 170917
rect 248860 170912 251791 170914
rect 248860 170856 251730 170912
rect 251786 170856 251791 170912
rect 248860 170854 251791 170856
rect 321908 170912 324379 170914
rect 321908 170856 324318 170912
rect 324374 170856 324379 170912
rect 321908 170854 324379 170856
rect 251725 170851 251791 170854
rect 324313 170851 324379 170854
rect 306741 170642 306807 170645
rect 306741 170640 310132 170642
rect 306741 170584 306746 170640
rect 306802 170584 310132 170640
rect 306741 170582 310132 170584
rect 306741 170579 306807 170582
rect 251817 170506 251883 170509
rect 248860 170504 251883 170506
rect 248860 170448 251822 170504
rect 251878 170448 251883 170504
rect 248860 170446 251883 170448
rect 251817 170443 251883 170446
rect 213913 170370 213979 170373
rect 213913 170368 217212 170370
rect 213913 170312 213918 170368
rect 213974 170312 217212 170368
rect 213913 170310 217212 170312
rect 213913 170307 213979 170310
rect 321318 170308 321324 170372
rect 321388 170370 321394 170372
rect 321388 170310 321938 170370
rect 321388 170308 321394 170310
rect 307661 170234 307727 170237
rect 307661 170232 310132 170234
rect 307661 170176 307666 170232
rect 307722 170176 310132 170232
rect 307661 170174 310132 170176
rect 307661 170171 307727 170174
rect 252502 170098 252508 170100
rect 248860 170038 252508 170098
rect 252502 170036 252508 170038
rect 252572 170036 252578 170100
rect 321878 170098 321938 170310
rect 324313 170098 324379 170101
rect 572621 170098 572687 170101
rect 321878 170096 324379 170098
rect 321878 170068 324318 170096
rect 321908 170040 324318 170068
rect 324374 170040 324379 170096
rect 321908 170038 324379 170040
rect 569940 170096 572687 170098
rect 569940 170040 572626 170096
rect 572682 170040 572687 170096
rect 569940 170038 572687 170040
rect 324313 170035 324379 170038
rect 572621 170035 572687 170038
rect 307293 169826 307359 169829
rect 307293 169824 310132 169826
rect 307293 169768 307298 169824
rect 307354 169768 310132 169824
rect 307293 169766 310132 169768
rect 307293 169763 307359 169766
rect 213913 169690 213979 169693
rect 213913 169688 217212 169690
rect 213913 169632 213918 169688
rect 213974 169632 217212 169688
rect 213913 169630 217212 169632
rect 213913 169627 213979 169630
rect 252737 169554 252803 169557
rect 248860 169552 252803 169554
rect 248860 169496 252742 169552
rect 252798 169496 252803 169552
rect 248860 169494 252803 169496
rect 252737 169491 252803 169494
rect 386873 169554 386939 169557
rect 386873 169552 390172 169554
rect 386873 169496 386878 169552
rect 386934 169496 390172 169552
rect 386873 169494 390172 169496
rect 386873 169491 386939 169494
rect 324313 169418 324379 169421
rect 321908 169416 324379 169418
rect 321908 169360 324318 169416
rect 324374 169360 324379 169416
rect 321908 169358 324379 169360
rect 324313 169355 324379 169358
rect 306741 169282 306807 169285
rect 306741 169280 310132 169282
rect 306741 169224 306746 169280
rect 306802 169224 310132 169280
rect 306741 169222 310132 169224
rect 306741 169219 306807 169222
rect 252461 169146 252527 169149
rect 248860 169144 252527 169146
rect 248860 169088 252466 169144
rect 252522 169088 252527 169144
rect 248860 169086 252527 169088
rect 252461 169083 252527 169086
rect 214005 169010 214071 169013
rect 214005 169008 217212 169010
rect 214005 168952 214010 169008
rect 214066 168952 217212 169008
rect 214005 168950 217212 168952
rect 214005 168947 214071 168950
rect 307569 168874 307635 168877
rect 307569 168872 310132 168874
rect 307569 168816 307574 168872
rect 307630 168816 310132 168872
rect 307569 168814 310132 168816
rect 307569 168811 307635 168814
rect 257838 168602 257844 168604
rect 248860 168542 257844 168602
rect 257838 168540 257844 168542
rect 257908 168540 257914 168604
rect 324497 168602 324563 168605
rect 321908 168600 324563 168602
rect 321908 168544 324502 168600
rect 324558 168544 324563 168600
rect 321908 168542 324563 168544
rect 324497 168539 324563 168542
rect 307293 168466 307359 168469
rect 307293 168464 310132 168466
rect 307293 168408 307298 168464
rect 307354 168408 310132 168464
rect 307293 168406 310132 168408
rect 307293 168403 307359 168406
rect 214005 168330 214071 168333
rect 214005 168328 217212 168330
rect 214005 168272 214010 168328
rect 214066 168272 217212 168328
rect 214005 168270 217212 168272
rect 214005 168267 214071 168270
rect 252461 168194 252527 168197
rect 248860 168192 252527 168194
rect 248860 168136 252466 168192
rect 252522 168136 252527 168192
rect 248860 168134 252527 168136
rect 252461 168131 252527 168134
rect 307293 168058 307359 168061
rect 307293 168056 310132 168058
rect 307293 168000 307298 168056
rect 307354 168000 310132 168056
rect 307293 167998 310132 168000
rect 307293 167995 307359 167998
rect 324405 167786 324471 167789
rect 321908 167784 324471 167786
rect 321908 167728 324410 167784
rect 324466 167728 324471 167784
rect 321908 167726 324471 167728
rect 324405 167723 324471 167726
rect 213913 167650 213979 167653
rect 252461 167650 252527 167653
rect 213913 167648 217212 167650
rect 213913 167592 213918 167648
rect 213974 167592 217212 167648
rect 213913 167590 217212 167592
rect 248860 167648 252527 167650
rect 248860 167592 252466 167648
rect 252522 167592 252527 167648
rect 248860 167590 252527 167592
rect 213913 167587 213979 167590
rect 252461 167587 252527 167590
rect 307661 167650 307727 167653
rect 307661 167648 310132 167650
rect 307661 167592 307666 167648
rect 307722 167592 310132 167648
rect 307661 167590 310132 167592
rect 307661 167587 307727 167590
rect 252369 167242 252435 167245
rect 248860 167240 252435 167242
rect 248860 167184 252374 167240
rect 252430 167184 252435 167240
rect 248860 167182 252435 167184
rect 252369 167179 252435 167182
rect 307477 167242 307543 167245
rect 307477 167240 310132 167242
rect 307477 167184 307482 167240
rect 307538 167184 310132 167240
rect 307477 167182 310132 167184
rect 307477 167179 307543 167182
rect 324313 167106 324379 167109
rect 321908 167104 324379 167106
rect 321908 167048 324318 167104
rect 324374 167048 324379 167104
rect 321908 167046 324379 167048
rect 324313 167043 324379 167046
rect 213913 166970 213979 166973
rect 213913 166968 217212 166970
rect 213913 166912 213918 166968
rect 213974 166912 217212 166968
rect 213913 166910 217212 166912
rect 213913 166907 213979 166910
rect 307661 166834 307727 166837
rect 307661 166832 310132 166834
rect 307661 166776 307666 166832
rect 307722 166776 310132 166832
rect 307661 166774 310132 166776
rect 307661 166771 307727 166774
rect 252369 166698 252435 166701
rect 572345 166698 572411 166701
rect 248860 166696 252435 166698
rect 248860 166640 252374 166696
rect 252430 166640 252435 166696
rect 248860 166638 252435 166640
rect 569940 166696 572411 166698
rect 569940 166640 572350 166696
rect 572406 166640 572411 166696
rect 569940 166638 572411 166640
rect 252369 166635 252435 166638
rect 572345 166635 572411 166638
rect 214097 166426 214163 166429
rect 306557 166426 306623 166429
rect 214097 166424 217212 166426
rect 214097 166368 214102 166424
rect 214158 166368 217212 166424
rect 214097 166366 217212 166368
rect 306557 166424 310132 166426
rect 306557 166368 306562 166424
rect 306618 166368 310132 166424
rect 306557 166366 310132 166368
rect 214097 166363 214163 166366
rect 306557 166363 306623 166366
rect 252461 166290 252527 166293
rect 324313 166290 324379 166293
rect 248860 166288 252527 166290
rect 248860 166232 252466 166288
rect 252522 166232 252527 166288
rect 248860 166230 252527 166232
rect 321908 166288 324379 166290
rect 321908 166232 324318 166288
rect 324374 166232 324379 166288
rect 321908 166230 324379 166232
rect 252461 166227 252527 166230
rect 324313 166227 324379 166230
rect 386873 166154 386939 166157
rect 386873 166152 390172 166154
rect 386873 166096 386878 166152
rect 386934 166096 390172 166152
rect 386873 166094 390172 166096
rect 386873 166091 386939 166094
rect 307477 165882 307543 165885
rect 582649 165882 582715 165885
rect 583520 165882 584960 165972
rect 307477 165880 310132 165882
rect 307477 165824 307482 165880
rect 307538 165824 310132 165880
rect 307477 165822 310132 165824
rect 582649 165880 584960 165882
rect 582649 165824 582654 165880
rect 582710 165824 584960 165880
rect 582649 165822 584960 165824
rect 307477 165819 307543 165822
rect 582649 165819 582715 165822
rect 214005 165746 214071 165749
rect 252277 165746 252343 165749
rect 214005 165744 217212 165746
rect 214005 165688 214010 165744
rect 214066 165688 217212 165744
rect 214005 165686 217212 165688
rect 248860 165744 252343 165746
rect 248860 165688 252282 165744
rect 252338 165688 252343 165744
rect 248860 165686 252343 165688
rect 214005 165683 214071 165686
rect 252277 165683 252343 165686
rect 321277 165746 321343 165749
rect 321277 165744 321570 165746
rect 321277 165688 321282 165744
rect 321338 165688 321570 165744
rect 583520 165732 584960 165822
rect 321277 165686 321570 165688
rect 321277 165683 321343 165686
rect 307569 165474 307635 165477
rect 321510 165474 321570 165686
rect 324313 165474 324379 165477
rect 307569 165472 310132 165474
rect 307569 165416 307574 165472
rect 307630 165416 310132 165472
rect 321510 165472 324379 165474
rect 321510 165444 324318 165472
rect 307569 165414 310132 165416
rect 321540 165416 324318 165444
rect 324374 165416 324379 165472
rect 321540 165414 324379 165416
rect 307569 165411 307635 165414
rect 324313 165411 324379 165414
rect 252461 165338 252527 165341
rect 248860 165336 252527 165338
rect 248860 165280 252466 165336
rect 252522 165280 252527 165336
rect 248860 165278 252527 165280
rect 252461 165275 252527 165278
rect 213913 165066 213979 165069
rect 307109 165066 307175 165069
rect 213913 165064 217212 165066
rect 213913 165008 213918 165064
rect 213974 165008 217212 165064
rect 213913 165006 217212 165008
rect 307109 165064 310132 165066
rect 307109 165008 307114 165064
rect 307170 165008 310132 165064
rect 307109 165006 310132 165008
rect 213913 165003 213979 165006
rect 307109 165003 307175 165006
rect 252461 164794 252527 164797
rect 323117 164794 323183 164797
rect 323393 164794 323459 164797
rect 248860 164792 252527 164794
rect 248860 164736 252466 164792
rect 252522 164736 252527 164792
rect 248860 164734 252527 164736
rect 321908 164792 323459 164794
rect 321908 164736 323122 164792
rect 323178 164736 323398 164792
rect 323454 164736 323459 164792
rect 321908 164734 323459 164736
rect 252461 164731 252527 164734
rect 323117 164731 323183 164734
rect 323393 164731 323459 164734
rect 307661 164658 307727 164661
rect 307661 164656 310132 164658
rect 307661 164600 307666 164656
rect 307722 164600 310132 164656
rect 307661 164598 310132 164600
rect 307661 164595 307727 164598
rect 166206 164324 166212 164388
rect 166276 164386 166282 164388
rect 250161 164386 250227 164389
rect 166276 164326 217212 164386
rect 248860 164384 250227 164386
rect 248860 164328 250166 164384
rect 250222 164328 250227 164384
rect 248860 164326 250227 164328
rect 166276 164324 166282 164326
rect 250161 164323 250227 164326
rect 307293 164250 307359 164253
rect 307293 164248 310132 164250
rect 307293 164192 307298 164248
rect 307354 164192 310132 164248
rect 307293 164190 310132 164192
rect 307293 164187 307359 164190
rect 253197 163978 253263 163981
rect 324313 163978 324379 163981
rect 248860 163976 253263 163978
rect 248860 163920 253202 163976
rect 253258 163920 253263 163976
rect 248860 163918 253263 163920
rect 321908 163976 324379 163978
rect 321908 163920 324318 163976
rect 324374 163920 324379 163976
rect 321908 163918 324379 163920
rect 253197 163915 253263 163918
rect 324313 163915 324379 163918
rect 307477 163842 307543 163845
rect 307477 163840 310132 163842
rect 307477 163784 307482 163840
rect 307538 163784 310132 163840
rect 307477 163782 310132 163784
rect 307477 163779 307543 163782
rect 214005 163706 214071 163709
rect 214005 163704 217212 163706
rect 214005 163648 214010 163704
rect 214066 163648 217212 163704
rect 214005 163646 217212 163648
rect 214005 163643 214071 163646
rect 307661 163434 307727 163437
rect 571333 163434 571399 163437
rect 248860 163374 258090 163434
rect 258030 163162 258090 163374
rect 307661 163432 310132 163434
rect 307661 163376 307666 163432
rect 307722 163376 310132 163432
rect 307661 163374 310132 163376
rect 569940 163432 571399 163434
rect 569940 163376 571338 163432
rect 571394 163376 571399 163432
rect 569940 163374 571399 163376
rect 307661 163371 307727 163374
rect 571333 163371 571399 163374
rect 269062 163162 269068 163164
rect 258030 163102 269068 163162
rect 269062 163100 269068 163102
rect 269132 163100 269138 163164
rect 324405 163162 324471 163165
rect 321908 163160 324471 163162
rect 321908 163104 324410 163160
rect 324466 163104 324471 163160
rect 321908 163102 324471 163104
rect 324405 163099 324471 163102
rect 213913 163026 213979 163029
rect 252185 163026 252251 163029
rect 213913 163024 217212 163026
rect 213913 162968 213918 163024
rect 213974 162968 217212 163024
rect 213913 162966 217212 162968
rect 248860 163024 252251 163026
rect 248860 162968 252190 163024
rect 252246 162968 252251 163024
rect 248860 162966 252251 162968
rect 213913 162963 213979 162966
rect 252185 162963 252251 162966
rect 253197 163026 253263 163029
rect 261150 163026 261156 163028
rect 253197 163024 261156 163026
rect 253197 162968 253202 163024
rect 253258 162968 261156 163024
rect 253197 162966 261156 162968
rect 253197 162963 253263 162966
rect 261150 162964 261156 162966
rect 261220 162964 261226 163028
rect 307201 163026 307267 163029
rect 307201 163024 310132 163026
rect 307201 162968 307206 163024
rect 307262 162968 310132 163024
rect 307201 162966 310132 162968
rect 307201 162963 307267 162966
rect 328678 162754 328684 162756
rect 321878 162694 328684 162754
rect 252093 162482 252159 162485
rect 248860 162480 252159 162482
rect 248860 162424 252098 162480
rect 252154 162424 252159 162480
rect 248860 162422 252159 162424
rect 252093 162419 252159 162422
rect 306741 162482 306807 162485
rect 306741 162480 310132 162482
rect 306741 162424 306746 162480
rect 306802 162424 310132 162480
rect 321878 162452 321938 162694
rect 328678 162692 328684 162694
rect 328748 162754 328754 162756
rect 386873 162754 386939 162757
rect 328748 162694 374010 162754
rect 328748 162692 328754 162694
rect 373950 162482 374010 162694
rect 386873 162752 390172 162754
rect 386873 162696 386878 162752
rect 386934 162696 390172 162752
rect 386873 162694 390172 162696
rect 386873 162691 386939 162694
rect 389817 162482 389883 162485
rect 373950 162480 389883 162482
rect 306741 162422 310132 162424
rect 373950 162424 389822 162480
rect 389878 162424 389883 162480
rect 373950 162422 389883 162424
rect 306741 162419 306807 162422
rect 389817 162419 389883 162422
rect 214557 162346 214623 162349
rect 214557 162344 217212 162346
rect 214557 162288 214562 162344
rect 214618 162288 217212 162344
rect 214557 162286 217212 162288
rect 214557 162283 214623 162286
rect 252461 162074 252527 162077
rect 248860 162072 252527 162074
rect 248860 162016 252466 162072
rect 252522 162016 252527 162072
rect 248860 162014 252527 162016
rect 252461 162011 252527 162014
rect 307661 162074 307727 162077
rect 307661 162072 310132 162074
rect 307661 162016 307666 162072
rect 307722 162016 310132 162072
rect 307661 162014 310132 162016
rect 307661 162011 307727 162014
rect 213913 161802 213979 161805
rect 213913 161800 217212 161802
rect 213913 161744 213918 161800
rect 213974 161744 217212 161800
rect 213913 161742 217212 161744
rect 213913 161739 213979 161742
rect 307477 161666 307543 161669
rect 325877 161666 325943 161669
rect 307477 161664 310132 161666
rect 307477 161608 307482 161664
rect 307538 161608 310132 161664
rect 307477 161606 310132 161608
rect 321908 161664 325943 161666
rect 321908 161608 325882 161664
rect 325938 161608 325943 161664
rect 321908 161606 325943 161608
rect 307477 161603 307543 161606
rect 325877 161603 325943 161606
rect 251541 161530 251607 161533
rect 248860 161528 251607 161530
rect 248860 161472 251546 161528
rect 251602 161472 251607 161528
rect 248860 161470 251607 161472
rect 251541 161467 251607 161470
rect 384481 161394 384547 161397
rect 335310 161392 384547 161394
rect 335310 161336 384486 161392
rect 384542 161336 384547 161392
rect 335310 161334 384547 161336
rect 306741 161258 306807 161261
rect 331489 161258 331555 161261
rect 331806 161258 331812 161260
rect 306741 161256 310132 161258
rect 306741 161200 306746 161256
rect 306802 161200 310132 161256
rect 306741 161198 310132 161200
rect 331489 161256 331812 161258
rect 331489 161200 331494 161256
rect 331550 161200 331812 161256
rect 331489 161198 331812 161200
rect 306741 161195 306807 161198
rect 331489 161195 331555 161198
rect 331806 161196 331812 161198
rect 331876 161258 331882 161260
rect 335310 161258 335370 161334
rect 384481 161331 384547 161334
rect 331876 161198 335370 161258
rect 331876 161196 331882 161198
rect 213913 161122 213979 161125
rect 256918 161122 256924 161124
rect 213913 161120 217212 161122
rect 213913 161064 213918 161120
rect 213974 161064 217212 161120
rect 213913 161062 217212 161064
rect 248860 161062 256924 161122
rect 213913 161059 213979 161062
rect 256918 161060 256924 161062
rect 256988 161060 256994 161124
rect 307569 160850 307635 160853
rect 324313 160850 324379 160853
rect 307569 160848 310132 160850
rect 307569 160792 307574 160848
rect 307630 160792 310132 160848
rect 307569 160790 310132 160792
rect 321908 160848 324379 160850
rect 321908 160792 324318 160848
rect 324374 160792 324379 160848
rect 321908 160790 324379 160792
rect 307569 160787 307635 160790
rect 324313 160787 324379 160790
rect 249149 160578 249215 160581
rect 248860 160576 249215 160578
rect 248860 160520 249154 160576
rect 249210 160520 249215 160576
rect 248860 160518 249215 160520
rect 249149 160515 249215 160518
rect 214005 160442 214071 160445
rect 307661 160442 307727 160445
rect 214005 160440 217212 160442
rect 214005 160384 214010 160440
rect 214066 160384 217212 160440
rect 214005 160382 217212 160384
rect 307661 160440 310132 160442
rect 307661 160384 307666 160440
rect 307722 160384 310132 160440
rect 307661 160382 310132 160384
rect 214005 160379 214071 160382
rect 307661 160379 307727 160382
rect 171174 160108 171180 160172
rect 171244 160170 171250 160172
rect 172329 160170 172395 160173
rect 251541 160170 251607 160173
rect 325601 160170 325667 160173
rect 171244 160168 172395 160170
rect 171244 160112 172334 160168
rect 172390 160112 172395 160168
rect 171244 160110 172395 160112
rect 248860 160168 251607 160170
rect 248860 160112 251546 160168
rect 251602 160112 251607 160168
rect 248860 160110 251607 160112
rect 321908 160168 325667 160170
rect 321908 160112 325606 160168
rect 325662 160112 325667 160168
rect 321908 160110 325667 160112
rect 171244 160108 171250 160110
rect 172329 160107 172395 160110
rect 251541 160107 251607 160110
rect 325601 160107 325667 160110
rect 307569 160034 307635 160037
rect 307569 160032 310132 160034
rect 307569 159976 307574 160032
rect 307630 159976 310132 160032
rect 307569 159974 310132 159976
rect 307569 159971 307635 159974
rect 572621 159898 572687 159901
rect 569940 159896 572687 159898
rect 569940 159840 572626 159896
rect 572682 159840 572687 159896
rect 569940 159838 572687 159840
rect 572621 159835 572687 159838
rect 217182 159218 217242 159732
rect 265014 159626 265020 159628
rect 248860 159566 265020 159626
rect 265014 159564 265020 159566
rect 265084 159564 265090 159628
rect 307477 159626 307543 159629
rect 307477 159624 310132 159626
rect 307477 159568 307482 159624
rect 307538 159568 310132 159624
rect 307477 159566 310132 159568
rect 307477 159563 307543 159566
rect 324313 159354 324379 159357
rect 321908 159352 324379 159354
rect 321908 159296 324318 159352
rect 324374 159296 324379 159352
rect 321908 159294 324379 159296
rect 324313 159291 324379 159294
rect 251449 159218 251515 159221
rect 200070 159158 217242 159218
rect 248860 159216 251515 159218
rect 248860 159160 251454 159216
rect 251510 159160 251515 159216
rect 248860 159158 251515 159160
rect 167678 158748 167684 158812
rect 167748 158810 167754 158812
rect 200070 158810 200130 159158
rect 251449 159155 251515 159158
rect 387057 159218 387123 159221
rect 387057 159216 390172 159218
rect 387057 159160 387062 159216
rect 387118 159160 390172 159216
rect 387057 159158 390172 159160
rect 387057 159155 387123 159158
rect 213913 159082 213979 159085
rect 307661 159082 307727 159085
rect 213913 159080 217212 159082
rect 213913 159024 213918 159080
rect 213974 159024 217212 159080
rect 213913 159022 217212 159024
rect 307661 159080 310132 159082
rect 307661 159024 307666 159080
rect 307722 159024 310132 159080
rect 307661 159022 310132 159024
rect 213913 159019 213979 159022
rect 307661 159019 307727 159022
rect 251357 158810 251423 158813
rect 167748 158750 200130 158810
rect 248860 158808 251423 158810
rect 248860 158752 251362 158808
rect 251418 158752 251423 158808
rect 248860 158750 251423 158752
rect 167748 158748 167754 158750
rect 251357 158747 251423 158750
rect 307661 158674 307727 158677
rect 307661 158672 310132 158674
rect 307661 158616 307666 158672
rect 307722 158616 310132 158672
rect 307661 158614 310132 158616
rect 307661 158611 307727 158614
rect 324313 158538 324379 158541
rect 321908 158536 324379 158538
rect 321908 158480 324318 158536
rect 324374 158480 324379 158536
rect 321908 158478 324379 158480
rect 324313 158475 324379 158478
rect 213913 158402 213979 158405
rect 213913 158400 217212 158402
rect 213913 158344 213918 158400
rect 213974 158344 217212 158400
rect 213913 158342 217212 158344
rect 213913 158339 213979 158342
rect 252461 158266 252527 158269
rect 248860 158264 252527 158266
rect 248860 158208 252466 158264
rect 252522 158208 252527 158264
rect 248860 158206 252527 158208
rect 252461 158203 252527 158206
rect 307477 158266 307543 158269
rect 307477 158264 310132 158266
rect 307477 158208 307482 158264
rect 307538 158208 310132 158264
rect 307477 158206 310132 158208
rect 307477 158203 307543 158206
rect 251909 157994 251975 157997
rect 262254 157994 262260 157996
rect 251909 157992 262260 157994
rect 251909 157936 251914 157992
rect 251970 157936 262260 157992
rect 251909 157934 262260 157936
rect 251909 157931 251975 157934
rect 262254 157932 262260 157934
rect 262324 157932 262330 157996
rect 251173 157858 251239 157861
rect 248860 157856 251239 157858
rect 248860 157800 251178 157856
rect 251234 157800 251239 157856
rect 248860 157798 251239 157800
rect 251173 157795 251239 157798
rect 307569 157858 307635 157861
rect 324405 157858 324471 157861
rect 307569 157856 310132 157858
rect 307569 157800 307574 157856
rect 307630 157800 310132 157856
rect 307569 157798 310132 157800
rect 321908 157856 324471 157858
rect 321908 157800 324410 157856
rect 324466 157800 324471 157856
rect 321908 157798 324471 157800
rect 307569 157795 307635 157798
rect 324405 157795 324471 157798
rect 214925 157722 214991 157725
rect 214925 157720 217212 157722
rect 214925 157664 214930 157720
rect 214986 157664 217212 157720
rect 214925 157662 217212 157664
rect 214925 157659 214991 157662
rect 307334 157388 307340 157452
rect 307404 157450 307410 157452
rect 307404 157390 310132 157450
rect 307404 157388 307410 157390
rect 252686 157314 252692 157316
rect 248860 157254 252692 157314
rect 252686 157252 252692 157254
rect 252756 157252 252762 157316
rect 213913 157178 213979 157181
rect 213913 157176 217212 157178
rect 213913 157120 213918 157176
rect 213974 157120 217212 157176
rect 213913 157118 217212 157120
rect 213913 157115 213979 157118
rect 306741 157042 306807 157045
rect 324313 157042 324379 157045
rect 306741 157040 310132 157042
rect 306741 156984 306746 157040
rect 306802 156984 310132 157040
rect 306741 156982 310132 156984
rect 321908 157040 324379 157042
rect 321908 156984 324318 157040
rect 324374 156984 324379 157040
rect 321908 156982 324379 156984
rect 306741 156979 306807 156982
rect 324313 156979 324379 156982
rect 251357 156906 251423 156909
rect 248860 156904 251423 156906
rect 248860 156848 251362 156904
rect 251418 156848 251423 156904
rect 248860 156846 251423 156848
rect 251357 156843 251423 156846
rect 307661 156634 307727 156637
rect 307661 156632 310132 156634
rect 307661 156576 307666 156632
rect 307722 156576 310132 156632
rect 307661 156574 310132 156576
rect 307661 156571 307727 156574
rect 214005 156498 214071 156501
rect 214005 156496 217212 156498
rect 214005 156440 214010 156496
rect 214066 156440 217212 156496
rect 214005 156438 217212 156440
rect 214005 156435 214071 156438
rect 251173 156362 251239 156365
rect 324405 156362 324471 156365
rect 248860 156360 251239 156362
rect 248860 156304 251178 156360
rect 251234 156304 251239 156360
rect 248860 156302 251239 156304
rect 321908 156360 324471 156362
rect 321908 156304 324410 156360
rect 324466 156304 324471 156360
rect 321908 156302 324471 156304
rect 251173 156299 251239 156302
rect 324405 156299 324471 156302
rect 306925 156226 306991 156229
rect 306925 156224 310132 156226
rect 306925 156168 306930 156224
rect 306986 156168 310132 156224
rect 306925 156166 310132 156168
rect 306925 156163 306991 156166
rect 569358 156093 569418 156468
rect 569309 156088 569418 156093
rect 569309 156032 569314 156088
rect 569370 156032 569418 156088
rect 569309 156030 569418 156032
rect 569309 156027 569375 156030
rect 252369 155954 252435 155957
rect 248860 155952 252435 155954
rect 248860 155896 252374 155952
rect 252430 155896 252435 155952
rect 248860 155894 252435 155896
rect 252369 155891 252435 155894
rect 388437 155954 388503 155957
rect 388437 155952 390172 155954
rect 388437 155896 388442 155952
rect 388498 155896 390172 155952
rect 388437 155894 390172 155896
rect 388437 155891 388503 155894
rect 213913 155818 213979 155821
rect 213913 155816 217212 155818
rect 213913 155760 213918 155816
rect 213974 155760 217212 155816
rect 213913 155758 217212 155760
rect 213913 155755 213979 155758
rect 307661 155682 307727 155685
rect 307661 155680 310132 155682
rect 307661 155624 307666 155680
rect 307722 155624 310132 155680
rect 307661 155622 310132 155624
rect 307661 155619 307727 155622
rect 324262 155546 324268 155548
rect 321908 155486 324268 155546
rect 324262 155484 324268 155486
rect 324332 155484 324338 155548
rect 252461 155410 252527 155413
rect 248860 155408 252527 155410
rect 248860 155352 252466 155408
rect 252522 155352 252527 155408
rect 248860 155350 252527 155352
rect 252461 155347 252527 155350
rect 307477 155274 307543 155277
rect 307477 155272 310132 155274
rect 307477 155216 307482 155272
rect 307538 155216 310132 155272
rect 307477 155214 310132 155216
rect 307477 155211 307543 155214
rect 166390 154532 166396 154596
rect 166460 154594 166466 154596
rect 217182 154594 217242 155108
rect 251817 155002 251883 155005
rect 248860 155000 251883 155002
rect 248860 154944 251822 155000
rect 251878 154944 251883 155000
rect 248860 154942 251883 154944
rect 251817 154939 251883 154942
rect 307293 154866 307359 154869
rect 307293 154864 310132 154866
rect 307293 154808 307298 154864
rect 307354 154808 310132 154864
rect 307293 154806 310132 154808
rect 307293 154803 307359 154806
rect 324313 154730 324379 154733
rect 321908 154728 324379 154730
rect 321908 154672 324318 154728
rect 324374 154672 324379 154728
rect 321908 154670 324379 154672
rect 324313 154667 324379 154670
rect 166460 154534 217242 154594
rect 166460 154532 166466 154534
rect 214005 154458 214071 154461
rect 252645 154458 252711 154461
rect 214005 154456 217212 154458
rect 214005 154400 214010 154456
rect 214066 154400 217212 154456
rect 214005 154398 217212 154400
rect 248860 154456 252711 154458
rect 248860 154400 252650 154456
rect 252706 154400 252711 154456
rect 248860 154398 252711 154400
rect 214005 154395 214071 154398
rect 252645 154395 252711 154398
rect 307569 154458 307635 154461
rect 307569 154456 310132 154458
rect 307569 154400 307574 154456
rect 307630 154400 310132 154456
rect 307569 154398 310132 154400
rect 307569 154395 307635 154398
rect 252461 154050 252527 154053
rect 248860 154048 252527 154050
rect 248860 153992 252466 154048
rect 252522 153992 252527 154048
rect 248860 153990 252527 153992
rect 252461 153987 252527 153990
rect 306557 154050 306623 154053
rect 324313 154050 324379 154053
rect 306557 154048 310132 154050
rect 306557 153992 306562 154048
rect 306618 153992 310132 154048
rect 306557 153990 310132 153992
rect 321908 154048 324379 154050
rect 321908 153992 324318 154048
rect 324374 153992 324379 154048
rect 321908 153990 324379 153992
rect 306557 153987 306623 153990
rect 324313 153987 324379 153990
rect 213913 153778 213979 153781
rect 213913 153776 217212 153778
rect 213913 153720 213918 153776
rect 213974 153720 217212 153776
rect 213913 153718 217212 153720
rect 213913 153715 213979 153718
rect 307017 153642 307083 153645
rect 307017 153640 310132 153642
rect 307017 153584 307022 153640
rect 307078 153584 310132 153640
rect 307017 153582 310132 153584
rect 307017 153579 307083 153582
rect 249793 153506 249859 153509
rect 248860 153504 249859 153506
rect 248860 153448 249798 153504
rect 249854 153448 249859 153504
rect 248860 153446 249859 153448
rect 249793 153443 249859 153446
rect 307661 153234 307727 153237
rect 324405 153234 324471 153237
rect 572621 153234 572687 153237
rect 307661 153232 310132 153234
rect 307661 153176 307666 153232
rect 307722 153176 310132 153232
rect 307661 153174 310132 153176
rect 321908 153232 324471 153234
rect 321908 153176 324410 153232
rect 324466 153176 324471 153232
rect 321908 153174 324471 153176
rect 569940 153232 572687 153234
rect 569940 153176 572626 153232
rect 572682 153176 572687 153232
rect 569940 153174 572687 153176
rect 307661 153171 307727 153174
rect 324405 153171 324471 153174
rect 572621 153171 572687 153174
rect 213913 153098 213979 153101
rect 252461 153098 252527 153101
rect 213913 153096 217212 153098
rect 213913 153040 213918 153096
rect 213974 153040 217212 153096
rect 213913 153038 217212 153040
rect 248860 153096 252527 153098
rect 248860 153040 252466 153096
rect 252522 153040 252527 153096
rect 248860 153038 252527 153040
rect 213913 153035 213979 153038
rect 252461 153035 252527 153038
rect 252369 152690 252435 152693
rect 248860 152688 252435 152690
rect 248860 152632 252374 152688
rect 252430 152632 252435 152688
rect 248860 152630 252435 152632
rect 252369 152627 252435 152630
rect 306557 152690 306623 152693
rect 581637 152690 581703 152693
rect 583520 152690 584960 152780
rect 306557 152688 310132 152690
rect 306557 152632 306562 152688
rect 306618 152632 310132 152688
rect 306557 152630 310132 152632
rect 581637 152688 584960 152690
rect 581637 152632 581642 152688
rect 581698 152632 584960 152688
rect 581637 152630 584960 152632
rect 306557 152627 306623 152630
rect 581637 152627 581703 152630
rect 214005 152554 214071 152557
rect 386873 152554 386939 152557
rect 214005 152552 217212 152554
rect 214005 152496 214010 152552
rect 214066 152496 217212 152552
rect 214005 152494 217212 152496
rect 386873 152552 390172 152554
rect 386873 152496 386878 152552
rect 386934 152496 390172 152552
rect 583520 152540 584960 152630
rect 386873 152494 390172 152496
rect 214005 152491 214071 152494
rect 386873 152491 386939 152494
rect 324957 152418 325023 152421
rect 321908 152416 325023 152418
rect 321908 152360 324962 152416
rect 325018 152360 325023 152416
rect 321908 152358 325023 152360
rect 324957 152355 325023 152358
rect 307569 152282 307635 152285
rect 307569 152280 310132 152282
rect 307569 152224 307574 152280
rect 307630 152224 310132 152280
rect 307569 152222 310132 152224
rect 307569 152219 307635 152222
rect 252277 152146 252343 152149
rect 248860 152144 252343 152146
rect 248860 152088 252282 152144
rect 252338 152088 252343 152144
rect 248860 152086 252343 152088
rect 252277 152083 252343 152086
rect 214649 151874 214715 151877
rect 307661 151874 307727 151877
rect 214649 151872 217212 151874
rect 214649 151816 214654 151872
rect 214710 151816 217212 151872
rect 214649 151814 217212 151816
rect 307661 151872 310132 151874
rect 307661 151816 307666 151872
rect 307722 151816 310132 151872
rect 307661 151814 310132 151816
rect 214649 151811 214715 151814
rect 307661 151811 307727 151814
rect 252461 151738 252527 151741
rect 324405 151738 324471 151741
rect 248860 151736 252527 151738
rect 248860 151680 252466 151736
rect 252522 151680 252527 151736
rect 248860 151678 252527 151680
rect 321908 151736 324471 151738
rect 321908 151680 324410 151736
rect 324466 151680 324471 151736
rect 321908 151678 324471 151680
rect 252461 151675 252527 151678
rect 324405 151675 324471 151678
rect 307477 151466 307543 151469
rect 307477 151464 310132 151466
rect 307477 151408 307482 151464
rect 307538 151408 310132 151464
rect 307477 151406 310132 151408
rect 307477 151403 307543 151406
rect 214005 151194 214071 151197
rect 249885 151194 249951 151197
rect 214005 151192 217212 151194
rect 214005 151136 214010 151192
rect 214066 151136 217212 151192
rect 214005 151134 217212 151136
rect 248860 151192 249951 151194
rect 248860 151136 249890 151192
rect 249946 151136 249951 151192
rect 248860 151134 249951 151136
rect 214005 151131 214071 151134
rect 249885 151131 249951 151134
rect 307569 151058 307635 151061
rect 307569 151056 310132 151058
rect 307569 151000 307574 151056
rect 307630 151000 310132 151056
rect 307569 150998 310132 151000
rect 307569 150995 307635 150998
rect 324313 150922 324379 150925
rect 321908 150920 324379 150922
rect 321908 150864 324318 150920
rect 324374 150864 324379 150920
rect 321908 150862 324379 150864
rect 324313 150859 324379 150862
rect 251909 150786 251975 150789
rect 248860 150784 251975 150786
rect 248860 150728 251914 150784
rect 251970 150728 251975 150784
rect 248860 150726 251975 150728
rect 251909 150723 251975 150726
rect 307661 150650 307727 150653
rect 307661 150648 310132 150650
rect 307661 150592 307666 150648
rect 307722 150592 310132 150648
rect 307661 150590 310132 150592
rect 307661 150587 307727 150590
rect 213913 150514 213979 150517
rect 572621 150514 572687 150517
rect 213913 150512 217212 150514
rect 213913 150456 213918 150512
rect 213974 150456 217212 150512
rect 213913 150454 217212 150456
rect 569940 150512 572687 150514
rect 569940 150456 572626 150512
rect 572682 150456 572687 150512
rect 569940 150454 572687 150456
rect 213913 150451 213979 150454
rect 572621 150451 572687 150454
rect 255446 150242 255452 150244
rect 248860 150182 255452 150242
rect 255446 150180 255452 150182
rect 255516 150180 255522 150244
rect 307150 150180 307156 150244
rect 307220 150242 307226 150244
rect 307220 150182 310132 150242
rect 307220 150180 307226 150182
rect 324313 150106 324379 150109
rect 321908 150104 324379 150106
rect 321908 150048 324318 150104
rect 324374 150048 324379 150104
rect 321908 150046 324379 150048
rect 324313 150043 324379 150046
rect 214005 149834 214071 149837
rect 251173 149834 251239 149837
rect 214005 149832 217212 149834
rect 214005 149776 214010 149832
rect 214066 149776 217212 149832
rect 214005 149774 217212 149776
rect 248860 149832 251239 149834
rect 248860 149776 251178 149832
rect 251234 149776 251239 149832
rect 248860 149774 251239 149776
rect 214005 149771 214071 149774
rect 251173 149771 251239 149774
rect 307477 149834 307543 149837
rect 307477 149832 310132 149834
rect 307477 149776 307482 149832
rect 307538 149776 310132 149832
rect 307477 149774 310132 149776
rect 307477 149771 307543 149774
rect 253197 149698 253263 149701
rect 306966 149698 306972 149700
rect 253197 149696 306972 149698
rect 253197 149640 253202 149696
rect 253258 149640 306972 149696
rect 253197 149638 306972 149640
rect 253197 149635 253263 149638
rect 306966 149636 306972 149638
rect 307036 149636 307042 149700
rect 324405 149426 324471 149429
rect 321908 149424 324471 149426
rect 321908 149368 324410 149424
rect 324466 149368 324471 149424
rect 321908 149366 324471 149368
rect 324405 149363 324471 149366
rect 251265 149290 251331 149293
rect 248860 149288 251331 149290
rect 248860 149232 251270 149288
rect 251326 149232 251331 149288
rect 248860 149230 251331 149232
rect 251265 149227 251331 149230
rect 306925 149290 306991 149293
rect 306925 149288 310132 149290
rect 306925 149232 306930 149288
rect 306986 149232 310132 149288
rect 306925 149230 310132 149232
rect 306925 149227 306991 149230
rect 213913 149154 213979 149157
rect 386597 149154 386663 149157
rect 213913 149152 217212 149154
rect 213913 149096 213918 149152
rect 213974 149096 217212 149152
rect 213913 149094 217212 149096
rect 386597 149152 390172 149154
rect 386597 149096 386602 149152
rect 386658 149096 390172 149152
rect 386597 149094 390172 149096
rect 213913 149091 213979 149094
rect 386597 149091 386663 149094
rect 251817 148882 251883 148885
rect 248860 148880 251883 148882
rect 248860 148824 251822 148880
rect 251878 148824 251883 148880
rect 248860 148822 251883 148824
rect 251817 148819 251883 148822
rect 307569 148882 307635 148885
rect 307569 148880 310132 148882
rect 307569 148824 307574 148880
rect 307630 148824 310132 148880
rect 307569 148822 310132 148824
rect 307569 148819 307635 148822
rect 322054 148746 322060 148748
rect 321878 148686 322060 148746
rect 321878 148610 321938 148686
rect 322054 148684 322060 148686
rect 322124 148684 322130 148748
rect 321540 148580 321938 148610
rect 321510 148550 321908 148580
rect 213913 148474 213979 148477
rect 307477 148474 307543 148477
rect 213913 148472 217212 148474
rect 213913 148416 213918 148472
rect 213974 148416 217212 148472
rect 213913 148414 217212 148416
rect 307477 148472 310132 148474
rect 307477 148416 307482 148472
rect 307538 148416 310132 148472
rect 307477 148414 310132 148416
rect 213913 148411 213979 148414
rect 307477 148411 307543 148414
rect 252461 148338 252527 148341
rect 248860 148336 252527 148338
rect 248860 148280 252466 148336
rect 252522 148280 252527 148336
rect 248860 148278 252527 148280
rect 252461 148275 252527 148278
rect 251950 148140 251956 148204
rect 252020 148202 252026 148204
rect 262949 148202 263015 148205
rect 252020 148200 263015 148202
rect 252020 148144 262954 148200
rect 263010 148144 263015 148200
rect 252020 148142 263015 148144
rect 252020 148140 252026 148142
rect 262949 148139 263015 148142
rect 307661 148066 307727 148069
rect 321510 148068 321570 148550
rect 321829 148338 321895 148341
rect 321829 148336 321938 148338
rect 321829 148280 321834 148336
rect 321890 148280 321938 148336
rect 321829 148275 321938 148280
rect 307661 148064 310132 148066
rect 307661 148008 307666 148064
rect 307722 148008 310132 148064
rect 307661 148006 310132 148008
rect 307661 148003 307727 148006
rect 321502 148004 321508 148068
rect 321572 148004 321578 148068
rect 214097 147930 214163 147933
rect 251214 147930 251220 147932
rect 214097 147928 217212 147930
rect 214097 147872 214102 147928
rect 214158 147872 217212 147928
rect 214097 147870 217212 147872
rect 248860 147870 251220 147930
rect 214097 147867 214163 147870
rect 251214 147868 251220 147870
rect 251284 147868 251290 147932
rect 321878 147794 321938 148275
rect 322841 147794 322907 147797
rect 321878 147792 322907 147794
rect 321878 147764 322846 147792
rect 321908 147736 322846 147764
rect 322902 147736 322907 147792
rect 321908 147734 322907 147736
rect 322841 147731 322907 147734
rect 307385 147658 307451 147661
rect 307385 147656 310132 147658
rect 307385 147600 307390 147656
rect 307446 147600 310132 147656
rect 307385 147598 310132 147600
rect 307385 147595 307451 147598
rect 252461 147522 252527 147525
rect 248860 147520 252527 147522
rect 248860 147464 252466 147520
rect 252522 147464 252527 147520
rect 248860 147462 252527 147464
rect 252461 147459 252527 147462
rect 214005 147250 214071 147253
rect 307477 147250 307543 147253
rect 214005 147248 217212 147250
rect 214005 147192 214010 147248
rect 214066 147192 217212 147248
rect 214005 147190 217212 147192
rect 307477 147248 310132 147250
rect 307477 147192 307482 147248
rect 307538 147192 310132 147248
rect 307477 147190 310132 147192
rect 214005 147187 214071 147190
rect 307477 147187 307543 147190
rect 324313 147114 324379 147117
rect 571701 147114 571767 147117
rect 321908 147112 324379 147114
rect 321908 147056 324318 147112
rect 324374 147056 324379 147112
rect 321908 147054 324379 147056
rect 569940 147112 571767 147114
rect 569940 147056 571706 147112
rect 571762 147056 571767 147112
rect 569940 147054 571767 147056
rect 324313 147051 324379 147054
rect 571701 147051 571767 147054
rect 251725 146978 251791 146981
rect 248860 146976 251791 146978
rect 248860 146920 251730 146976
rect 251786 146920 251791 146976
rect 248860 146918 251791 146920
rect 251725 146915 251791 146918
rect 307569 146842 307635 146845
rect 307569 146840 310132 146842
rect 307569 146784 307574 146840
rect 307630 146784 310132 146840
rect 307569 146782 310132 146784
rect 307569 146779 307635 146782
rect 213913 146570 213979 146573
rect 252369 146570 252435 146573
rect 213913 146568 217212 146570
rect 213913 146512 213918 146568
rect 213974 146512 217212 146568
rect 213913 146510 217212 146512
rect 248860 146568 252435 146570
rect 248860 146512 252374 146568
rect 252430 146512 252435 146568
rect 248860 146510 252435 146512
rect 213913 146507 213979 146510
rect 252369 146507 252435 146510
rect 307661 146434 307727 146437
rect 307661 146432 310132 146434
rect 307661 146376 307666 146432
rect 307722 146376 310132 146432
rect 307661 146374 310132 146376
rect 307661 146371 307727 146374
rect 251766 146236 251772 146300
rect 251836 146298 251842 146300
rect 254117 146298 254183 146301
rect 251836 146296 254183 146298
rect 251836 146240 254122 146296
rect 254178 146240 254183 146296
rect 251836 146238 254183 146240
rect 251836 146236 251842 146238
rect 254117 146235 254183 146238
rect 255814 146236 255820 146300
rect 255884 146298 255890 146300
rect 256233 146298 256299 146301
rect 255884 146296 256299 146298
rect 255884 146240 256238 146296
rect 256294 146240 256299 146296
rect 255884 146238 256299 146240
rect 255884 146236 255890 146238
rect 256233 146235 256299 146238
rect 252093 146026 252159 146029
rect 248860 146024 252159 146026
rect 248860 145968 252098 146024
rect 252154 145968 252159 146024
rect 248860 145966 252159 145968
rect 252093 145963 252159 145966
rect 214005 145890 214071 145893
rect 306557 145890 306623 145893
rect 214005 145888 217212 145890
rect 214005 145832 214010 145888
rect 214066 145832 217212 145888
rect 214005 145830 217212 145832
rect 306557 145888 310132 145890
rect 306557 145832 306562 145888
rect 306618 145832 310132 145888
rect 306557 145830 310132 145832
rect 214005 145827 214071 145830
rect 306557 145827 306623 145830
rect 266302 145618 266308 145620
rect 248860 145558 266308 145618
rect 266302 145556 266308 145558
rect 266372 145556 266378 145620
rect 287973 145618 288039 145621
rect 307334 145618 307340 145620
rect 287973 145616 307340 145618
rect 287973 145560 287978 145616
rect 288034 145560 307340 145616
rect 287973 145558 307340 145560
rect 287973 145555 288039 145558
rect 307334 145556 307340 145558
rect 307404 145556 307410 145620
rect 321878 145618 321938 146268
rect 328494 145618 328500 145620
rect 321878 145558 328500 145618
rect 328494 145556 328500 145558
rect 328564 145556 328570 145620
rect 386597 145618 386663 145621
rect 386597 145616 390172 145618
rect 386597 145560 386602 145616
rect 386658 145560 390172 145616
rect 386597 145558 390172 145560
rect 386597 145555 386663 145558
rect 305729 145482 305795 145485
rect 324313 145482 324379 145485
rect 305729 145480 310132 145482
rect 305729 145424 305734 145480
rect 305790 145424 310132 145480
rect 305729 145422 310132 145424
rect 321908 145480 324379 145482
rect 321908 145424 324318 145480
rect 324374 145424 324379 145480
rect 321908 145422 324379 145424
rect 305729 145419 305795 145422
rect 324313 145419 324379 145422
rect 213913 145210 213979 145213
rect 213913 145208 217212 145210
rect 213913 145152 213918 145208
rect 213974 145152 217212 145208
rect 213913 145150 217212 145152
rect 213913 145147 213979 145150
rect 252277 145074 252343 145077
rect 248860 145072 252343 145074
rect 248860 145016 252282 145072
rect 252338 145016 252343 145072
rect 248860 145014 252343 145016
rect 252277 145011 252343 145014
rect 306925 145074 306991 145077
rect 306925 145072 310132 145074
rect 306925 145016 306930 145072
rect 306986 145016 310132 145072
rect 306925 145014 310132 145016
rect 306925 145011 306991 145014
rect 324313 144802 324379 144805
rect 321908 144800 324379 144802
rect 321908 144744 324318 144800
rect 324374 144744 324379 144800
rect 321908 144742 324379 144744
rect 324313 144739 324379 144742
rect 251541 144666 251607 144669
rect 248860 144664 251607 144666
rect 248860 144608 251546 144664
rect 251602 144608 251607 144664
rect 248860 144606 251607 144608
rect 251541 144603 251607 144606
rect 306925 144666 306991 144669
rect 306925 144664 310132 144666
rect 306925 144608 306930 144664
rect 306986 144608 310132 144664
rect 306925 144606 310132 144608
rect 306925 144603 306991 144606
rect 213913 144530 213979 144533
rect 213913 144528 217212 144530
rect 213913 144472 213918 144528
rect 213974 144472 217212 144528
rect 213913 144470 217212 144472
rect 213913 144467 213979 144470
rect 306557 144258 306623 144261
rect 306557 144256 310132 144258
rect 306557 144200 306562 144256
rect 306618 144200 310132 144256
rect 306557 144198 310132 144200
rect 306557 144195 306623 144198
rect 251909 144122 251975 144125
rect 248860 144120 251975 144122
rect 248860 144064 251914 144120
rect 251970 144064 251975 144120
rect 248860 144062 251975 144064
rect 251909 144059 251975 144062
rect 324405 143986 324471 143989
rect 321908 143984 324471 143986
rect 321908 143928 324410 143984
rect 324466 143928 324471 143984
rect 321908 143926 324471 143928
rect 324405 143923 324471 143926
rect 214649 143850 214715 143853
rect 307661 143850 307727 143853
rect 214649 143848 217212 143850
rect 214649 143792 214654 143848
rect 214710 143792 217212 143848
rect 214649 143790 217212 143792
rect 307661 143848 310132 143850
rect 307661 143792 307666 143848
rect 307722 143792 310132 143848
rect 307661 143790 310132 143792
rect 214649 143787 214715 143790
rect 307661 143787 307727 143790
rect 252461 143714 252527 143717
rect 248860 143712 252527 143714
rect 248860 143656 252466 143712
rect 252522 143656 252527 143712
rect 248860 143654 252527 143656
rect 252461 143651 252527 143654
rect 572621 143578 572687 143581
rect 569940 143576 572687 143578
rect 569940 143520 572626 143576
rect 572682 143520 572687 143576
rect 569940 143518 572687 143520
rect 572621 143515 572687 143518
rect 307661 143442 307727 143445
rect 307661 143440 310132 143442
rect 307661 143384 307666 143440
rect 307722 143384 310132 143440
rect 307661 143382 310132 143384
rect 307661 143379 307727 143382
rect 213913 143306 213979 143309
rect 213913 143304 217212 143306
rect 213913 143248 213918 143304
rect 213974 143248 217212 143304
rect 213913 143246 217212 143248
rect 213913 143243 213979 143246
rect 250621 143170 250687 143173
rect 324313 143170 324379 143173
rect 248860 143168 250687 143170
rect 248860 143112 250626 143168
rect 250682 143112 250687 143168
rect 248860 143110 250687 143112
rect 321908 143168 324379 143170
rect 321908 143112 324318 143168
rect 324374 143112 324379 143168
rect 321908 143110 324379 143112
rect 250621 143107 250687 143110
rect 324313 143107 324379 143110
rect 307477 143034 307543 143037
rect 307477 143032 310132 143034
rect 307477 142976 307482 143032
rect 307538 142976 310132 143032
rect 307477 142974 310132 142976
rect 307477 142971 307543 142974
rect 387609 142898 387675 142901
rect 387609 142896 390172 142898
rect 387609 142840 387614 142896
rect 387670 142840 390172 142896
rect 387609 142838 390172 142840
rect 387609 142835 387675 142838
rect 252461 142762 252527 142765
rect 248860 142760 252527 142762
rect 248860 142704 252466 142760
rect 252522 142704 252527 142760
rect 248860 142702 252527 142704
rect 252461 142699 252527 142702
rect 214557 142626 214623 142629
rect 251081 142626 251147 142629
rect 259678 142626 259684 142628
rect 214557 142624 217212 142626
rect 214557 142568 214562 142624
rect 214618 142568 217212 142624
rect 214557 142566 217212 142568
rect 251081 142624 259684 142626
rect 251081 142568 251086 142624
rect 251142 142568 259684 142624
rect 251081 142566 259684 142568
rect 214557 142563 214623 142566
rect 251081 142563 251147 142566
rect 259678 142564 259684 142566
rect 259748 142564 259754 142628
rect 306741 142490 306807 142493
rect 324405 142490 324471 142493
rect 306741 142488 310132 142490
rect 306741 142432 306746 142488
rect 306802 142432 310132 142488
rect 306741 142430 310132 142432
rect 321908 142488 324471 142490
rect 321908 142432 324410 142488
rect 324466 142432 324471 142488
rect 321908 142430 324471 142432
rect 306741 142427 306807 142430
rect 324405 142427 324471 142430
rect 252369 142218 252435 142221
rect 248860 142216 252435 142218
rect 248860 142160 252374 142216
rect 252430 142160 252435 142216
rect 248860 142158 252435 142160
rect 252369 142155 252435 142158
rect 307702 142020 307708 142084
rect 307772 142082 307778 142084
rect 307772 142022 310132 142082
rect 307772 142020 307778 142022
rect 214005 141946 214071 141949
rect 214005 141944 217212 141946
rect 214005 141888 214010 141944
rect 214066 141888 217212 141944
rect 214005 141886 217212 141888
rect 214005 141883 214071 141886
rect 256734 141810 256740 141812
rect 248860 141750 256740 141810
rect 256734 141748 256740 141750
rect 256804 141748 256810 141812
rect 307385 141674 307451 141677
rect 324313 141674 324379 141677
rect 307385 141672 310132 141674
rect 307385 141616 307390 141672
rect 307446 141616 310132 141672
rect 307385 141614 310132 141616
rect 321908 141672 324379 141674
rect 321908 141616 324318 141672
rect 324374 141616 324379 141672
rect 321908 141614 324379 141616
rect 307385 141611 307451 141614
rect 324313 141611 324379 141614
rect 252461 141402 252527 141405
rect 248860 141400 252527 141402
rect 248860 141344 252466 141400
rect 252522 141344 252527 141400
rect 248860 141342 252527 141344
rect 252461 141339 252527 141342
rect 213913 141266 213979 141269
rect 307661 141266 307727 141269
rect 213913 141264 217212 141266
rect 213913 141208 213918 141264
rect 213974 141208 217212 141264
rect 213913 141206 217212 141208
rect 307661 141264 310132 141266
rect 307661 141208 307666 141264
rect 307722 141208 310132 141264
rect 307661 141206 310132 141208
rect 213913 141203 213979 141206
rect 307661 141203 307727 141206
rect 255262 140858 255268 140860
rect 248860 140798 255268 140858
rect 255262 140796 255268 140798
rect 255332 140796 255338 140860
rect 306005 140858 306071 140861
rect 324405 140858 324471 140861
rect 306005 140856 310132 140858
rect 306005 140800 306010 140856
rect 306066 140800 310132 140856
rect 306005 140798 310132 140800
rect 321908 140856 324471 140858
rect 321908 140800 324410 140856
rect 324466 140800 324471 140856
rect 321908 140798 324471 140800
rect 306005 140795 306071 140798
rect 324405 140795 324471 140798
rect 213913 140586 213979 140589
rect 213913 140584 217212 140586
rect 213913 140528 213918 140584
rect 213974 140528 217212 140584
rect 213913 140526 217212 140528
rect 213913 140523 213979 140526
rect 252093 140450 252159 140453
rect 248860 140448 252159 140450
rect 248860 140392 252098 140448
rect 252154 140392 252159 140448
rect 248860 140390 252159 140392
rect 252093 140387 252159 140390
rect 307569 140450 307635 140453
rect 307569 140448 310132 140450
rect 307569 140392 307574 140448
rect 307630 140392 310132 140448
rect 307569 140390 310132 140392
rect 307569 140387 307635 140390
rect 324313 140178 324379 140181
rect 572621 140178 572687 140181
rect 321908 140176 324379 140178
rect 321908 140120 324318 140176
rect 324374 140120 324379 140176
rect 321908 140118 324379 140120
rect 569940 140176 572687 140178
rect 569940 140120 572626 140176
rect 572682 140120 572687 140176
rect 569940 140118 572687 140120
rect 324313 140115 324379 140118
rect 572621 140115 572687 140118
rect 297725 140042 297791 140045
rect 307702 140042 307708 140044
rect 297725 140040 307708 140042
rect 297725 139984 297730 140040
rect 297786 139984 307708 140040
rect 297725 139982 307708 139984
rect 297725 139979 297791 139982
rect 307702 139980 307708 139982
rect 307772 139980 307778 140044
rect 308262 139982 310132 140042
rect 214649 139906 214715 139909
rect 251725 139906 251791 139909
rect 214649 139904 217212 139906
rect 214649 139848 214654 139904
rect 214710 139848 217212 139904
rect 214649 139846 217212 139848
rect 248860 139904 251791 139906
rect 248860 139848 251730 139904
rect 251786 139848 251791 139904
rect 248860 139846 251791 139848
rect 214649 139843 214715 139846
rect 251725 139843 251791 139846
rect 305494 139708 305500 139772
rect 305564 139770 305570 139772
rect 308262 139770 308322 139982
rect 305564 139710 308322 139770
rect 305564 139708 305570 139710
rect 307661 139634 307727 139637
rect 307661 139632 310132 139634
rect 307661 139576 307666 139632
rect 307722 139576 310132 139632
rect 307661 139574 310132 139576
rect 307661 139571 307727 139574
rect 251725 139498 251791 139501
rect 248860 139496 251791 139498
rect 248860 139440 251730 139496
rect 251786 139440 251791 139496
rect 248860 139438 251791 139440
rect 251725 139435 251791 139438
rect 387149 139498 387215 139501
rect 387149 139496 390172 139498
rect 387149 139440 387154 139496
rect 387210 139440 390172 139496
rect 387149 139438 390172 139440
rect 387149 139435 387215 139438
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 214005 139226 214071 139229
rect 214005 139224 217212 139226
rect 214005 139168 214010 139224
rect 214066 139168 217212 139224
rect 214005 139166 217212 139168
rect 214005 139163 214071 139166
rect 306925 139090 306991 139093
rect 321737 139090 321803 139093
rect 306925 139088 310132 139090
rect 306925 139032 306930 139088
rect 306986 139032 310132 139088
rect 306925 139030 310132 139032
rect 321694 139088 321803 139090
rect 321694 139032 321742 139088
rect 321798 139032 321803 139088
rect 306925 139027 306991 139030
rect 321694 139027 321803 139032
rect 248860 138894 253122 138954
rect 213913 138682 213979 138685
rect 213913 138680 217212 138682
rect 213913 138624 213918 138680
rect 213974 138624 217212 138680
rect 213913 138622 217212 138624
rect 213913 138619 213979 138622
rect 251357 138546 251423 138549
rect 248860 138544 251423 138546
rect 248860 138488 251362 138544
rect 251418 138488 251423 138544
rect 248860 138486 251423 138488
rect 251357 138483 251423 138486
rect 253062 138274 253122 138894
rect 296670 138622 310132 138682
rect 253238 138348 253244 138412
rect 253308 138410 253314 138412
rect 296670 138410 296730 138622
rect 321694 138546 321754 139027
rect 321878 138682 321938 139332
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect 332542 138682 332548 138684
rect 321878 138622 332548 138682
rect 332542 138620 332548 138622
rect 332612 138620 332618 138684
rect 322841 138546 322907 138549
rect 321694 138544 322907 138546
rect 321694 138516 322846 138544
rect 321724 138488 322846 138516
rect 322902 138488 322907 138544
rect 321724 138486 322907 138488
rect 322841 138483 322907 138486
rect 253308 138350 296730 138410
rect 253308 138348 253314 138350
rect 259494 138274 259500 138276
rect 253062 138214 259500 138274
rect 259494 138212 259500 138214
rect 259564 138212 259570 138276
rect 307201 138274 307267 138277
rect 307201 138272 310132 138274
rect 307201 138216 307206 138272
rect 307262 138216 310132 138272
rect 307201 138214 310132 138216
rect 307201 138211 307267 138214
rect 263542 138002 263548 138004
rect 217182 137458 217242 137972
rect 248860 137942 263548 138002
rect 263542 137940 263548 137942
rect 263612 137940 263618 138004
rect 306925 137866 306991 137869
rect 324313 137866 324379 137869
rect 306925 137864 310132 137866
rect 306925 137808 306930 137864
rect 306986 137808 310132 137864
rect 306925 137806 310132 137808
rect 321908 137864 324379 137866
rect 321908 137808 324318 137864
rect 324374 137808 324379 137864
rect 321908 137806 324379 137808
rect 306925 137803 306991 137806
rect 324313 137803 324379 137806
rect 252093 137594 252159 137597
rect 248860 137592 252159 137594
rect 248860 137536 252098 137592
rect 252154 137536 252159 137592
rect 248860 137534 252159 137536
rect 252093 137531 252159 137534
rect 200070 137398 217242 137458
rect 307661 137458 307727 137461
rect 307661 137456 310132 137458
rect 307661 137400 307666 137456
rect 307722 137400 310132 137456
rect 307661 137398 310132 137400
rect 171910 136852 171916 136916
rect 171980 136914 171986 136916
rect 200070 136914 200130 137398
rect 307661 137395 307727 137398
rect 214649 137322 214715 137325
rect 214649 137320 217212 137322
rect 214649 137264 214654 137320
rect 214710 137264 217212 137320
rect 214649 137262 217212 137264
rect 214649 137259 214715 137262
rect 252461 137050 252527 137053
rect 248860 137048 252527 137050
rect 248860 136992 252466 137048
rect 252522 136992 252527 137048
rect 248860 136990 252527 136992
rect 252461 136987 252527 136990
rect 307293 137050 307359 137053
rect 324405 137050 324471 137053
rect 307293 137048 310132 137050
rect 307293 136992 307298 137048
rect 307354 136992 310132 137048
rect 307293 136990 310132 136992
rect 321908 137048 324471 137050
rect 321908 136992 324410 137048
rect 324466 136992 324471 137048
rect 321908 136990 324471 136992
rect 307293 136987 307359 136990
rect 324405 136987 324471 136990
rect 572621 136914 572687 136917
rect 171980 136854 200130 136914
rect 569940 136912 572687 136914
rect 569940 136856 572626 136912
rect 572682 136856 572687 136912
rect 569940 136854 572687 136856
rect 171980 136852 171986 136854
rect 572621 136851 572687 136854
rect 214741 136642 214807 136645
rect 260966 136642 260972 136644
rect 214741 136640 217212 136642
rect 214741 136584 214746 136640
rect 214802 136584 217212 136640
rect 214741 136582 217212 136584
rect 248860 136582 260972 136642
rect 214741 136579 214807 136582
rect 260966 136580 260972 136582
rect 261036 136580 261042 136644
rect 306925 136642 306991 136645
rect 306925 136640 310132 136642
rect 306925 136584 306930 136640
rect 306986 136584 310132 136640
rect 306925 136582 310132 136584
rect 306925 136579 306991 136582
rect 324313 136370 324379 136373
rect 321908 136368 324379 136370
rect 321908 136312 324318 136368
rect 324374 136312 324379 136368
rect 321908 136310 324379 136312
rect 324313 136307 324379 136310
rect 252093 136234 252159 136237
rect 248860 136232 252159 136234
rect 248860 136176 252098 136232
rect 252154 136176 252159 136232
rect 248860 136174 252159 136176
rect 252093 136171 252159 136174
rect 307477 136234 307543 136237
rect 307477 136232 310132 136234
rect 307477 136176 307482 136232
rect 307538 136176 310132 136232
rect 307477 136174 310132 136176
rect 307477 136171 307543 136174
rect 386689 136098 386755 136101
rect 386689 136096 390172 136098
rect 386689 136040 386694 136096
rect 386750 136040 390172 136096
rect 386689 136038 390172 136040
rect 386689 136035 386755 136038
rect 214005 135962 214071 135965
rect 214005 135960 217212 135962
rect 214005 135904 214010 135960
rect 214066 135904 217212 135960
rect 214005 135902 217212 135904
rect 214005 135899 214071 135902
rect 251725 135690 251791 135693
rect 248860 135688 251791 135690
rect 248860 135632 251730 135688
rect 251786 135632 251791 135688
rect 248860 135630 251791 135632
rect 251725 135627 251791 135630
rect 307569 135690 307635 135693
rect 307569 135688 310132 135690
rect 307569 135632 307574 135688
rect 307630 135632 310132 135688
rect 307569 135630 310132 135632
rect 307569 135627 307635 135630
rect 324405 135554 324471 135557
rect 321908 135552 324471 135554
rect 321908 135496 324410 135552
rect 324466 135496 324471 135552
rect 321908 135494 324471 135496
rect 324405 135491 324471 135494
rect 213913 135282 213979 135285
rect 252369 135282 252435 135285
rect 213913 135280 217212 135282
rect 213913 135224 213918 135280
rect 213974 135224 217212 135280
rect 213913 135222 217212 135224
rect 248860 135280 252435 135282
rect 248860 135224 252374 135280
rect 252430 135224 252435 135280
rect 248860 135222 252435 135224
rect 213913 135219 213979 135222
rect 252369 135219 252435 135222
rect 307661 135282 307727 135285
rect 307661 135280 310132 135282
rect 307661 135224 307666 135280
rect 307722 135224 310132 135280
rect 307661 135222 310132 135224
rect 307661 135219 307727 135222
rect 306741 134874 306807 134877
rect 306741 134872 310132 134874
rect 306741 134816 306746 134872
rect 306802 134816 310132 134872
rect 306741 134814 310132 134816
rect 306741 134811 306807 134814
rect 252461 134738 252527 134741
rect 324313 134738 324379 134741
rect 248860 134736 252527 134738
rect 248860 134680 252466 134736
rect 252522 134680 252527 134736
rect 248860 134678 252527 134680
rect 321908 134736 324379 134738
rect 321908 134680 324318 134736
rect 324374 134680 324379 134736
rect 321908 134678 324379 134680
rect 252461 134675 252527 134678
rect 324313 134675 324379 134678
rect 213913 134602 213979 134605
rect 213913 134600 217212 134602
rect 213913 134544 213918 134600
rect 213974 134544 217212 134600
rect 213913 134542 217212 134544
rect 213913 134539 213979 134542
rect 283925 134466 283991 134469
rect 307150 134466 307156 134468
rect 283925 134464 307156 134466
rect 283925 134408 283930 134464
rect 283986 134408 307156 134464
rect 283925 134406 307156 134408
rect 283925 134403 283991 134406
rect 307150 134404 307156 134406
rect 307220 134404 307226 134468
rect 307661 134466 307727 134469
rect 307661 134464 310132 134466
rect 307661 134408 307666 134464
rect 307722 134408 310132 134464
rect 307661 134406 310132 134408
rect 307661 134403 307727 134406
rect 252277 134330 252343 134333
rect 248860 134328 252343 134330
rect 248860 134272 252282 134328
rect 252338 134272 252343 134328
rect 248860 134270 252343 134272
rect 252277 134267 252343 134270
rect 306966 133996 306972 134060
rect 307036 134058 307042 134060
rect 324405 134058 324471 134061
rect 307036 133998 310132 134058
rect 321908 134056 324471 134058
rect 321908 134000 324410 134056
rect 324466 134000 324471 134056
rect 321908 133998 324471 134000
rect 307036 133996 307042 133998
rect 324405 133995 324471 133998
rect 166390 133860 166396 133924
rect 166460 133922 166466 133924
rect 166460 133862 217212 133922
rect 166460 133860 166466 133862
rect 252461 133786 252527 133789
rect 248860 133784 252527 133786
rect 248860 133728 252466 133784
rect 252522 133728 252527 133784
rect 248860 133726 252527 133728
rect 252461 133723 252527 133726
rect 306925 133650 306991 133653
rect 306925 133648 310132 133650
rect 306925 133592 306930 133648
rect 306986 133592 310132 133648
rect 306925 133590 310132 133592
rect 306925 133587 306991 133590
rect 213913 133378 213979 133381
rect 252369 133378 252435 133381
rect 572713 133378 572779 133381
rect 213913 133376 217212 133378
rect 213913 133320 213918 133376
rect 213974 133320 217212 133376
rect 213913 133318 217212 133320
rect 248860 133376 252435 133378
rect 248860 133320 252374 133376
rect 252430 133320 252435 133376
rect 248860 133318 252435 133320
rect 569940 133376 572779 133378
rect 569940 133320 572718 133376
rect 572774 133320 572779 133376
rect 569940 133318 572779 133320
rect 213913 133315 213979 133318
rect 252369 133315 252435 133318
rect 572713 133315 572779 133318
rect 307477 133242 307543 133245
rect 324313 133242 324379 133245
rect 307477 133240 310132 133242
rect 307477 133184 307482 133240
rect 307538 133184 310132 133240
rect 307477 133182 310132 133184
rect 321908 133240 324379 133242
rect 321908 133184 324318 133240
rect 324374 133184 324379 133240
rect 321908 133182 324379 133184
rect 307477 133179 307543 133182
rect 324313 133179 324379 133182
rect 251725 132834 251791 132837
rect 248860 132832 251791 132834
rect 248860 132776 251730 132832
rect 251786 132776 251791 132832
rect 248860 132774 251791 132776
rect 251725 132771 251791 132774
rect 389081 132834 389147 132837
rect 389081 132832 390172 132834
rect 389081 132776 389086 132832
rect 389142 132776 390172 132832
rect 389081 132774 390172 132776
rect 389081 132771 389147 132774
rect 214414 132636 214420 132700
rect 214484 132698 214490 132700
rect 214484 132638 217212 132698
rect 214484 132636 214490 132638
rect 299974 132636 299980 132700
rect 300044 132698 300050 132700
rect 300044 132638 310132 132698
rect 300044 132636 300050 132638
rect 252461 132426 252527 132429
rect 324313 132426 324379 132429
rect 248860 132424 252527 132426
rect 248860 132368 252466 132424
rect 252522 132368 252527 132424
rect 248860 132366 252527 132368
rect 321908 132424 324379 132426
rect 321908 132368 324318 132424
rect 324374 132368 324379 132424
rect 321908 132366 324379 132368
rect 252461 132363 252527 132366
rect 324313 132363 324379 132366
rect 307477 132290 307543 132293
rect 307477 132288 310132 132290
rect 307477 132232 307482 132288
rect 307538 132232 310132 132288
rect 307477 132230 310132 132232
rect 307477 132227 307543 132230
rect 166206 131412 166212 131476
rect 166276 131474 166282 131476
rect 217182 131474 217242 131988
rect 252461 131882 252527 131885
rect 248860 131880 252527 131882
rect 248860 131824 252466 131880
rect 252522 131824 252527 131880
rect 248860 131822 252527 131824
rect 252461 131819 252527 131822
rect 307569 131882 307635 131885
rect 307569 131880 310132 131882
rect 307569 131824 307574 131880
rect 307630 131824 310132 131880
rect 307569 131822 310132 131824
rect 307569 131819 307635 131822
rect 324405 131746 324471 131749
rect 321908 131744 324471 131746
rect 321908 131688 324410 131744
rect 324466 131688 324471 131744
rect 321908 131686 324471 131688
rect 324405 131683 324471 131686
rect 251909 131474 251975 131477
rect 166276 131414 217242 131474
rect 248860 131472 251975 131474
rect 248860 131416 251914 131472
rect 251970 131416 251975 131472
rect 248860 131414 251975 131416
rect 166276 131412 166282 131414
rect 251909 131411 251975 131414
rect 307661 131474 307727 131477
rect 307661 131472 310132 131474
rect 307661 131416 307666 131472
rect 307722 131416 310132 131472
rect 307661 131414 310132 131416
rect 307661 131411 307727 131414
rect 213913 131338 213979 131341
rect 213913 131336 217212 131338
rect 213913 131280 213918 131336
rect 213974 131280 217212 131336
rect 213913 131278 217212 131280
rect 213913 131275 213979 131278
rect 306741 131066 306807 131069
rect 306741 131064 310132 131066
rect 306741 131008 306746 131064
rect 306802 131008 310132 131064
rect 306741 131006 310132 131008
rect 306741 131003 306807 131006
rect 252461 130930 252527 130933
rect 324313 130930 324379 130933
rect 248860 130928 252527 130930
rect 248860 130872 252466 130928
rect 252522 130872 252527 130928
rect 248860 130870 252527 130872
rect 321908 130928 324379 130930
rect 321908 130872 324318 130928
rect 324374 130872 324379 130928
rect 321908 130870 324379 130872
rect 252461 130867 252527 130870
rect 324313 130867 324379 130870
rect 307569 130658 307635 130661
rect 307569 130656 310132 130658
rect 170254 130052 170260 130116
rect 170324 130114 170330 130116
rect 217182 130114 217242 130628
rect 307569 130600 307574 130656
rect 307630 130600 310132 130656
rect 307569 130598 310132 130600
rect 307569 130595 307635 130598
rect 252369 130522 252435 130525
rect 248860 130520 252435 130522
rect 248860 130464 252374 130520
rect 252430 130464 252435 130520
rect 248860 130462 252435 130464
rect 252369 130459 252435 130462
rect 307661 130250 307727 130253
rect 307661 130248 310132 130250
rect 307661 130192 307666 130248
rect 307722 130192 310132 130248
rect 307661 130190 310132 130192
rect 307661 130187 307727 130190
rect 252185 130114 252251 130117
rect 324405 130114 324471 130117
rect 572621 130114 572687 130117
rect 170324 130054 217242 130114
rect 248860 130112 252251 130114
rect 248860 130056 252190 130112
rect 252246 130056 252251 130112
rect 248860 130054 252251 130056
rect 321908 130112 324471 130114
rect 321908 130056 324410 130112
rect 324466 130056 324471 130112
rect 321908 130054 324471 130056
rect 569940 130112 572687 130114
rect 569940 130056 572626 130112
rect 572682 130056 572687 130112
rect 569940 130054 572687 130056
rect 170324 130052 170330 130054
rect 252185 130051 252251 130054
rect 324405 130051 324471 130054
rect 572621 130051 572687 130054
rect 171726 129916 171732 129980
rect 171796 129978 171802 129980
rect 171796 129918 217212 129978
rect 171796 129916 171802 129918
rect 307109 129842 307175 129845
rect 307109 129840 310132 129842
rect 307109 129784 307114 129840
rect 307170 129784 310132 129840
rect 307109 129782 310132 129784
rect 307109 129779 307175 129782
rect 252461 129570 252527 129573
rect 248860 129568 252527 129570
rect 248860 129512 252466 129568
rect 252522 129512 252527 129568
rect 248860 129510 252527 129512
rect 252461 129507 252527 129510
rect 323025 129434 323091 129437
rect 325049 129434 325115 129437
rect 321908 129432 325115 129434
rect 321908 129376 323030 129432
rect 323086 129376 325054 129432
rect 325110 129376 325115 129432
rect 321908 129374 325115 129376
rect 323025 129371 323091 129374
rect 325049 129371 325115 129374
rect 386597 129434 386663 129437
rect 386597 129432 390172 129434
rect 386597 129376 386602 129432
rect 386658 129376 390172 129432
rect 386597 129374 390172 129376
rect 386597 129371 386663 129374
rect 66069 129298 66135 129301
rect 68142 129298 68816 129304
rect 66069 129296 68816 129298
rect 66069 129240 66074 129296
rect 66130 129244 68816 129296
rect 66130 129240 68202 129244
rect 66069 129238 68202 129240
rect 66069 129235 66135 129238
rect 214005 129298 214071 129301
rect 307477 129298 307543 129301
rect 214005 129296 217212 129298
rect 214005 129240 214010 129296
rect 214066 129240 217212 129296
rect 214005 129238 217212 129240
rect 307477 129296 310132 129298
rect 307477 129240 307482 129296
rect 307538 129240 310132 129296
rect 307477 129238 310132 129240
rect 214005 129235 214071 129238
rect 307477 129235 307543 129238
rect 251725 129162 251791 129165
rect 248860 129160 251791 129162
rect 248860 129104 251730 129160
rect 251786 129104 251791 129160
rect 248860 129102 251791 129104
rect 251725 129099 251791 129102
rect 257838 128964 257844 129028
rect 257908 129026 257914 129028
rect 300853 129026 300919 129029
rect 257908 129024 300919 129026
rect 257908 128968 300858 129024
rect 300914 128968 300919 129024
rect 257908 128966 300919 128968
rect 257908 128964 257914 128966
rect 300853 128963 300919 128966
rect 340781 129026 340847 129029
rect 342294 129026 342300 129028
rect 340781 129024 342300 129026
rect 340781 128968 340786 129024
rect 340842 128968 342300 129024
rect 340781 128966 342300 128968
rect 340781 128963 340847 128966
rect 342294 128964 342300 128966
rect 342364 129026 342370 129028
rect 373441 129026 373507 129029
rect 342364 129024 373507 129026
rect 342364 128968 373446 129024
rect 373502 128968 373507 129024
rect 342364 128966 373507 128968
rect 342364 128964 342370 128966
rect 373441 128963 373507 128966
rect 307661 128890 307727 128893
rect 307661 128888 310132 128890
rect 307661 128832 307666 128888
rect 307722 128832 310132 128888
rect 307661 128830 310132 128832
rect 307661 128827 307727 128830
rect 213913 128754 213979 128757
rect 213913 128752 217212 128754
rect 213913 128696 213918 128752
rect 213974 128696 217212 128752
rect 213913 128694 217212 128696
rect 213913 128691 213979 128694
rect 252369 128618 252435 128621
rect 324313 128618 324379 128621
rect 248860 128616 252435 128618
rect 248860 128560 252374 128616
rect 252430 128560 252435 128616
rect 248860 128558 252435 128560
rect 321908 128616 324379 128618
rect 321908 128560 324318 128616
rect 324374 128560 324379 128616
rect 321908 128558 324379 128560
rect 252369 128555 252435 128558
rect 324313 128555 324379 128558
rect 301446 128420 301452 128484
rect 301516 128482 301522 128484
rect 301516 128422 310132 128482
rect 301516 128420 301522 128422
rect 252461 128210 252527 128213
rect 248860 128208 252527 128210
rect 248860 128152 252466 128208
rect 252522 128152 252527 128208
rect 248860 128150 252527 128152
rect 252461 128147 252527 128150
rect 67633 128074 67699 128077
rect 68142 128074 68816 128080
rect 67633 128072 68816 128074
rect 67633 128016 67638 128072
rect 67694 128020 68816 128072
rect 67694 128016 68202 128020
rect 67633 128014 68202 128016
rect 67633 128011 67699 128014
rect 213913 128074 213979 128077
rect 307477 128074 307543 128077
rect 213913 128072 217212 128074
rect 213913 128016 213918 128072
rect 213974 128016 217212 128072
rect 213913 128014 217212 128016
rect 307477 128072 310132 128074
rect 307477 128016 307482 128072
rect 307538 128016 310132 128072
rect 307477 128014 310132 128016
rect 213913 128011 213979 128014
rect 307477 128011 307543 128014
rect 324313 127802 324379 127805
rect 321908 127800 324379 127802
rect 321908 127744 324318 127800
rect 324374 127744 324379 127800
rect 321908 127742 324379 127744
rect 324313 127739 324379 127742
rect 251950 127666 251956 127668
rect 248860 127606 251956 127666
rect 251950 127604 251956 127606
rect 252020 127604 252026 127668
rect 307661 127666 307727 127669
rect 307661 127664 310132 127666
rect 307661 127608 307666 127664
rect 307722 127608 310132 127664
rect 307661 127606 310132 127608
rect 307661 127603 307727 127606
rect 200070 127334 217212 127394
rect 167678 127196 167684 127260
rect 167748 127258 167754 127260
rect 200070 127258 200130 127334
rect 252369 127258 252435 127261
rect 167748 127198 200130 127258
rect 248860 127256 252435 127258
rect 248860 127200 252374 127256
rect 252430 127200 252435 127256
rect 248860 127198 252435 127200
rect 167748 127196 167754 127198
rect 252369 127195 252435 127198
rect 307569 127258 307635 127261
rect 307569 127256 310132 127258
rect 307569 127200 307574 127256
rect 307630 127200 310132 127256
rect 307569 127198 310132 127200
rect 307569 127195 307635 127198
rect 324497 127122 324563 127125
rect 321908 127120 324563 127122
rect 321908 127064 324502 127120
rect 324558 127064 324563 127120
rect 321908 127062 324563 127064
rect 324497 127059 324563 127062
rect 296670 126790 310132 126850
rect 214005 126714 214071 126717
rect 252461 126714 252527 126717
rect 214005 126712 217212 126714
rect 214005 126656 214010 126712
rect 214066 126656 217212 126712
rect 214005 126654 217212 126656
rect 248860 126712 252527 126714
rect 248860 126656 252466 126712
rect 252522 126656 252527 126712
rect 248860 126654 252527 126656
rect 214005 126651 214071 126654
rect 252461 126651 252527 126654
rect 66161 126306 66227 126309
rect 68142 126306 68816 126312
rect 66161 126304 68816 126306
rect 66161 126248 66166 126304
rect 66222 126252 68816 126304
rect 252461 126306 252527 126309
rect 66222 126248 68202 126252
rect 66161 126246 68202 126248
rect 66161 126243 66227 126246
rect 248860 126304 252527 126306
rect 248860 126248 252466 126304
rect 252522 126248 252527 126304
rect 248860 126246 252527 126248
rect 252461 126243 252527 126246
rect 213913 126034 213979 126037
rect 213913 126032 217212 126034
rect 213913 125976 213918 126032
rect 213974 125976 217212 126032
rect 213913 125974 217212 125976
rect 213913 125971 213979 125974
rect 287646 125836 287652 125900
rect 287716 125898 287722 125900
rect 296670 125898 296730 126790
rect 571333 126578 571399 126581
rect 569940 126576 571399 126578
rect 569940 126520 571338 126576
rect 571394 126520 571399 126576
rect 569940 126518 571399 126520
rect 571333 126515 571399 126518
rect 307569 126442 307635 126445
rect 307569 126440 310132 126442
rect 307569 126384 307574 126440
rect 307630 126384 310132 126440
rect 307569 126382 310132 126384
rect 307569 126379 307635 126382
rect 324313 126306 324379 126309
rect 321908 126304 324379 126306
rect 321908 126248 324318 126304
rect 324374 126248 324379 126304
rect 321908 126246 324379 126248
rect 324313 126243 324379 126246
rect 387609 126034 387675 126037
rect 579613 126034 579679 126037
rect 583520 126034 584960 126124
rect 387609 126032 390172 126034
rect 387609 125976 387614 126032
rect 387670 125976 390172 126032
rect 387609 125974 390172 125976
rect 579613 126032 584960 126034
rect 579613 125976 579618 126032
rect 579674 125976 584960 126032
rect 579613 125974 584960 125976
rect 387609 125971 387675 125974
rect 579613 125971 579679 125974
rect 287716 125838 296730 125898
rect 307661 125898 307727 125901
rect 307661 125896 310132 125898
rect 307661 125840 307666 125896
rect 307722 125840 310132 125896
rect 583520 125884 584960 125974
rect 307661 125838 310132 125840
rect 287716 125836 287722 125838
rect 307661 125835 307727 125838
rect 252369 125762 252435 125765
rect 248860 125760 252435 125762
rect 248860 125704 252374 125760
rect 252430 125704 252435 125760
rect 248860 125702 252435 125704
rect 252369 125699 252435 125702
rect 306741 125490 306807 125493
rect 324313 125490 324379 125493
rect 306741 125488 310132 125490
rect 306741 125432 306746 125488
rect 306802 125432 310132 125488
rect 306741 125430 310132 125432
rect 321908 125488 324379 125490
rect 321908 125432 324318 125488
rect 324374 125432 324379 125488
rect 321908 125430 324379 125432
rect 306741 125427 306807 125430
rect 324313 125427 324379 125430
rect 214005 125354 214071 125357
rect 251173 125354 251239 125357
rect 214005 125352 217212 125354
rect 214005 125296 214010 125352
rect 214066 125296 217212 125352
rect 214005 125294 217212 125296
rect 248860 125352 251239 125354
rect 248860 125296 251178 125352
rect 251234 125296 251239 125352
rect 248860 125294 251239 125296
rect 214005 125291 214071 125294
rect 251173 125291 251239 125294
rect 66161 125218 66227 125221
rect 68142 125218 68816 125224
rect 66161 125216 68816 125218
rect 66161 125160 66166 125216
rect 66222 125164 68816 125216
rect 66222 125160 68202 125164
rect 66161 125158 68202 125160
rect 66161 125155 66227 125158
rect 64781 124266 64847 124269
rect 66161 124266 66227 124269
rect 64781 124264 66227 124266
rect 64781 124208 64786 124264
rect 64842 124208 66166 124264
rect 66222 124208 66227 124264
rect 64781 124206 66227 124208
rect 64781 124203 64847 124206
rect 66161 124203 66227 124206
rect -960 123572 480 123812
rect 307477 125082 307543 125085
rect 307477 125080 310132 125082
rect 307477 125024 307482 125080
rect 307538 125024 310132 125080
rect 307477 125022 310132 125024
rect 307477 125019 307543 125022
rect 252461 124810 252527 124813
rect 324405 124810 324471 124813
rect 248860 124808 252527 124810
rect 248860 124752 252466 124808
rect 252522 124752 252527 124808
rect 248860 124750 252527 124752
rect 321908 124808 324471 124810
rect 321908 124752 324410 124808
rect 324466 124752 324471 124808
rect 321908 124750 324471 124752
rect 252461 124747 252527 124750
rect 324405 124747 324471 124750
rect 213913 124674 213979 124677
rect 305637 124674 305703 124677
rect 213913 124672 217212 124674
rect 213913 124616 213918 124672
rect 213974 124616 217212 124672
rect 213913 124614 217212 124616
rect 305637 124672 310132 124674
rect 305637 124616 305642 124672
rect 305698 124616 310132 124672
rect 305637 124614 310132 124616
rect 213913 124611 213979 124614
rect 305637 124611 305703 124614
rect 252369 124402 252435 124405
rect 248860 124400 252435 124402
rect 248860 124344 252374 124400
rect 252430 124344 252435 124400
rect 248860 124342 252435 124344
rect 252369 124339 252435 124342
rect 307661 124266 307727 124269
rect 307661 124264 310132 124266
rect 307661 124208 307666 124264
rect 307722 124208 310132 124264
rect 307661 124206 310132 124208
rect 307661 124203 307727 124206
rect 214005 124130 214071 124133
rect 214005 124128 217212 124130
rect 214005 124072 214010 124128
rect 214066 124072 217212 124128
rect 214005 124070 217212 124072
rect 214005 124067 214071 124070
rect 252461 123994 252527 123997
rect 324313 123994 324379 123997
rect 248860 123992 252527 123994
rect 248860 123936 252466 123992
rect 252522 123936 252527 123992
rect 248860 123934 252527 123936
rect 321908 123992 324379 123994
rect 321908 123936 324318 123992
rect 324374 123936 324379 123992
rect 321908 123934 324379 123936
rect 252461 123931 252527 123934
rect 324313 123931 324379 123934
rect 307477 123858 307543 123861
rect 307477 123856 310132 123858
rect 307477 123800 307482 123856
rect 307538 123800 310132 123856
rect 307477 123798 310132 123800
rect 307477 123795 307543 123798
rect 66069 123586 66135 123589
rect 68142 123586 68816 123592
rect 66069 123584 68816 123586
rect 66069 123528 66074 123584
rect 66130 123532 68816 123584
rect 66130 123528 68202 123532
rect 66069 123526 68202 123528
rect 66069 123523 66135 123526
rect 213913 123450 213979 123453
rect 252369 123450 252435 123453
rect 213913 123448 217212 123450
rect 213913 123392 213918 123448
rect 213974 123392 217212 123448
rect 213913 123390 217212 123392
rect 248860 123448 252435 123450
rect 248860 123392 252374 123448
rect 252430 123392 252435 123448
rect 248860 123390 252435 123392
rect 213913 123387 213979 123390
rect 252369 123387 252435 123390
rect 307661 123450 307727 123453
rect 307661 123448 310132 123450
rect 307661 123392 307666 123448
rect 307722 123392 310132 123448
rect 307661 123390 310132 123392
rect 307661 123387 307727 123390
rect 572621 123314 572687 123317
rect 569940 123312 572687 123314
rect 569940 123256 572626 123312
rect 572682 123256 572687 123312
rect 569940 123254 572687 123256
rect 572621 123251 572687 123254
rect 324405 123178 324471 123181
rect 321908 123176 324471 123178
rect 321908 123120 324410 123176
rect 324466 123120 324471 123176
rect 321908 123118 324471 123120
rect 324405 123115 324471 123118
rect 252277 123042 252343 123045
rect 248860 123040 252343 123042
rect 248860 122984 252282 123040
rect 252338 122984 252343 123040
rect 248860 122982 252343 122984
rect 252277 122979 252343 122982
rect 307109 123042 307175 123045
rect 307109 123040 310132 123042
rect 307109 122984 307114 123040
rect 307170 122984 310132 123040
rect 307109 122982 310132 122984
rect 307109 122979 307175 122982
rect 214005 122770 214071 122773
rect 214005 122768 217212 122770
rect 214005 122712 214010 122768
rect 214066 122712 217212 122768
rect 214005 122710 217212 122712
rect 214005 122707 214071 122710
rect 66161 122634 66227 122637
rect 68142 122634 68816 122640
rect 66161 122632 68816 122634
rect 66161 122576 66166 122632
rect 66222 122580 68816 122632
rect 66222 122576 68202 122580
rect 66161 122574 68202 122576
rect 66161 122571 66227 122574
rect 386781 122634 386847 122637
rect 386781 122632 390172 122634
rect 386781 122576 386786 122632
rect 386842 122576 390172 122632
rect 386781 122574 390172 122576
rect 386781 122571 386847 122574
rect 252461 122498 252527 122501
rect 248860 122496 252527 122498
rect 248860 122440 252466 122496
rect 252522 122440 252527 122496
rect 248860 122438 252527 122440
rect 252461 122435 252527 122438
rect 307477 122498 307543 122501
rect 324313 122498 324379 122501
rect 307477 122496 310132 122498
rect 307477 122440 307482 122496
rect 307538 122440 310132 122496
rect 307477 122438 310132 122440
rect 321908 122496 324379 122498
rect 321908 122440 324318 122496
rect 324374 122440 324379 122496
rect 321908 122438 324379 122440
rect 307477 122435 307543 122438
rect 324313 122435 324379 122438
rect 321645 122226 321711 122229
rect 321645 122224 321754 122226
rect 321645 122168 321650 122224
rect 321706 122168 321754 122224
rect 321645 122163 321754 122168
rect 213913 122090 213979 122093
rect 252369 122090 252435 122093
rect 213913 122088 217212 122090
rect 213913 122032 213918 122088
rect 213974 122032 217212 122088
rect 213913 122030 217212 122032
rect 248860 122088 252435 122090
rect 248860 122032 252374 122088
rect 252430 122032 252435 122088
rect 248860 122030 252435 122032
rect 213913 122027 213979 122030
rect 252369 122027 252435 122030
rect 307569 122090 307635 122093
rect 307569 122088 310132 122090
rect 307569 122032 307574 122088
rect 307630 122032 310132 122088
rect 307569 122030 310132 122032
rect 307569 122027 307635 122030
rect 307661 121682 307727 121685
rect 307661 121680 310132 121682
rect 307661 121624 307666 121680
rect 307722 121624 310132 121680
rect 321694 121652 321754 122163
rect 307661 121622 310132 121624
rect 307661 121619 307727 121622
rect 252461 121546 252527 121549
rect 248860 121544 252527 121546
rect 248860 121488 252466 121544
rect 252522 121488 252527 121544
rect 248860 121486 252527 121488
rect 252461 121483 252527 121486
rect 214005 121410 214071 121413
rect 327533 121412 327599 121413
rect 327533 121410 327580 121412
rect 214005 121408 217212 121410
rect 214005 121352 214010 121408
rect 214066 121352 217212 121408
rect 214005 121350 217212 121352
rect 327452 121408 327580 121410
rect 327644 121410 327650 121412
rect 385534 121410 385540 121412
rect 327452 121352 327538 121408
rect 327452 121350 327580 121352
rect 214005 121347 214071 121350
rect 327533 121348 327580 121350
rect 327644 121350 385540 121410
rect 327644 121348 327650 121350
rect 385534 121348 385540 121350
rect 385604 121348 385610 121412
rect 327533 121347 327599 121348
rect 306741 121274 306807 121277
rect 306741 121272 310132 121274
rect 306741 121216 306746 121272
rect 306802 121216 310132 121272
rect 306741 121214 310132 121216
rect 306741 121211 306807 121214
rect 252461 121138 252527 121141
rect 248860 121136 252527 121138
rect 248860 121080 252466 121136
rect 252522 121080 252527 121136
rect 248860 121078 252527 121080
rect 252461 121075 252527 121078
rect 67449 120866 67515 120869
rect 68142 120866 68816 120872
rect 67449 120864 68816 120866
rect 67449 120808 67454 120864
rect 67510 120812 68816 120864
rect 67510 120808 68202 120812
rect 67449 120806 68202 120808
rect 67449 120803 67515 120806
rect 307569 120866 307635 120869
rect 324313 120866 324379 120869
rect 307569 120864 310132 120866
rect 307569 120808 307574 120864
rect 307630 120808 310132 120864
rect 307569 120806 310132 120808
rect 321908 120864 324379 120866
rect 321908 120808 324318 120864
rect 324374 120808 324379 120864
rect 321908 120806 324379 120808
rect 307569 120803 307635 120806
rect 324313 120803 324379 120806
rect 213913 120730 213979 120733
rect 213913 120728 217212 120730
rect 213913 120672 213918 120728
rect 213974 120672 217212 120728
rect 213913 120670 217212 120672
rect 213913 120667 213979 120670
rect 251541 120594 251607 120597
rect 248860 120592 251607 120594
rect 248860 120536 251546 120592
rect 251602 120536 251607 120592
rect 248860 120534 251607 120536
rect 251541 120531 251607 120534
rect 307661 120458 307727 120461
rect 307661 120456 310132 120458
rect 307661 120400 307666 120456
rect 307722 120400 310132 120456
rect 307661 120398 310132 120400
rect 307661 120395 307727 120398
rect 252369 120186 252435 120189
rect 324405 120186 324471 120189
rect 248860 120184 252435 120186
rect 248860 120128 252374 120184
rect 252430 120128 252435 120184
rect 248860 120126 252435 120128
rect 321908 120184 324471 120186
rect 321908 120128 324410 120184
rect 324466 120128 324471 120184
rect 321908 120126 324471 120128
rect 252369 120123 252435 120126
rect 324405 120123 324471 120126
rect 214097 120050 214163 120053
rect 307661 120050 307727 120053
rect 214097 120048 217212 120050
rect 214097 119992 214102 120048
rect 214158 119992 217212 120048
rect 214097 119990 217212 119992
rect 307661 120048 310132 120050
rect 307661 119992 307666 120048
rect 307722 119992 310132 120048
rect 307661 119990 310132 119992
rect 214097 119987 214163 119990
rect 307661 119987 307727 119990
rect 571425 119778 571491 119781
rect 569940 119776 571491 119778
rect 569940 119720 571430 119776
rect 571486 119720 571491 119776
rect 569940 119718 571491 119720
rect 571425 119715 571491 119718
rect 252461 119642 252527 119645
rect 248860 119640 252527 119642
rect 248860 119584 252466 119640
rect 252522 119584 252527 119640
rect 248860 119582 252527 119584
rect 252461 119579 252527 119582
rect 306557 119642 306623 119645
rect 306557 119640 310132 119642
rect 306557 119584 306562 119640
rect 306618 119584 310132 119640
rect 306557 119582 310132 119584
rect 306557 119579 306623 119582
rect 214005 119506 214071 119509
rect 214005 119504 217212 119506
rect 214005 119448 214010 119504
rect 214066 119448 217212 119504
rect 214005 119446 217212 119448
rect 214005 119443 214071 119446
rect 324313 119370 324379 119373
rect 321908 119368 324379 119370
rect 321908 119312 324318 119368
rect 324374 119312 324379 119368
rect 321908 119310 324379 119312
rect 324313 119307 324379 119310
rect 252093 119234 252159 119237
rect 248860 119232 252159 119234
rect 248860 119176 252098 119232
rect 252154 119176 252159 119232
rect 248860 119174 252159 119176
rect 252093 119171 252159 119174
rect 386873 119234 386939 119237
rect 386873 119232 390172 119234
rect 386873 119176 386878 119232
rect 386934 119176 390172 119232
rect 386873 119174 390172 119176
rect 386873 119171 386939 119174
rect 307109 119098 307175 119101
rect 307109 119096 310132 119098
rect 307109 119040 307114 119096
rect 307170 119040 310132 119096
rect 307109 119038 310132 119040
rect 307109 119035 307175 119038
rect 213913 118826 213979 118829
rect 252369 118826 252435 118829
rect 213913 118824 217212 118826
rect 213913 118768 213918 118824
rect 213974 118768 217212 118824
rect 213913 118766 217212 118768
rect 248860 118824 252435 118826
rect 248860 118768 252374 118824
rect 252430 118768 252435 118824
rect 248860 118766 252435 118768
rect 213913 118763 213979 118766
rect 252369 118763 252435 118766
rect 306925 118690 306991 118693
rect 306925 118688 310132 118690
rect 306925 118632 306930 118688
rect 306986 118632 310132 118688
rect 306925 118630 310132 118632
rect 306925 118627 306991 118630
rect 324313 118554 324379 118557
rect 321908 118552 324379 118554
rect 321908 118496 324318 118552
rect 324374 118496 324379 118552
rect 321908 118494 324379 118496
rect 324313 118491 324379 118494
rect 252461 118282 252527 118285
rect 248860 118280 252527 118282
rect 248860 118224 252466 118280
rect 252522 118224 252527 118280
rect 248860 118222 252527 118224
rect 252461 118219 252527 118222
rect 306557 118282 306623 118285
rect 306557 118280 310132 118282
rect 306557 118224 306562 118280
rect 306618 118224 310132 118280
rect 306557 118222 310132 118224
rect 306557 118219 306623 118222
rect 214005 118146 214071 118149
rect 214005 118144 217212 118146
rect 214005 118088 214010 118144
rect 214066 118088 217212 118144
rect 214005 118086 217212 118088
rect 214005 118083 214071 118086
rect 251817 117874 251883 117877
rect 248860 117872 251883 117874
rect 248860 117816 251822 117872
rect 251878 117816 251883 117872
rect 248860 117814 251883 117816
rect 251817 117811 251883 117814
rect 304206 117812 304212 117876
rect 304276 117874 304282 117876
rect 324405 117874 324471 117877
rect 304276 117814 310132 117874
rect 321908 117872 324471 117874
rect 321908 117816 324410 117872
rect 324466 117816 324471 117872
rect 321908 117814 324471 117816
rect 304276 117812 304282 117814
rect 324405 117811 324471 117814
rect 213913 117466 213979 117469
rect 307661 117466 307727 117469
rect 213913 117464 217212 117466
rect 213913 117408 213918 117464
rect 213974 117408 217212 117464
rect 213913 117406 217212 117408
rect 307661 117464 310132 117466
rect 307661 117408 307666 117464
rect 307722 117408 310132 117464
rect 307661 117406 310132 117408
rect 213913 117403 213979 117406
rect 307661 117403 307727 117406
rect 252369 117330 252435 117333
rect 248860 117328 252435 117330
rect 248860 117272 252374 117328
rect 252430 117272 252435 117328
rect 248860 117270 252435 117272
rect 252369 117267 252435 117270
rect 307569 117058 307635 117061
rect 324313 117058 324379 117061
rect 307569 117056 310132 117058
rect 307569 117000 307574 117056
rect 307630 117000 310132 117056
rect 307569 116998 310132 117000
rect 321908 117056 324379 117058
rect 321908 117000 324318 117056
rect 324374 117000 324379 117056
rect 321908 116998 324379 117000
rect 307569 116995 307635 116998
rect 324313 116995 324379 116998
rect 252461 116922 252527 116925
rect 248860 116920 252527 116922
rect 248860 116864 252466 116920
rect 252522 116864 252527 116920
rect 248860 116862 252527 116864
rect 252461 116859 252527 116862
rect 213177 116786 213243 116789
rect 213177 116784 217212 116786
rect 213177 116728 213182 116784
rect 213238 116728 217212 116784
rect 213177 116726 217212 116728
rect 213177 116723 213243 116726
rect 307477 116650 307543 116653
rect 307477 116648 310132 116650
rect 307477 116592 307482 116648
rect 307538 116592 310132 116648
rect 307477 116590 310132 116592
rect 307477 116587 307543 116590
rect 357341 116514 357407 116517
rect 387190 116514 387196 116516
rect 357341 116512 387196 116514
rect 357341 116456 357346 116512
rect 357402 116456 387196 116512
rect 357341 116454 387196 116456
rect 357341 116451 357407 116454
rect 387190 116452 387196 116454
rect 387260 116452 387266 116516
rect 572621 116514 572687 116517
rect 569940 116512 572687 116514
rect 569940 116456 572626 116512
rect 572682 116456 572687 116512
rect 569940 116454 572687 116456
rect 572621 116451 572687 116454
rect 252001 116378 252067 116381
rect 324497 116378 324563 116381
rect 248860 116376 252067 116378
rect 248860 116320 252006 116376
rect 252062 116320 252067 116376
rect 248860 116318 252067 116320
rect 321908 116376 324563 116378
rect 321908 116320 324502 116376
rect 324558 116320 324563 116376
rect 321908 116318 324563 116320
rect 252001 116315 252067 116318
rect 324497 116315 324563 116318
rect 307661 116242 307727 116245
rect 307661 116240 310132 116242
rect 307661 116184 307666 116240
rect 307722 116184 310132 116240
rect 307661 116182 310132 116184
rect 307661 116179 307727 116182
rect 213913 116106 213979 116109
rect 213913 116104 217212 116106
rect 213913 116048 213918 116104
rect 213974 116048 217212 116104
rect 213913 116046 217212 116048
rect 213913 116043 213979 116046
rect 251909 115970 251975 115973
rect 248860 115968 251975 115970
rect 248860 115912 251914 115968
rect 251970 115912 251975 115968
rect 248860 115910 251975 115912
rect 251909 115907 251975 115910
rect 307017 115698 307083 115701
rect 386873 115698 386939 115701
rect 307017 115696 310132 115698
rect 307017 115640 307022 115696
rect 307078 115640 310132 115696
rect 307017 115638 310132 115640
rect 386873 115696 390172 115698
rect 386873 115640 386878 115696
rect 386934 115640 390172 115696
rect 386873 115638 390172 115640
rect 307017 115635 307083 115638
rect 386873 115635 386939 115638
rect 324313 115562 324379 115565
rect 321908 115560 324379 115562
rect 321908 115504 324318 115560
rect 324374 115504 324379 115560
rect 321908 115502 324379 115504
rect 324313 115499 324379 115502
rect 214005 115426 214071 115429
rect 252277 115426 252343 115429
rect 214005 115424 217212 115426
rect 214005 115368 214010 115424
rect 214066 115368 217212 115424
rect 214005 115366 217212 115368
rect 248860 115424 252343 115426
rect 248860 115368 252282 115424
rect 252338 115368 252343 115424
rect 248860 115366 252343 115368
rect 214005 115363 214071 115366
rect 252277 115363 252343 115366
rect 307477 115290 307543 115293
rect 307477 115288 310132 115290
rect 307477 115232 307482 115288
rect 307538 115232 310132 115288
rect 307477 115230 310132 115232
rect 307477 115227 307543 115230
rect 346301 115154 346367 115157
rect 389766 115154 389772 115156
rect 346301 115152 389772 115154
rect 346301 115096 346306 115152
rect 346362 115096 389772 115152
rect 346301 115094 389772 115096
rect 346301 115091 346367 115094
rect 389766 115092 389772 115094
rect 389836 115092 389842 115156
rect 252001 115018 252067 115021
rect 248860 115016 252067 115018
rect 248860 114960 252006 115016
rect 252062 114960 252067 115016
rect 248860 114958 252067 114960
rect 252001 114955 252067 114958
rect 213913 114882 213979 114885
rect 307109 114882 307175 114885
rect 213913 114880 217212 114882
rect 213913 114824 213918 114880
rect 213974 114824 217212 114880
rect 213913 114822 217212 114824
rect 307109 114880 310132 114882
rect 307109 114824 307114 114880
rect 307170 114824 310132 114880
rect 307109 114822 310132 114824
rect 213913 114819 213979 114822
rect 307109 114819 307175 114822
rect 324405 114746 324471 114749
rect 321908 114744 324471 114746
rect 321908 114688 324410 114744
rect 324466 114688 324471 114744
rect 321908 114686 324471 114688
rect 324405 114683 324471 114686
rect 252461 114474 252527 114477
rect 248860 114472 252527 114474
rect 248860 114416 252466 114472
rect 252522 114416 252527 114472
rect 248860 114414 252527 114416
rect 252461 114411 252527 114414
rect 307569 114474 307635 114477
rect 307569 114472 310132 114474
rect 307569 114416 307574 114472
rect 307630 114416 310132 114472
rect 307569 114414 310132 114416
rect 307569 114411 307635 114414
rect 214005 114202 214071 114205
rect 214005 114200 217212 114202
rect 214005 114144 214010 114200
rect 214066 114144 217212 114200
rect 214005 114142 217212 114144
rect 214005 114139 214071 114142
rect 251541 114066 251607 114069
rect 248860 114064 251607 114066
rect 248860 114008 251546 114064
rect 251602 114008 251607 114064
rect 248860 114006 251607 114008
rect 251541 114003 251607 114006
rect 306557 114066 306623 114069
rect 324313 114066 324379 114069
rect 306557 114064 310132 114066
rect 306557 114008 306562 114064
rect 306618 114008 310132 114064
rect 306557 114006 310132 114008
rect 321908 114064 324379 114066
rect 321908 114008 324318 114064
rect 324374 114008 324379 114064
rect 321908 114006 324379 114008
rect 306557 114003 306623 114006
rect 324313 114003 324379 114006
rect 301630 113596 301636 113660
rect 301700 113658 301706 113660
rect 301700 113598 310132 113658
rect 301700 113596 301706 113598
rect 213913 113522 213979 113525
rect 251817 113522 251883 113525
rect 213913 113520 217212 113522
rect 213913 113464 213918 113520
rect 213974 113464 217212 113520
rect 213913 113462 217212 113464
rect 248860 113520 251883 113522
rect 248860 113464 251822 113520
rect 251878 113464 251883 113520
rect 248860 113462 251883 113464
rect 213913 113459 213979 113462
rect 251817 113459 251883 113462
rect 307661 113250 307727 113253
rect 324405 113250 324471 113253
rect 307661 113248 310132 113250
rect 307661 113192 307666 113248
rect 307722 113192 310132 113248
rect 307661 113190 310132 113192
rect 321908 113248 324471 113250
rect 321908 113192 324410 113248
rect 324466 113192 324471 113248
rect 321908 113190 324471 113192
rect 307661 113187 307727 113190
rect 324405 113187 324471 113190
rect 252369 113114 252435 113117
rect 248860 113112 252435 113114
rect 248860 113056 252374 113112
rect 252430 113056 252435 113112
rect 248860 113054 252435 113056
rect 252369 113051 252435 113054
rect 571517 112978 571583 112981
rect 569940 112976 571583 112978
rect 569940 112920 571522 112976
rect 571578 112920 571583 112976
rect 569940 112918 571583 112920
rect 571517 112915 571583 112918
rect 214005 112842 214071 112845
rect 579889 112842 579955 112845
rect 583520 112842 584960 112932
rect 214005 112840 217212 112842
rect 214005 112784 214010 112840
rect 214066 112784 217212 112840
rect 214005 112782 217212 112784
rect 579889 112840 584960 112842
rect 579889 112784 579894 112840
rect 579950 112784 584960 112840
rect 579889 112782 584960 112784
rect 214005 112779 214071 112782
rect 579889 112779 579955 112782
rect 252461 112706 252527 112709
rect 248860 112704 252527 112706
rect 248860 112648 252466 112704
rect 252522 112648 252527 112704
rect 248860 112646 252527 112648
rect 252461 112643 252527 112646
rect 296670 112646 310132 112706
rect 583520 112692 584960 112782
rect 213913 112162 213979 112165
rect 251541 112162 251607 112165
rect 213913 112160 217212 112162
rect 213913 112104 213918 112160
rect 213974 112104 217212 112160
rect 213913 112102 217212 112104
rect 248860 112160 251607 112162
rect 248860 112104 251546 112160
rect 251602 112104 251607 112160
rect 248860 112102 251607 112104
rect 213913 112099 213979 112102
rect 251541 112099 251607 112102
rect 283414 112100 283420 112164
rect 283484 112162 283490 112164
rect 296670 112162 296730 112646
rect 324313 112434 324379 112437
rect 321908 112432 324379 112434
rect 321908 112376 324318 112432
rect 324374 112376 324379 112432
rect 321908 112374 324379 112376
rect 324313 112371 324379 112374
rect 387558 112372 387564 112436
rect 387628 112434 387634 112436
rect 387628 112374 390172 112434
rect 387628 112372 387634 112374
rect 307569 112298 307635 112301
rect 307569 112296 310132 112298
rect 307569 112240 307574 112296
rect 307630 112240 310132 112296
rect 307569 112238 310132 112240
rect 307569 112235 307635 112238
rect 283484 112102 296730 112162
rect 283484 112100 283490 112102
rect 307661 111890 307727 111893
rect 307661 111888 310132 111890
rect 307661 111832 307666 111888
rect 307722 111832 310132 111888
rect 307661 111830 310132 111832
rect 307661 111827 307727 111830
rect 167913 111754 167979 111757
rect 252369 111754 252435 111757
rect 324405 111754 324471 111757
rect 164694 111752 167979 111754
rect 164694 111696 167918 111752
rect 167974 111696 167979 111752
rect 164694 111694 167979 111696
rect 248860 111752 252435 111754
rect 248860 111696 252374 111752
rect 252430 111696 252435 111752
rect 248860 111694 252435 111696
rect 321908 111752 324471 111754
rect 321908 111696 324410 111752
rect 324466 111696 324471 111752
rect 321908 111694 324471 111696
rect -960 110666 480 110756
rect 2773 110666 2839 110669
rect -960 110664 2839 110666
rect -960 110608 2778 110664
rect 2834 110608 2839 110664
rect -960 110606 2839 110608
rect -960 110516 480 110606
rect 2773 110603 2839 110606
rect 167913 111691 167979 111694
rect 252369 111691 252435 111694
rect 324405 111691 324471 111694
rect 214005 111482 214071 111485
rect 307477 111482 307543 111485
rect 214005 111480 217212 111482
rect 214005 111424 214010 111480
rect 214066 111424 217212 111480
rect 214005 111422 217212 111424
rect 307477 111480 310132 111482
rect 307477 111424 307482 111480
rect 307538 111424 310132 111480
rect 307477 111422 310132 111424
rect 214005 111419 214071 111422
rect 307477 111419 307543 111422
rect 251766 111210 251772 111212
rect 248860 111150 251772 111210
rect 251766 111148 251772 111150
rect 251836 111148 251842 111212
rect 307661 111074 307727 111077
rect 307661 111072 310132 111074
rect 307661 111016 307666 111072
rect 307722 111016 310132 111072
rect 307661 111014 310132 111016
rect 307661 111011 307727 111014
rect 324313 110938 324379 110941
rect 321908 110936 324379 110938
rect 321908 110880 324318 110936
rect 324374 110880 324379 110936
rect 321908 110878 324379 110880
rect 324313 110875 324379 110878
rect 213913 110802 213979 110805
rect 252461 110802 252527 110805
rect 213913 110800 217212 110802
rect 213913 110744 213918 110800
rect 213974 110744 217212 110800
rect 213913 110742 217212 110744
rect 248860 110800 252527 110802
rect 248860 110744 252466 110800
rect 252522 110744 252527 110800
rect 248860 110742 252527 110744
rect 213913 110739 213979 110742
rect 252461 110739 252527 110742
rect 307569 110666 307635 110669
rect 307569 110664 310132 110666
rect 307569 110608 307574 110664
rect 307630 110608 310132 110664
rect 307569 110606 310132 110608
rect 307569 110603 307635 110606
rect 214005 110258 214071 110261
rect 252461 110258 252527 110261
rect 214005 110256 217212 110258
rect 214005 110200 214010 110256
rect 214066 110200 217212 110256
rect 214005 110198 217212 110200
rect 248860 110256 252527 110258
rect 248860 110200 252466 110256
rect 252522 110200 252527 110256
rect 248860 110198 252527 110200
rect 214005 110195 214071 110198
rect 252461 110195 252527 110198
rect 306925 110258 306991 110261
rect 306925 110256 310132 110258
rect 306925 110200 306930 110256
rect 306986 110200 310132 110256
rect 306925 110198 310132 110200
rect 306925 110195 306991 110198
rect 167821 110122 167887 110125
rect 324773 110122 324839 110125
rect 164694 110120 167887 110122
rect 164694 110064 167826 110120
rect 167882 110064 167887 110120
rect 164694 110062 167887 110064
rect 321908 110120 324839 110122
rect 321908 110064 324778 110120
rect 324834 110064 324839 110120
rect 321908 110062 324839 110064
rect 167821 110059 167887 110062
rect 324773 110059 324839 110062
rect 252093 109850 252159 109853
rect 248860 109848 252159 109850
rect 248860 109792 252098 109848
rect 252154 109792 252159 109848
rect 248860 109790 252159 109792
rect 252093 109787 252159 109790
rect 307661 109850 307727 109853
rect 307661 109848 310132 109850
rect 307661 109792 307666 109848
rect 307722 109792 310132 109848
rect 307661 109790 310132 109792
rect 307661 109787 307727 109790
rect 329925 109714 329991 109717
rect 387006 109714 387012 109716
rect 329925 109712 387012 109714
rect 329925 109656 329930 109712
rect 329986 109656 387012 109712
rect 329925 109654 387012 109656
rect 329925 109651 329991 109654
rect 387006 109652 387012 109654
rect 387076 109652 387082 109716
rect 570086 109714 570092 109716
rect 569940 109654 570092 109714
rect 570086 109652 570092 109654
rect 570156 109652 570162 109716
rect 213913 109578 213979 109581
rect 213913 109576 217212 109578
rect 213913 109520 213918 109576
rect 213974 109520 217212 109576
rect 213913 109518 217212 109520
rect 213913 109515 213979 109518
rect 324313 109442 324379 109445
rect 321908 109440 324379 109442
rect 321908 109384 324318 109440
rect 324374 109384 324379 109440
rect 321908 109382 324379 109384
rect 324313 109379 324379 109382
rect 252369 109306 252435 109309
rect 248860 109304 252435 109306
rect 248860 109248 252374 109304
rect 252430 109248 252435 109304
rect 248860 109246 252435 109248
rect 252369 109243 252435 109246
rect 307569 109306 307635 109309
rect 307569 109304 310132 109306
rect 307569 109248 307574 109304
rect 307630 109248 310132 109304
rect 307569 109246 310132 109248
rect 307569 109243 307635 109246
rect 386597 109034 386663 109037
rect 386597 109032 390172 109034
rect 386597 108976 386602 109032
rect 386658 108976 390172 109032
rect 386597 108974 390172 108976
rect 386597 108971 386663 108974
rect 214005 108898 214071 108901
rect 252461 108898 252527 108901
rect 214005 108896 217212 108898
rect 214005 108840 214010 108896
rect 214066 108840 217212 108896
rect 214005 108838 217212 108840
rect 248860 108896 252527 108898
rect 248860 108840 252466 108896
rect 252522 108840 252527 108896
rect 248860 108838 252527 108840
rect 214005 108835 214071 108838
rect 252461 108835 252527 108838
rect 307385 108898 307451 108901
rect 307385 108896 310132 108898
rect 307385 108840 307390 108896
rect 307446 108840 310132 108896
rect 307385 108838 310132 108840
rect 307385 108835 307451 108838
rect 168097 108762 168163 108765
rect 164694 108760 168163 108762
rect 164694 108704 168102 108760
rect 168158 108704 168163 108760
rect 164694 108702 168163 108704
rect 168097 108699 168163 108702
rect 324405 108626 324471 108629
rect 321908 108624 324471 108626
rect 321908 108568 324410 108624
rect 324466 108568 324471 108624
rect 321908 108566 324471 108568
rect 324405 108563 324471 108566
rect 307477 108490 307543 108493
rect 307477 108488 310132 108490
rect 307477 108432 307482 108488
rect 307538 108432 310132 108488
rect 307477 108430 310132 108432
rect 307477 108427 307543 108430
rect 252369 108354 252435 108357
rect 248860 108352 252435 108354
rect 248860 108296 252374 108352
rect 252430 108296 252435 108352
rect 248860 108294 252435 108296
rect 252369 108291 252435 108294
rect 213913 108218 213979 108221
rect 213913 108216 217212 108218
rect 213913 108160 213918 108216
rect 213974 108160 217212 108216
rect 213913 108158 217212 108160
rect 213913 108155 213979 108158
rect 307661 108082 307727 108085
rect 307661 108080 310132 108082
rect 307661 108024 307666 108080
rect 307722 108024 310132 108080
rect 307661 108022 310132 108024
rect 307661 108019 307727 108022
rect 252093 107946 252159 107949
rect 248860 107944 252159 107946
rect 248860 107888 252098 107944
rect 252154 107888 252159 107944
rect 248860 107886 252159 107888
rect 252093 107883 252159 107886
rect 324313 107810 324379 107813
rect 321908 107808 324379 107810
rect 321908 107752 324318 107808
rect 324374 107752 324379 107808
rect 321908 107750 324379 107752
rect 324313 107747 324379 107750
rect 307569 107674 307635 107677
rect 307569 107672 310132 107674
rect 307569 107616 307574 107672
rect 307630 107616 310132 107672
rect 307569 107614 310132 107616
rect 307569 107611 307635 107614
rect 214005 107538 214071 107541
rect 252461 107538 252527 107541
rect 214005 107536 217212 107538
rect 214005 107480 214010 107536
rect 214066 107480 217212 107536
rect 214005 107478 217212 107480
rect 248860 107536 252527 107538
rect 248860 107480 252466 107536
rect 252522 107480 252527 107536
rect 248860 107478 252527 107480
rect 214005 107475 214071 107478
rect 252461 107475 252527 107478
rect 307477 107266 307543 107269
rect 307477 107264 310132 107266
rect 307477 107208 307482 107264
rect 307538 107208 310132 107264
rect 307477 107206 310132 107208
rect 307477 107203 307543 107206
rect 325509 107130 325575 107133
rect 321908 107128 325575 107130
rect 321908 107100 325514 107128
rect 321878 107072 325514 107100
rect 325570 107072 325575 107128
rect 321878 107070 325575 107072
rect 251541 106994 251607 106997
rect 248860 106992 251607 106994
rect 248860 106936 251546 106992
rect 251602 106936 251607 106992
rect 248860 106934 251607 106936
rect 251541 106931 251607 106934
rect 213913 106858 213979 106861
rect 307569 106858 307635 106861
rect 321553 106858 321619 106861
rect 213913 106856 217212 106858
rect 213913 106800 213918 106856
rect 213974 106800 217212 106856
rect 213913 106798 217212 106800
rect 307569 106856 310132 106858
rect 307569 106800 307574 106856
rect 307630 106800 310132 106856
rect 307569 106798 310132 106800
rect 321510 106856 321619 106858
rect 321510 106800 321558 106856
rect 321614 106800 321619 106856
rect 213913 106795 213979 106798
rect 307569 106795 307635 106798
rect 321510 106795 321619 106800
rect 321737 106858 321803 106861
rect 321878 106858 321938 107070
rect 325509 107067 325575 107070
rect 570045 106858 570111 106861
rect 321737 106856 321938 106858
rect 321737 106800 321742 106856
rect 321798 106800 321938 106856
rect 321737 106798 321938 106800
rect 569910 106856 570111 106858
rect 569910 106800 570050 106856
rect 570106 106800 570111 106856
rect 569910 106798 570111 106800
rect 321737 106795 321803 106798
rect 252369 106586 252435 106589
rect 248860 106584 252435 106586
rect 248860 106528 252374 106584
rect 252430 106528 252435 106584
rect 248860 106526 252435 106528
rect 252369 106523 252435 106526
rect 307661 106450 307727 106453
rect 307661 106448 310132 106450
rect 307661 106392 307666 106448
rect 307722 106392 310132 106448
rect 307661 106390 310132 106392
rect 307661 106387 307727 106390
rect 305821 106314 305887 106317
rect 307477 106314 307543 106317
rect 305821 106312 307543 106314
rect 305821 106256 305826 106312
rect 305882 106256 307482 106312
rect 307538 106256 307543 106312
rect 321510 106284 321570 106795
rect 569910 106314 569970 106798
rect 570045 106795 570111 106798
rect 571241 106314 571307 106317
rect 569910 106312 571307 106314
rect 569910 106284 571246 106312
rect 305821 106254 307543 106256
rect 569940 106256 571246 106284
rect 571302 106256 571307 106312
rect 569940 106254 571307 106256
rect 305821 106251 305887 106254
rect 307477 106251 307543 106254
rect 571241 106251 571307 106254
rect 214005 106178 214071 106181
rect 387057 106178 387123 106181
rect 387609 106178 387675 106181
rect 214005 106176 217212 106178
rect 214005 106120 214010 106176
rect 214066 106120 217212 106176
rect 214005 106118 217212 106120
rect 387057 106176 387675 106178
rect 387057 106120 387062 106176
rect 387118 106120 387614 106176
rect 387670 106120 387675 106176
rect 387057 106118 387675 106120
rect 214005 106115 214071 106118
rect 387057 106115 387123 106118
rect 387609 106115 387675 106118
rect 251633 106042 251699 106045
rect 248860 106040 251699 106042
rect 248860 105984 251638 106040
rect 251694 105984 251699 106040
rect 248860 105982 251699 105984
rect 251633 105979 251699 105982
rect 305678 105844 305684 105908
rect 305748 105906 305754 105908
rect 305748 105846 310132 105906
rect 305748 105844 305754 105846
rect 214097 105634 214163 105637
rect 252461 105634 252527 105637
rect 214097 105632 217212 105634
rect 214097 105576 214102 105632
rect 214158 105576 217212 105632
rect 214097 105574 217212 105576
rect 248860 105632 252527 105634
rect 248860 105576 252466 105632
rect 252522 105576 252527 105632
rect 248860 105574 252527 105576
rect 214097 105571 214163 105574
rect 252461 105571 252527 105574
rect 387609 105634 387675 105637
rect 387609 105632 390172 105634
rect 387609 105576 387614 105632
rect 387670 105576 390172 105632
rect 387609 105574 390172 105576
rect 387609 105571 387675 105574
rect 307569 105498 307635 105501
rect 324313 105498 324379 105501
rect 307569 105496 310132 105498
rect 307569 105440 307574 105496
rect 307630 105440 310132 105496
rect 307569 105438 310132 105440
rect 321908 105496 324379 105498
rect 321908 105440 324318 105496
rect 324374 105440 324379 105496
rect 321908 105438 324379 105440
rect 307569 105435 307635 105438
rect 324313 105435 324379 105438
rect 252093 105090 252159 105093
rect 248860 105088 252159 105090
rect 248860 105032 252098 105088
rect 252154 105032 252159 105088
rect 248860 105030 252159 105032
rect 252093 105027 252159 105030
rect 307661 105090 307727 105093
rect 307661 105088 310132 105090
rect 307661 105032 307666 105088
rect 307722 105032 310132 105088
rect 307661 105030 310132 105032
rect 307661 105027 307727 105030
rect 213913 104954 213979 104957
rect 213913 104952 217212 104954
rect 213913 104896 213918 104952
rect 213974 104896 217212 104952
rect 213913 104894 217212 104896
rect 213913 104891 213979 104894
rect 324262 104818 324268 104820
rect 321908 104758 324268 104818
rect 324262 104756 324268 104758
rect 324332 104756 324338 104820
rect 251817 104682 251883 104685
rect 248860 104680 251883 104682
rect 248860 104624 251822 104680
rect 251878 104624 251883 104680
rect 248860 104622 251883 104624
rect 251817 104619 251883 104622
rect 307477 104682 307543 104685
rect 307477 104680 310132 104682
rect 307477 104624 307482 104680
rect 307538 104624 310132 104680
rect 307477 104622 310132 104624
rect 307477 104619 307543 104622
rect 214005 104274 214071 104277
rect 252277 104274 252343 104277
rect 214005 104272 217212 104274
rect 214005 104216 214010 104272
rect 214066 104216 217212 104272
rect 214005 104214 217212 104216
rect 251038 104272 252343 104274
rect 251038 104216 252282 104272
rect 252338 104216 252343 104272
rect 251038 104214 252343 104216
rect 214005 104211 214071 104214
rect 251038 104138 251098 104214
rect 252277 104211 252343 104214
rect 307661 104274 307727 104277
rect 307661 104272 310132 104274
rect 307661 104216 307666 104272
rect 307722 104216 310132 104272
rect 307661 104214 310132 104216
rect 307661 104211 307727 104214
rect 248860 104078 251098 104138
rect 251265 104138 251331 104141
rect 295374 104138 295380 104140
rect 251265 104136 295380 104138
rect 251265 104080 251270 104136
rect 251326 104080 295380 104136
rect 251265 104078 295380 104080
rect 251265 104075 251331 104078
rect 295374 104076 295380 104078
rect 295444 104076 295450 104140
rect 322933 104002 322999 104005
rect 321908 104000 322999 104002
rect 321908 103944 322938 104000
rect 322994 103944 322999 104000
rect 321908 103942 322999 103944
rect 322933 103939 322999 103942
rect 305913 103866 305979 103869
rect 305913 103864 310132 103866
rect 305913 103808 305918 103864
rect 305974 103808 310132 103864
rect 305913 103806 310132 103808
rect 305913 103803 305979 103806
rect 252093 103730 252159 103733
rect 248860 103728 252159 103730
rect 248860 103672 252098 103728
rect 252154 103672 252159 103728
rect 248860 103670 252159 103672
rect 252093 103667 252159 103670
rect 213913 103594 213979 103597
rect 213913 103592 217212 103594
rect 213913 103536 213918 103592
rect 213974 103536 217212 103592
rect 213913 103534 217212 103536
rect 213913 103531 213979 103534
rect 306741 103458 306807 103461
rect 306741 103456 310132 103458
rect 306741 103400 306746 103456
rect 306802 103400 310132 103456
rect 306741 103398 310132 103400
rect 306741 103395 306807 103398
rect 252185 103186 252251 103189
rect 325601 103186 325667 103189
rect 248860 103184 252251 103186
rect 248860 103128 252190 103184
rect 252246 103128 252251 103184
rect 248860 103126 252251 103128
rect 321908 103184 325667 103186
rect 321908 103128 325606 103184
rect 325662 103128 325667 103184
rect 321908 103126 325667 103128
rect 252185 103123 252251 103126
rect 325601 103123 325667 103126
rect 307477 103050 307543 103053
rect 307477 103048 310132 103050
rect 307477 102992 307482 103048
rect 307538 102992 310132 103048
rect 307477 102990 310132 102992
rect 307477 102987 307543 102990
rect 214005 102914 214071 102917
rect 214005 102912 217212 102914
rect 214005 102856 214010 102912
rect 214066 102856 217212 102912
rect 214005 102854 217212 102856
rect 214005 102851 214071 102854
rect 251909 102778 251975 102781
rect 572621 102778 572687 102781
rect 248860 102776 251975 102778
rect 248860 102720 251914 102776
rect 251970 102720 251975 102776
rect 248860 102718 251975 102720
rect 569940 102776 572687 102778
rect 569940 102720 572626 102776
rect 572682 102720 572687 102776
rect 569940 102718 572687 102720
rect 251909 102715 251975 102718
rect 572621 102715 572687 102718
rect 307661 102506 307727 102509
rect 324405 102506 324471 102509
rect 307661 102504 310132 102506
rect 307661 102448 307666 102504
rect 307722 102448 310132 102504
rect 307661 102446 310132 102448
rect 321908 102504 324471 102506
rect 321908 102448 324410 102504
rect 324466 102448 324471 102504
rect 321908 102446 324471 102448
rect 307661 102443 307727 102446
rect 324405 102443 324471 102446
rect 68142 102316 68816 102376
rect 64689 102234 64755 102237
rect 68142 102234 68202 102316
rect 64689 102232 68202 102234
rect 64689 102176 64694 102232
rect 64750 102176 68202 102232
rect 64689 102174 68202 102176
rect 64689 102171 64755 102174
rect 213913 102234 213979 102237
rect 252461 102234 252527 102237
rect 213913 102232 217212 102234
rect 213913 102176 213918 102232
rect 213974 102176 217212 102232
rect 213913 102174 217212 102176
rect 248860 102232 252527 102234
rect 248860 102176 252466 102232
rect 252522 102176 252527 102232
rect 248860 102174 252527 102176
rect 213913 102171 213979 102174
rect 252461 102171 252527 102174
rect 335854 102172 335860 102236
rect 335924 102234 335930 102236
rect 335924 102174 390172 102234
rect 335924 102172 335930 102174
rect 306741 102098 306807 102101
rect 306741 102096 310132 102098
rect 306741 102040 306746 102096
rect 306802 102040 310132 102096
rect 306741 102038 310132 102040
rect 306741 102035 306807 102038
rect 252369 101826 252435 101829
rect 248860 101824 252435 101826
rect 248860 101768 252374 101824
rect 252430 101768 252435 101824
rect 248860 101766 252435 101768
rect 252369 101763 252435 101766
rect 307477 101690 307543 101693
rect 307477 101688 310132 101690
rect 307477 101632 307482 101688
rect 307538 101632 310132 101688
rect 307477 101630 310132 101632
rect 307477 101627 307543 101630
rect 214598 101492 214604 101556
rect 214668 101554 214674 101556
rect 214668 101494 217212 101554
rect 214668 101492 214674 101494
rect 251817 101418 251883 101421
rect 248860 101416 251883 101418
rect 248860 101360 251822 101416
rect 251878 101360 251883 101416
rect 248860 101358 251883 101360
rect 251817 101355 251883 101358
rect 252461 101418 252527 101421
rect 271086 101418 271092 101420
rect 252461 101416 271092 101418
rect 252461 101360 252466 101416
rect 252522 101360 271092 101416
rect 252461 101358 271092 101360
rect 252461 101355 252527 101358
rect 271086 101356 271092 101358
rect 271156 101356 271162 101420
rect 307569 101282 307635 101285
rect 307569 101280 310132 101282
rect 307569 101224 307574 101280
rect 307630 101224 310132 101280
rect 307569 101222 310132 101224
rect 307569 101219 307635 101222
rect 321694 101149 321754 101660
rect 321645 101144 321754 101149
rect 321645 101088 321650 101144
rect 321706 101088 321754 101144
rect 321645 101086 321754 101088
rect 321645 101083 321711 101086
rect 213913 101010 213979 101013
rect 213913 101008 217212 101010
rect 213913 100952 213918 101008
rect 213974 100952 217212 101008
rect 213913 100950 217212 100952
rect 213913 100947 213979 100950
rect 252093 100874 252159 100877
rect 248860 100872 252159 100874
rect 248860 100816 252098 100872
rect 252154 100816 252159 100872
rect 248860 100814 252159 100816
rect 252093 100811 252159 100814
rect 307661 100874 307727 100877
rect 324589 100874 324655 100877
rect 307661 100872 310132 100874
rect 307661 100816 307666 100872
rect 307722 100816 310132 100872
rect 307661 100814 310132 100816
rect 321908 100872 324655 100874
rect 321908 100816 324594 100872
rect 324650 100816 324655 100872
rect 321908 100814 324655 100816
rect 307661 100811 307727 100814
rect 324589 100811 324655 100814
rect 67725 100738 67791 100741
rect 68142 100738 68816 100744
rect 67725 100736 68816 100738
rect 67725 100680 67730 100736
rect 67786 100684 68816 100736
rect 67786 100680 68202 100684
rect 67725 100678 68202 100680
rect 67725 100675 67791 100678
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 252001 100466 252067 100469
rect 248860 100464 252067 100466
rect 248860 100408 252006 100464
rect 252062 100408 252067 100464
rect 248860 100406 252067 100408
rect 252001 100403 252067 100406
rect 307661 100466 307727 100469
rect 307661 100464 310132 100466
rect 307661 100408 307666 100464
rect 307722 100408 310132 100464
rect 307661 100406 310132 100408
rect 307661 100403 307727 100406
rect 214005 100330 214071 100333
rect 214005 100328 217212 100330
rect 214005 100272 214010 100328
rect 214066 100272 217212 100328
rect 214005 100270 217212 100272
rect 214005 100267 214071 100270
rect 322933 100194 322999 100197
rect 321908 100192 322999 100194
rect 321908 100136 322938 100192
rect 322994 100136 322999 100192
rect 321908 100134 322999 100136
rect 322933 100131 322999 100134
rect 307477 100058 307543 100061
rect 307477 100056 310132 100058
rect 307477 100000 307482 100056
rect 307538 100000 310132 100056
rect 307477 99998 310132 100000
rect 307477 99995 307543 99998
rect 251909 99922 251975 99925
rect 248860 99920 251975 99922
rect 248860 99864 251914 99920
rect 251970 99864 251975 99920
rect 248860 99862 251975 99864
rect 251909 99859 251975 99862
rect 214097 99650 214163 99653
rect 214097 99648 217212 99650
rect 214097 99592 214102 99648
rect 214158 99592 217212 99648
rect 214097 99590 217212 99592
rect 214097 99587 214163 99590
rect 302734 99588 302740 99652
rect 302804 99650 302810 99652
rect 302804 99590 310132 99650
rect 302804 99588 302810 99590
rect 252093 99514 252159 99517
rect 248860 99512 252159 99514
rect 248860 99456 252098 99512
rect 252154 99456 252159 99512
rect 248860 99454 252159 99456
rect 252093 99451 252159 99454
rect 305729 99514 305795 99517
rect 307661 99514 307727 99517
rect 305729 99512 307727 99514
rect 305729 99456 305734 99512
rect 305790 99456 307666 99512
rect 307722 99456 307727 99512
rect 305729 99454 307727 99456
rect 569910 99514 569970 100028
rect 570045 99514 570111 99517
rect 569910 99512 570111 99514
rect 569910 99456 570050 99512
rect 570106 99456 570111 99512
rect 569910 99454 570111 99456
rect 305729 99451 305795 99454
rect 307661 99451 307727 99454
rect 570045 99451 570111 99454
rect 580349 99514 580415 99517
rect 583520 99514 584960 99604
rect 580349 99512 584960 99514
rect 580349 99456 580354 99512
rect 580410 99456 584960 99512
rect 580349 99454 584960 99456
rect 580349 99451 580415 99454
rect 324313 99378 324379 99381
rect 321908 99376 324379 99378
rect 321908 99320 324318 99376
rect 324374 99320 324379 99376
rect 583520 99364 584960 99454
rect 321908 99318 324379 99320
rect 324313 99315 324379 99318
rect 306557 99106 306623 99109
rect 306557 99104 310132 99106
rect 306557 99048 306562 99104
rect 306618 99048 310132 99104
rect 306557 99046 310132 99048
rect 306557 99043 306623 99046
rect 213913 98970 213979 98973
rect 251173 98970 251239 98973
rect 213913 98968 217212 98970
rect 213913 98912 213918 98968
rect 213974 98912 217212 98968
rect 213913 98910 217212 98912
rect 248860 98968 251239 98970
rect 248860 98912 251178 98968
rect 251234 98912 251239 98968
rect 248860 98910 251239 98912
rect 213913 98907 213979 98910
rect 251173 98907 251239 98910
rect 386873 98834 386939 98837
rect 386873 98832 390172 98834
rect 386873 98776 386878 98832
rect 386934 98776 390172 98832
rect 386873 98774 390172 98776
rect 386873 98771 386939 98774
rect 307569 98698 307635 98701
rect 307569 98696 310132 98698
rect 307569 98640 307574 98696
rect 307630 98640 310132 98696
rect 307569 98638 310132 98640
rect 307569 98635 307635 98638
rect 252369 98562 252435 98565
rect 324405 98562 324471 98565
rect 248860 98560 252435 98562
rect 248860 98504 252374 98560
rect 252430 98504 252435 98560
rect 248860 98502 252435 98504
rect 321908 98560 324471 98562
rect 321908 98504 324410 98560
rect 324466 98504 324471 98560
rect 321908 98502 324471 98504
rect 252369 98499 252435 98502
rect 324405 98499 324471 98502
rect 214557 98290 214623 98293
rect 307661 98290 307727 98293
rect 214557 98288 217212 98290
rect 214557 98232 214562 98288
rect 214618 98232 217212 98288
rect 214557 98230 217212 98232
rect 307661 98288 310132 98290
rect 307661 98232 307666 98288
rect 307722 98232 310132 98288
rect 307661 98230 310132 98232
rect 214557 98227 214623 98230
rect 307661 98227 307727 98230
rect 252277 98018 252343 98021
rect 248860 98016 252343 98018
rect 248860 97960 252282 98016
rect 252338 97960 252343 98016
rect 248860 97958 252343 97960
rect 252277 97955 252343 97958
rect 251817 97882 251883 97885
rect 273846 97882 273852 97884
rect 251817 97880 273852 97882
rect 251817 97824 251822 97880
rect 251878 97824 273852 97880
rect 251817 97822 273852 97824
rect 251817 97819 251883 97822
rect 273846 97820 273852 97822
rect 273916 97820 273922 97884
rect 307017 97882 307083 97885
rect 324589 97882 324655 97885
rect 307017 97880 310132 97882
rect 307017 97824 307022 97880
rect 307078 97824 310132 97880
rect 307017 97822 310132 97824
rect 321908 97880 324655 97882
rect 321908 97824 324594 97880
rect 324650 97824 324655 97880
rect 321908 97822 324655 97824
rect 307017 97819 307083 97822
rect 324589 97819 324655 97822
rect 213913 97610 213979 97613
rect 251909 97610 251975 97613
rect 213913 97608 217212 97610
rect 213913 97552 213918 97608
rect 213974 97552 217212 97608
rect 213913 97550 217212 97552
rect 248860 97608 251975 97610
rect 248860 97552 251914 97608
rect 251970 97552 251975 97608
rect 248860 97550 251975 97552
rect 213913 97547 213979 97550
rect 251909 97547 251975 97550
rect 307477 97474 307543 97477
rect 307477 97472 310132 97474
rect 307477 97416 307482 97472
rect 307538 97416 310132 97472
rect 307477 97414 310132 97416
rect 307477 97411 307543 97414
rect 167310 97140 167316 97204
rect 167380 97202 167386 97204
rect 214925 97202 214991 97205
rect 167380 97200 214991 97202
rect 167380 97144 214930 97200
rect 214986 97144 214991 97200
rect 167380 97142 214991 97144
rect 167380 97140 167386 97142
rect 214925 97139 214991 97142
rect 569309 97202 569375 97205
rect 579654 97202 579660 97204
rect 569309 97200 579660 97202
rect 569309 97144 569314 97200
rect 569370 97144 579660 97200
rect 569309 97142 579660 97144
rect 569309 97139 569375 97142
rect 579654 97140 579660 97142
rect 579724 97140 579730 97204
rect 249241 97066 249307 97069
rect 251817 97066 251883 97069
rect 248860 97064 251883 97066
rect 248860 97008 249246 97064
rect 249302 97008 251822 97064
rect 251878 97008 251883 97064
rect 248860 97006 251883 97008
rect 249241 97003 249307 97006
rect 251817 97003 251883 97006
rect 307150 97004 307156 97068
rect 307220 97066 307226 97068
rect 307220 97006 310132 97066
rect 307220 97004 307226 97006
rect 214833 96930 214899 96933
rect 214833 96928 217212 96930
rect 214833 96872 214838 96928
rect 214894 96872 217212 96928
rect 214833 96870 217212 96872
rect 214833 96867 214899 96870
rect 321510 96661 321570 97036
rect 251173 96658 251239 96661
rect 252461 96658 252527 96661
rect 248860 96656 252527 96658
rect 248860 96600 251178 96656
rect 251234 96600 252466 96656
rect 252522 96600 252527 96656
rect 248860 96598 252527 96600
rect 251173 96595 251239 96598
rect 252461 96595 252527 96598
rect 307661 96658 307727 96661
rect 321510 96658 321619 96661
rect 324446 96658 324452 96660
rect 307661 96656 310132 96658
rect 307661 96600 307666 96656
rect 307722 96600 310132 96656
rect 307661 96598 310132 96600
rect 321510 96656 324452 96658
rect 321510 96600 321558 96656
rect 321614 96600 324452 96656
rect 321510 96598 324452 96600
rect 307661 96595 307727 96598
rect 321553 96595 321619 96598
rect 324446 96596 324452 96598
rect 324516 96596 324522 96660
rect 571609 96658 571675 96661
rect 569940 96656 571675 96658
rect 569940 96600 571614 96656
rect 571670 96600 571675 96656
rect 569940 96598 571675 96600
rect 571609 96595 571675 96598
rect 322054 96460 322060 96524
rect 322124 96522 322130 96524
rect 574093 96522 574159 96525
rect 322124 96520 574159 96522
rect 322124 96464 574098 96520
rect 574154 96464 574159 96520
rect 322124 96462 574159 96464
rect 322124 96460 322130 96462
rect 574093 96459 574159 96462
rect 213913 96386 213979 96389
rect 324313 96386 324379 96389
rect 213913 96384 217212 96386
rect 213913 96328 213918 96384
rect 213974 96328 217212 96384
rect 213913 96326 217212 96328
rect 321908 96384 324379 96386
rect 321908 96328 324318 96384
rect 324374 96328 324379 96384
rect 321908 96326 324379 96328
rect 213913 96323 213979 96326
rect 324313 96323 324379 96326
rect 324446 96324 324452 96388
rect 324516 96386 324522 96388
rect 362217 96386 362283 96389
rect 324516 96384 362283 96386
rect 324516 96328 362222 96384
rect 362278 96328 362283 96384
rect 324516 96326 362283 96328
rect 324516 96324 324522 96326
rect 362217 96323 362283 96326
rect 387190 96324 387196 96388
rect 387260 96386 387266 96388
rect 571558 96386 571564 96388
rect 387260 96326 571564 96386
rect 387260 96324 387266 96326
rect 571558 96324 571564 96326
rect 571628 96324 571634 96388
rect 307661 96250 307727 96253
rect 307661 96248 310132 96250
rect 218053 95978 218119 95981
rect 219198 95978 219204 95980
rect 218053 95976 219204 95978
rect 218053 95920 218058 95976
rect 218114 95920 219204 95976
rect 218053 95918 219204 95920
rect 218053 95915 218119 95918
rect 219198 95916 219204 95918
rect 219268 95916 219274 95980
rect 248830 95706 248890 96220
rect 307661 96192 307666 96248
rect 307722 96192 310132 96248
rect 307661 96190 310132 96192
rect 307661 96187 307727 96190
rect 389766 96188 389772 96252
rect 389836 96250 389842 96252
rect 571333 96250 571399 96253
rect 389836 96248 571399 96250
rect 389836 96192 571338 96248
rect 571394 96192 571399 96248
rect 389836 96190 571399 96192
rect 389836 96188 389842 96190
rect 571333 96187 571399 96190
rect 250989 95706 251055 95709
rect 248830 95704 251055 95706
rect 248830 95648 250994 95704
rect 251050 95648 251055 95704
rect 248830 95646 251055 95648
rect 250989 95643 251055 95646
rect 173157 95162 173223 95165
rect 321553 95162 321619 95165
rect 173157 95160 321619 95162
rect 173157 95104 173162 95160
rect 173218 95104 321558 95160
rect 321614 95104 321619 95160
rect 173157 95102 321619 95104
rect 173157 95099 173223 95102
rect 321553 95099 321619 95102
rect 376109 95162 376175 95165
rect 582649 95162 582715 95165
rect 376109 95160 582715 95162
rect 376109 95104 376114 95160
rect 376170 95104 582654 95160
rect 582710 95104 582715 95160
rect 376109 95102 582715 95104
rect 376109 95099 376175 95102
rect 582649 95099 582715 95102
rect 380157 95026 380223 95029
rect 575473 95026 575539 95029
rect 380157 95024 575539 95026
rect 380157 94968 380162 95024
rect 380218 94968 575478 95024
rect 575534 94968 575539 95024
rect 380157 94966 575539 94968
rect 380157 94963 380223 94966
rect 575473 94963 575539 94966
rect 60641 94890 60707 94893
rect 191189 94890 191255 94893
rect 60641 94888 191255 94890
rect 60641 94832 60646 94888
rect 60702 94832 191194 94888
rect 191250 94832 191255 94888
rect 60641 94830 191255 94832
rect 60641 94827 60707 94830
rect 191189 94827 191255 94830
rect 112345 94756 112411 94757
rect 113173 94756 113239 94757
rect 123201 94756 123267 94757
rect 151905 94756 151971 94757
rect 112320 94692 112326 94756
rect 112390 94754 112411 94756
rect 112390 94752 112482 94754
rect 112406 94696 112482 94752
rect 112390 94694 112482 94696
rect 112390 94692 112411 94694
rect 113136 94692 113142 94756
rect 113206 94754 113239 94756
rect 113206 94752 113298 94754
rect 113234 94696 113298 94752
rect 113206 94694 113298 94696
rect 113206 94692 113239 94694
rect 119392 94692 119398 94756
rect 119462 94754 119468 94756
rect 119838 94754 119844 94756
rect 119462 94694 119844 94754
rect 119462 94692 119468 94694
rect 119838 94692 119844 94694
rect 119908 94692 119914 94756
rect 123200 94754 123206 94756
rect 123114 94694 123206 94754
rect 123200 94692 123206 94694
rect 123270 94692 123276 94756
rect 151302 94692 151308 94756
rect 151372 94754 151378 94756
rect 151624 94754 151630 94756
rect 151372 94694 151630 94754
rect 151372 94692 151378 94694
rect 151624 94692 151630 94694
rect 151694 94692 151700 94756
rect 151896 94692 151902 94756
rect 151966 94754 151972 94756
rect 151966 94694 152058 94754
rect 151966 94692 151972 94694
rect 112345 94691 112411 94692
rect 113173 94691 113239 94692
rect 123201 94691 123267 94692
rect 151905 94691 151971 94692
rect 125593 94482 125659 94485
rect 167494 94482 167500 94484
rect 125593 94480 167500 94482
rect 125593 94424 125598 94480
rect 125654 94424 167500 94480
rect 125593 94422 167500 94424
rect 125593 94419 125659 94422
rect 167494 94420 167500 94422
rect 167564 94420 167570 94484
rect 116710 93740 116716 93804
rect 116780 93802 116786 93804
rect 116780 93742 122850 93802
rect 116780 93740 116786 93742
rect 121729 93668 121795 93669
rect 121678 93666 121684 93668
rect 121638 93606 121684 93666
rect 121748 93664 121795 93668
rect 121790 93608 121795 93664
rect 121678 93604 121684 93606
rect 121748 93604 121795 93608
rect 122790 93666 122850 93742
rect 169150 93740 169156 93804
rect 169220 93802 169226 93804
rect 324497 93802 324563 93805
rect 169220 93800 324563 93802
rect 169220 93744 324502 93800
rect 324558 93744 324563 93800
rect 169220 93742 324563 93744
rect 169220 93740 169226 93742
rect 324497 93739 324563 93742
rect 389633 93802 389699 93805
rect 571517 93802 571583 93805
rect 389633 93800 571583 93802
rect 389633 93744 389638 93800
rect 389694 93744 571522 93800
rect 571578 93744 571583 93800
rect 389633 93742 571583 93744
rect 389633 93739 389699 93742
rect 571517 93739 571583 93742
rect 171910 93666 171916 93668
rect 122790 93606 171916 93666
rect 171910 93604 171916 93606
rect 171980 93604 171986 93668
rect 538765 93666 538831 93669
rect 574686 93666 574692 93668
rect 538765 93664 574692 93666
rect 538765 93608 538770 93664
rect 538826 93608 574692 93664
rect 538765 93606 574692 93608
rect 121729 93603 121795 93604
rect 538765 93603 538831 93606
rect 574686 93604 574692 93606
rect 574756 93604 574762 93668
rect 93945 93532 94011 93533
rect 107745 93532 107811 93533
rect 151537 93532 151603 93533
rect 93894 93530 93900 93532
rect 93854 93470 93900 93530
rect 93964 93528 94011 93532
rect 107694 93530 107700 93532
rect 94006 93472 94011 93528
rect 93894 93468 93900 93470
rect 93964 93468 94011 93472
rect 107654 93470 107700 93530
rect 107764 93528 107811 93532
rect 151486 93530 151492 93532
rect 107806 93472 107811 93528
rect 107694 93468 107700 93470
rect 107764 93468 107811 93472
rect 151446 93470 151492 93530
rect 151556 93528 151603 93532
rect 151598 93472 151603 93528
rect 151486 93468 151492 93470
rect 151556 93468 151603 93472
rect 93945 93467 94011 93468
rect 107745 93467 107811 93468
rect 151537 93467 151603 93468
rect 110137 93260 110203 93261
rect 128169 93260 128235 93261
rect 324313 93260 324379 93261
rect 110086 93258 110092 93260
rect 110046 93198 110092 93258
rect 110156 93256 110203 93260
rect 128118 93258 128124 93260
rect 110198 93200 110203 93256
rect 110086 93196 110092 93198
rect 110156 93196 110203 93200
rect 128078 93198 128124 93258
rect 128188 93256 128235 93260
rect 324262 93258 324268 93260
rect 128230 93200 128235 93256
rect 128118 93196 128124 93198
rect 128188 93196 128235 93200
rect 324222 93198 324268 93258
rect 324332 93256 324379 93260
rect 324374 93200 324379 93256
rect 324262 93196 324268 93198
rect 324332 93196 324379 93200
rect 110137 93195 110203 93196
rect 128169 93195 128235 93196
rect 324313 93195 324379 93196
rect 128353 93122 128419 93125
rect 214414 93122 214420 93124
rect 128353 93120 214420 93122
rect 128353 93064 128358 93120
rect 128414 93064 214420 93120
rect 128353 93062 214420 93064
rect 128353 93059 128419 93062
rect 214414 93060 214420 93062
rect 214484 93060 214490 93124
rect 85614 92380 85620 92444
rect 85684 92442 85690 92444
rect 85757 92442 85823 92445
rect 85684 92440 85823 92442
rect 85684 92384 85762 92440
rect 85818 92384 85823 92440
rect 85684 92382 85823 92384
rect 85684 92380 85690 92382
rect 85757 92379 85823 92382
rect 87086 92380 87092 92444
rect 87156 92442 87162 92444
rect 87229 92442 87295 92445
rect 88977 92444 89043 92445
rect 88926 92442 88932 92444
rect 87156 92440 87295 92442
rect 87156 92384 87234 92440
rect 87290 92384 87295 92440
rect 87156 92382 87295 92384
rect 88886 92382 88932 92442
rect 88996 92440 89043 92444
rect 89038 92384 89043 92440
rect 87156 92380 87162 92382
rect 87229 92379 87295 92382
rect 88926 92380 88932 92382
rect 88996 92380 89043 92384
rect 99598 92380 99604 92444
rect 99668 92442 99674 92444
rect 100477 92442 100543 92445
rect 99668 92440 100543 92442
rect 99668 92384 100482 92440
rect 100538 92384 100543 92440
rect 99668 92382 100543 92384
rect 99668 92380 99674 92382
rect 88977 92379 89043 92380
rect 100477 92379 100543 92382
rect 106774 92380 106780 92444
rect 106844 92442 106850 92444
rect 107469 92442 107535 92445
rect 106844 92440 107535 92442
rect 106844 92384 107474 92440
rect 107530 92384 107535 92440
rect 106844 92382 107535 92384
rect 106844 92380 106850 92382
rect 107469 92379 107535 92382
rect 109166 92380 109172 92444
rect 109236 92442 109242 92444
rect 109677 92442 109743 92445
rect 109236 92440 109743 92442
rect 109236 92384 109682 92440
rect 109738 92384 109743 92440
rect 109236 92382 109743 92384
rect 109236 92380 109242 92382
rect 109677 92379 109743 92382
rect 111190 92380 111196 92444
rect 111260 92442 111266 92444
rect 111609 92442 111675 92445
rect 114185 92444 114251 92445
rect 118049 92444 118115 92445
rect 124489 92444 124555 92445
rect 125409 92444 125475 92445
rect 125777 92444 125843 92445
rect 129457 92444 129523 92445
rect 135713 92444 135779 92445
rect 114134 92442 114140 92444
rect 111260 92440 111675 92442
rect 111260 92384 111614 92440
rect 111670 92384 111675 92440
rect 111260 92382 111675 92384
rect 114094 92382 114140 92442
rect 114204 92440 114251 92444
rect 117998 92442 118004 92444
rect 114246 92384 114251 92440
rect 111260 92380 111266 92382
rect 111609 92379 111675 92382
rect 114134 92380 114140 92382
rect 114204 92380 114251 92384
rect 117958 92382 118004 92442
rect 118068 92440 118115 92444
rect 124438 92442 124444 92444
rect 118110 92384 118115 92440
rect 117998 92380 118004 92382
rect 118068 92380 118115 92384
rect 124398 92382 124444 92442
rect 124508 92440 124555 92444
rect 125358 92442 125364 92444
rect 124550 92384 124555 92440
rect 124438 92380 124444 92382
rect 124508 92380 124555 92384
rect 125318 92382 125364 92442
rect 125428 92440 125475 92444
rect 125726 92442 125732 92444
rect 125470 92384 125475 92440
rect 125358 92380 125364 92382
rect 125428 92380 125475 92384
rect 125686 92382 125732 92442
rect 125796 92440 125843 92444
rect 129406 92442 129412 92444
rect 125838 92384 125843 92440
rect 125726 92380 125732 92382
rect 125796 92380 125843 92384
rect 129366 92382 129412 92442
rect 129476 92440 129523 92444
rect 135662 92442 135668 92444
rect 129518 92384 129523 92440
rect 129406 92380 129412 92382
rect 129476 92380 129523 92384
rect 135622 92382 135668 92442
rect 135732 92440 135779 92444
rect 135774 92384 135779 92440
rect 135662 92380 135668 92382
rect 135732 92380 135779 92384
rect 114185 92379 114251 92380
rect 118049 92379 118115 92380
rect 124489 92379 124555 92380
rect 125409 92379 125475 92380
rect 125777 92379 125843 92380
rect 129457 92379 129523 92380
rect 135713 92379 135779 92380
rect 374637 92442 374703 92445
rect 405457 92442 405523 92445
rect 374637 92440 405523 92442
rect 374637 92384 374642 92440
rect 374698 92384 405462 92440
rect 405518 92384 405523 92440
rect 374637 92382 405523 92384
rect 374637 92379 374703 92382
rect 405457 92379 405523 92382
rect 115422 92244 115428 92308
rect 115492 92306 115498 92308
rect 167310 92306 167316 92308
rect 115492 92246 167316 92306
rect 115492 92244 115498 92246
rect 167310 92244 167316 92246
rect 167380 92244 167386 92308
rect 151721 92172 151787 92173
rect 151670 92170 151676 92172
rect 151630 92110 151676 92170
rect 151740 92168 151787 92172
rect 151782 92112 151787 92168
rect 151670 92108 151676 92110
rect 151740 92108 151787 92112
rect 151721 92107 151787 92108
rect 115054 91700 115060 91764
rect 115124 91762 115130 91764
rect 115381 91762 115447 91765
rect 115124 91760 115447 91762
rect 115124 91704 115386 91760
rect 115442 91704 115447 91760
rect 115124 91702 115447 91704
rect 115124 91700 115130 91702
rect 115381 91699 115447 91702
rect 104249 91628 104315 91629
rect 104198 91626 104204 91628
rect 104158 91566 104204 91626
rect 104268 91624 104315 91628
rect 104310 91568 104315 91624
rect 104198 91564 104204 91566
rect 104268 91564 104315 91568
rect 131982 91564 131988 91628
rect 132052 91626 132058 91628
rect 132217 91626 132283 91629
rect 151353 91628 151419 91629
rect 151302 91626 151308 91628
rect 132052 91624 132283 91626
rect 132052 91568 132222 91624
rect 132278 91568 132283 91624
rect 132052 91566 132283 91568
rect 151262 91566 151308 91626
rect 151372 91624 151419 91628
rect 151414 91568 151419 91624
rect 132052 91564 132058 91566
rect 104249 91563 104315 91564
rect 132217 91563 132283 91566
rect 151302 91564 151308 91566
rect 151372 91564 151419 91568
rect 151353 91563 151419 91564
rect 98494 91428 98500 91492
rect 98564 91490 98570 91492
rect 99281 91490 99347 91493
rect 101857 91492 101923 91493
rect 101806 91490 101812 91492
rect 98564 91488 99347 91490
rect 98564 91432 99286 91488
rect 99342 91432 99347 91488
rect 98564 91430 99347 91432
rect 101766 91430 101812 91490
rect 101876 91488 101923 91492
rect 101918 91432 101923 91488
rect 98564 91428 98570 91430
rect 99281 91427 99347 91430
rect 101806 91428 101812 91430
rect 101876 91428 101923 91432
rect 122782 91428 122788 91492
rect 122852 91490 122858 91492
rect 124121 91490 124187 91493
rect 122852 91488 124187 91490
rect 122852 91432 124126 91488
rect 124182 91432 124187 91488
rect 122852 91430 124187 91432
rect 122852 91428 122858 91430
rect 101857 91427 101923 91428
rect 124121 91427 124187 91430
rect 98126 91292 98132 91356
rect 98196 91354 98202 91356
rect 99097 91354 99163 91357
rect 98196 91352 99163 91354
rect 98196 91296 99102 91352
rect 99158 91296 99163 91352
rect 98196 91294 99163 91296
rect 98196 91292 98202 91294
rect 99097 91291 99163 91294
rect 101622 91292 101628 91356
rect 101692 91354 101698 91356
rect 102041 91354 102107 91357
rect 101692 91352 102107 91354
rect 101692 91296 102046 91352
rect 102102 91296 102107 91352
rect 101692 91294 102107 91296
rect 101692 91292 101698 91294
rect 102041 91291 102107 91294
rect 102910 91292 102916 91356
rect 102980 91354 102986 91356
rect 103329 91354 103395 91357
rect 102980 91352 103395 91354
rect 102980 91296 103334 91352
rect 103390 91296 103395 91352
rect 102980 91294 103395 91296
rect 102980 91292 102986 91294
rect 103329 91291 103395 91294
rect 105118 91292 105124 91356
rect 105188 91354 105194 91356
rect 106181 91354 106247 91357
rect 119889 91356 119955 91357
rect 119838 91354 119844 91356
rect 105188 91352 106247 91354
rect 105188 91296 106186 91352
rect 106242 91296 106247 91352
rect 105188 91294 106247 91296
rect 119798 91294 119844 91354
rect 119908 91352 119955 91356
rect 119950 91296 119955 91352
rect 105188 91292 105194 91294
rect 106181 91291 106247 91294
rect 119838 91292 119844 91294
rect 119908 91292 119955 91296
rect 120574 91292 120580 91356
rect 120644 91354 120650 91356
rect 120717 91354 120783 91357
rect 120644 91352 120783 91354
rect 120644 91296 120722 91352
rect 120778 91296 120783 91352
rect 120644 91294 120783 91296
rect 120644 91292 120650 91294
rect 119889 91291 119955 91292
rect 120717 91291 120783 91294
rect 126646 91292 126652 91356
rect 126716 91354 126722 91356
rect 126881 91354 126947 91357
rect 126716 91352 126947 91354
rect 126716 91296 126886 91352
rect 126942 91296 126947 91352
rect 126716 91294 126947 91296
rect 126716 91292 126722 91294
rect 126881 91291 126947 91294
rect 74758 91156 74764 91220
rect 74828 91218 74834 91220
rect 75821 91218 75887 91221
rect 74828 91216 75887 91218
rect 74828 91160 75826 91216
rect 75882 91160 75887 91216
rect 74828 91158 75887 91160
rect 74828 91156 74834 91158
rect 75821 91155 75887 91158
rect 84326 91156 84332 91220
rect 84396 91218 84402 91220
rect 85481 91218 85547 91221
rect 84396 91216 85547 91218
rect 84396 91160 85486 91216
rect 85542 91160 85547 91216
rect 84396 91158 85547 91160
rect 84396 91156 84402 91158
rect 85481 91155 85547 91158
rect 86718 91156 86724 91220
rect 86788 91218 86794 91220
rect 86861 91218 86927 91221
rect 86788 91216 86927 91218
rect 86788 91160 86866 91216
rect 86922 91160 86927 91216
rect 86788 91158 86927 91160
rect 86788 91156 86794 91158
rect 86861 91155 86927 91158
rect 90214 91156 90220 91220
rect 90284 91218 90290 91220
rect 90725 91218 90791 91221
rect 90284 91216 90791 91218
rect 90284 91160 90730 91216
rect 90786 91160 90791 91216
rect 90284 91158 90791 91160
rect 90284 91156 90290 91158
rect 90725 91155 90791 91158
rect 91318 91156 91324 91220
rect 91388 91218 91394 91220
rect 92381 91218 92447 91221
rect 91388 91216 92447 91218
rect 91388 91160 92386 91216
rect 92442 91160 92447 91216
rect 91388 91158 92447 91160
rect 91388 91156 91394 91158
rect 92381 91155 92447 91158
rect 92606 91156 92612 91220
rect 92676 91218 92682 91220
rect 93761 91218 93827 91221
rect 92676 91216 93827 91218
rect 92676 91160 93766 91216
rect 93822 91160 93827 91216
rect 92676 91158 93827 91160
rect 92676 91156 92682 91158
rect 93761 91155 93827 91158
rect 94998 91156 95004 91220
rect 95068 91218 95074 91220
rect 95141 91218 95207 91221
rect 95068 91216 95207 91218
rect 95068 91160 95146 91216
rect 95202 91160 95207 91216
rect 95068 91158 95207 91160
rect 95068 91156 95074 91158
rect 95141 91155 95207 91158
rect 96102 91156 96108 91220
rect 96172 91218 96178 91220
rect 96521 91218 96587 91221
rect 97073 91220 97139 91221
rect 97022 91218 97028 91220
rect 96172 91216 96587 91218
rect 96172 91160 96526 91216
rect 96582 91160 96587 91216
rect 96172 91158 96587 91160
rect 96982 91158 97028 91218
rect 97092 91216 97139 91220
rect 97134 91160 97139 91216
rect 96172 91156 96178 91158
rect 96521 91155 96587 91158
rect 97022 91156 97028 91158
rect 97092 91156 97139 91160
rect 97206 91156 97212 91220
rect 97276 91218 97282 91220
rect 97901 91218 97967 91221
rect 99189 91220 99255 91221
rect 100569 91220 100635 91221
rect 99189 91218 99236 91220
rect 97276 91216 97967 91218
rect 97276 91160 97906 91216
rect 97962 91160 97967 91216
rect 97276 91158 97967 91160
rect 99144 91216 99236 91218
rect 99144 91160 99194 91216
rect 99144 91158 99236 91160
rect 97276 91156 97282 91158
rect 97073 91155 97139 91156
rect 97901 91155 97967 91158
rect 99189 91156 99236 91158
rect 99300 91156 99306 91220
rect 100518 91218 100524 91220
rect 100478 91158 100524 91218
rect 100588 91216 100635 91220
rect 101949 91220 102015 91221
rect 101949 91218 101996 91220
rect 100630 91160 100635 91216
rect 100518 91156 100524 91158
rect 100588 91156 100635 91160
rect 101904 91216 101996 91218
rect 101904 91160 101954 91216
rect 101904 91158 101996 91160
rect 99189 91155 99255 91156
rect 100569 91155 100635 91156
rect 101949 91156 101996 91158
rect 102060 91156 102066 91220
rect 103278 91156 103284 91220
rect 103348 91218 103354 91220
rect 103421 91218 103487 91221
rect 103348 91216 103487 91218
rect 103348 91160 103426 91216
rect 103482 91160 103487 91216
rect 103348 91158 103487 91160
rect 103348 91156 103354 91158
rect 101949 91155 102015 91156
rect 103421 91155 103487 91158
rect 104566 91156 104572 91220
rect 104636 91218 104642 91220
rect 104801 91218 104867 91221
rect 106089 91220 106155 91221
rect 106038 91218 106044 91220
rect 104636 91216 104867 91218
rect 104636 91160 104806 91216
rect 104862 91160 104867 91216
rect 104636 91158 104867 91160
rect 105998 91158 106044 91218
rect 106108 91216 106155 91220
rect 106150 91160 106155 91216
rect 104636 91156 104642 91158
rect 104801 91155 104867 91158
rect 106038 91156 106044 91158
rect 106108 91156 106155 91160
rect 106406 91156 106412 91220
rect 106476 91218 106482 91220
rect 107561 91218 107627 91221
rect 106476 91216 107627 91218
rect 106476 91160 107566 91216
rect 107622 91160 107627 91216
rect 106476 91158 107627 91160
rect 106476 91156 106482 91158
rect 106089 91155 106155 91156
rect 107561 91155 107627 91158
rect 108062 91156 108068 91220
rect 108132 91218 108138 91220
rect 108481 91218 108547 91221
rect 108132 91216 108547 91218
rect 108132 91160 108486 91216
rect 108542 91160 108547 91216
rect 108132 91158 108547 91160
rect 108132 91156 108138 91158
rect 108481 91155 108547 91158
rect 109534 91156 109540 91220
rect 109604 91218 109610 91220
rect 110229 91218 110295 91221
rect 109604 91216 110295 91218
rect 109604 91160 110234 91216
rect 110290 91160 110295 91216
rect 109604 91158 110295 91160
rect 109604 91156 109610 91158
rect 110229 91155 110295 91158
rect 110638 91156 110644 91220
rect 110708 91218 110714 91220
rect 111701 91218 111767 91221
rect 110708 91216 111767 91218
rect 110708 91160 111706 91216
rect 111762 91160 111767 91216
rect 110708 91158 111767 91160
rect 110708 91156 110714 91158
rect 111701 91155 111767 91158
rect 111926 91156 111932 91220
rect 111996 91218 112002 91220
rect 113081 91218 113147 91221
rect 111996 91216 113147 91218
rect 111996 91160 113086 91216
rect 113142 91160 113147 91216
rect 111996 91158 113147 91160
rect 111996 91156 112002 91158
rect 113081 91155 113147 91158
rect 113766 91156 113772 91220
rect 113836 91218 113842 91220
rect 113909 91218 113975 91221
rect 115841 91220 115907 91221
rect 117129 91220 117195 91221
rect 118233 91220 118299 91221
rect 115790 91218 115796 91220
rect 113836 91216 113975 91218
rect 113836 91160 113914 91216
rect 113970 91160 113975 91216
rect 113836 91158 113975 91160
rect 115750 91158 115796 91218
rect 115860 91216 115907 91220
rect 117078 91218 117084 91220
rect 115902 91160 115907 91216
rect 113836 91156 113842 91158
rect 113909 91155 113975 91158
rect 115790 91156 115796 91158
rect 115860 91156 115907 91160
rect 117038 91158 117084 91218
rect 117148 91216 117195 91220
rect 118182 91218 118188 91220
rect 117190 91160 117195 91216
rect 117078 91156 117084 91158
rect 117148 91156 117195 91160
rect 118142 91158 118188 91218
rect 118252 91216 118299 91220
rect 118294 91160 118299 91216
rect 118182 91156 118188 91158
rect 118252 91156 118299 91160
rect 119654 91156 119660 91220
rect 119724 91218 119730 91220
rect 119981 91218 120047 91221
rect 119724 91216 120047 91218
rect 119724 91160 119986 91216
rect 120042 91160 120047 91216
rect 119724 91158 120047 91160
rect 119724 91156 119730 91158
rect 115841 91155 115907 91156
rect 117129 91155 117195 91156
rect 118233 91155 118299 91156
rect 119981 91155 120047 91158
rect 120206 91156 120212 91220
rect 120276 91218 120282 91220
rect 121361 91218 121427 91221
rect 120276 91216 121427 91218
rect 120276 91160 121366 91216
rect 121422 91160 121427 91216
rect 120276 91158 121427 91160
rect 120276 91156 120282 91158
rect 121361 91155 121427 91158
rect 122046 91156 122052 91220
rect 122116 91218 122122 91220
rect 122741 91218 122807 91221
rect 122116 91216 122807 91218
rect 122116 91160 122746 91216
rect 122802 91160 122807 91216
rect 122116 91158 122807 91160
rect 122116 91156 122122 91158
rect 122741 91155 122807 91158
rect 124029 91220 124095 91221
rect 124029 91216 124076 91220
rect 124140 91218 124146 91220
rect 124029 91160 124034 91216
rect 124029 91156 124076 91160
rect 124140 91158 124186 91218
rect 124140 91156 124146 91158
rect 126462 91156 126468 91220
rect 126532 91218 126538 91220
rect 126789 91218 126855 91221
rect 130745 91220 130811 91221
rect 133137 91220 133203 91221
rect 130694 91218 130700 91220
rect 126532 91216 126855 91218
rect 126532 91160 126794 91216
rect 126850 91160 126855 91216
rect 126532 91158 126855 91160
rect 130654 91158 130700 91218
rect 130764 91216 130811 91220
rect 133086 91218 133092 91220
rect 130806 91160 130811 91216
rect 126532 91156 126538 91158
rect 124029 91155 124095 91156
rect 126789 91155 126855 91158
rect 130694 91156 130700 91158
rect 130764 91156 130811 91160
rect 133046 91158 133092 91218
rect 133156 91216 133203 91220
rect 133198 91160 133203 91216
rect 133086 91156 133092 91158
rect 133156 91156 133203 91160
rect 134374 91156 134380 91220
rect 134444 91218 134450 91220
rect 134701 91218 134767 91221
rect 134444 91216 134767 91218
rect 134444 91160 134706 91216
rect 134762 91160 134767 91216
rect 134444 91158 134767 91160
rect 134444 91156 134450 91158
rect 130745 91155 130811 91156
rect 133137 91155 133203 91156
rect 134701 91155 134767 91158
rect 179270 91020 179276 91084
rect 179340 91082 179346 91084
rect 383561 91082 383627 91085
rect 408677 91082 408743 91085
rect 179340 91080 408743 91082
rect 179340 91024 383566 91080
rect 383622 91024 408682 91080
rect 408738 91024 408743 91080
rect 179340 91022 408743 91024
rect 179340 91020 179346 91022
rect 383561 91019 383627 91022
rect 408677 91019 408743 91022
rect 67449 90946 67515 90949
rect 214598 90946 214604 90948
rect 67449 90944 214604 90946
rect 67449 90888 67454 90944
rect 67510 90888 214604 90944
rect 67449 90886 214604 90888
rect 67449 90883 67515 90886
rect 214598 90884 214604 90886
rect 214668 90884 214674 90948
rect 57881 89722 57947 89725
rect 194041 89722 194107 89725
rect 57881 89720 194107 89722
rect 57881 89664 57886 89720
rect 57942 89664 194046 89720
rect 194102 89664 194107 89720
rect 57881 89662 194107 89664
rect 57881 89659 57947 89662
rect 194041 89659 194107 89662
rect 110229 88226 110295 88229
rect 166390 88226 166396 88228
rect 110229 88224 166396 88226
rect 110229 88168 110234 88224
rect 110290 88168 166396 88224
rect 110229 88166 166396 88168
rect 110229 88163 110295 88166
rect 166390 88164 166396 88166
rect 166460 88164 166466 88228
rect 97073 86866 97139 86869
rect 167678 86866 167684 86868
rect 97073 86864 167684 86866
rect 97073 86808 97078 86864
rect 97134 86808 167684 86864
rect 97073 86806 167684 86808
rect 97073 86803 97139 86806
rect 167678 86804 167684 86806
rect 167748 86804 167754 86868
rect 265566 86804 265572 86868
rect 265636 86866 265642 86868
rect 535453 86866 535519 86869
rect 265636 86864 535519 86866
rect 265636 86808 535458 86864
rect 535514 86808 535519 86864
rect 265636 86806 535519 86808
rect 265636 86804 265642 86806
rect 535453 86803 535519 86806
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect 55121 85506 55187 85509
rect 327901 85506 327967 85509
rect 55121 85504 327967 85506
rect 55121 85448 55126 85504
rect 55182 85448 327906 85504
rect 327962 85448 327967 85504
rect 55121 85446 327967 85448
rect 55121 85443 55187 85446
rect 327901 85443 327967 85446
rect 192477 84826 192543 84829
rect 307150 84826 307156 84828
rect 192477 84824 307156 84826
rect -960 84690 480 84780
rect 192477 84768 192482 84824
rect 192538 84768 307156 84824
rect 192477 84766 307156 84768
rect 192477 84763 192543 84766
rect 307150 84764 307156 84766
rect 307220 84764 307226 84828
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 106089 84146 106155 84149
rect 166206 84146 166212 84148
rect 106089 84144 166212 84146
rect 106089 84088 106094 84144
rect 106150 84088 166212 84144
rect 106089 84086 166212 84088
rect 106089 84083 106155 84086
rect 166206 84084 166212 84086
rect 166276 84084 166282 84148
rect 387006 84084 387012 84148
rect 387076 84146 387082 84148
rect 571374 84146 571380 84148
rect 387076 84086 571380 84146
rect 387076 84084 387082 84086
rect 571374 84084 571380 84086
rect 571444 84084 571450 84148
rect 101949 82786 102015 82789
rect 171726 82786 171732 82788
rect 101949 82784 171732 82786
rect 101949 82728 101954 82784
rect 102010 82728 171732 82784
rect 101949 82726 171732 82728
rect 101949 82723 102015 82726
rect 171726 82724 171732 82726
rect 171796 82724 171802 82788
rect 103421 81426 103487 81429
rect 170254 81426 170260 81428
rect 103421 81424 170260 81426
rect 103421 81368 103426 81424
rect 103482 81368 170260 81424
rect 103421 81366 170260 81368
rect 103421 81363 103487 81366
rect 170254 81364 170260 81366
rect 170324 81364 170330 81428
rect 17953 75170 18019 75173
rect 301630 75170 301636 75172
rect 17953 75168 301636 75170
rect 17953 75112 17958 75168
rect 18014 75112 301636 75168
rect 17953 75110 301636 75112
rect 17953 75107 18019 75110
rect 301630 75108 301636 75110
rect 301700 75108 301706 75172
rect 579981 72994 580047 72997
rect 583520 72994 584960 73084
rect 579981 72992 584960 72994
rect 579981 72936 579986 72992
rect 580042 72936 584960 72992
rect 579981 72934 584960 72936
rect 579981 72931 580047 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 13813 66874 13879 66877
rect 287646 66874 287652 66876
rect 13813 66872 287652 66874
rect 13813 66816 13818 66872
rect 13874 66816 287652 66872
rect 13813 66814 287652 66816
rect 13813 66811 13879 66814
rect 287646 66812 287652 66814
rect 287716 66812 287722 66876
rect 2773 64154 2839 64157
rect 305494 64154 305500 64156
rect 2773 64152 305500 64154
rect 2773 64096 2778 64152
rect 2834 64096 305500 64152
rect 2773 64094 305500 64096
rect 2773 64091 2839 64094
rect 305494 64092 305500 64094
rect 305564 64092 305570 64156
rect 67633 59938 67699 59941
rect 299974 59938 299980 59940
rect 67633 59936 299980 59938
rect 67633 59880 67638 59936
rect 67694 59880 299980 59936
rect 67633 59878 299980 59880
rect 67633 59875 67699 59878
rect 299974 59876 299980 59878
rect 300044 59876 300050 59940
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 69013 54498 69079 54501
rect 305678 54498 305684 54500
rect 69013 54496 305684 54498
rect 69013 54440 69018 54496
rect 69074 54440 305684 54496
rect 69013 54438 305684 54440
rect 69013 54435 69079 54438
rect 305678 54436 305684 54438
rect 305748 54436 305754 54500
rect 177062 51716 177068 51780
rect 177132 51778 177138 51780
rect 339493 51778 339559 51781
rect 177132 51776 339559 51778
rect 177132 51720 339498 51776
rect 339554 51720 339559 51776
rect 177132 51718 339559 51720
rect 177132 51716 177138 51718
rect 339493 51715 339559 51718
rect 176326 50220 176332 50284
rect 176396 50282 176402 50284
rect 313273 50282 313339 50285
rect 176396 50280 313339 50282
rect 176396 50224 313278 50280
rect 313334 50224 313339 50280
rect 176396 50222 313339 50224
rect 176396 50220 176402 50222
rect 313273 50219 313339 50222
rect 583753 46882 583819 46885
rect 583710 46880 583819 46882
rect 583710 46824 583758 46880
rect 583814 46824 583819 46880
rect 583710 46819 583819 46824
rect 583710 46474 583770 46819
rect 583342 46428 583770 46474
rect 583342 46414 584960 46428
rect 583342 46338 583402 46414
rect 583520 46338 584960 46414
rect 583342 46278 584960 46338
rect 11053 46202 11119 46205
rect 302734 46202 302740 46204
rect 11053 46200 302740 46202
rect 11053 46144 11058 46200
rect 11114 46144 302740 46200
rect 11053 46142 302740 46144
rect 11053 46139 11119 46142
rect 302734 46140 302740 46142
rect 302804 46140 302810 46204
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 175038 42060 175044 42124
rect 175108 42122 175114 42124
rect 336733 42122 336799 42125
rect 175108 42120 336799 42122
rect 175108 42064 336738 42120
rect 336794 42064 336799 42120
rect 175108 42062 336799 42064
rect 175108 42060 175114 42062
rect 336733 42059 336799 42062
rect 8293 40626 8359 40629
rect 283414 40626 283420 40628
rect 8293 40624 283420 40626
rect 8293 40568 8298 40624
rect 8354 40568 283420 40624
rect 8293 40566 283420 40568
rect 8293 40563 8359 40566
rect 283414 40564 283420 40566
rect 283484 40564 283490 40628
rect 55213 36546 55279 36549
rect 304206 36546 304212 36548
rect 55213 36544 304212 36546
rect 55213 36488 55218 36544
rect 55274 36488 304212 36544
rect 55213 36486 304212 36488
rect 55213 36483 55279 36486
rect 304206 36484 304212 36486
rect 304276 36484 304282 36548
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 179822 26964 179828 27028
rect 179892 27026 179898 27028
rect 287053 27026 287119 27029
rect 179892 27024 287119 27026
rect 179892 26968 287058 27024
rect 287114 26968 287119 27024
rect 179892 26966 287119 26968
rect 179892 26964 179898 26966
rect 287053 26963 287119 26966
rect 117313 26890 117379 26893
rect 253054 26890 253060 26892
rect 117313 26888 253060 26890
rect 117313 26832 117318 26888
rect 117374 26832 253060 26888
rect 117313 26830 253060 26832
rect 117313 26827 117379 26830
rect 253054 26828 253060 26830
rect 253124 26828 253130 26892
rect 285765 26890 285831 26893
rect 293902 26890 293908 26892
rect 285765 26888 293908 26890
rect 285765 26832 285770 26888
rect 285826 26832 293908 26888
rect 285765 26830 293908 26832
rect 285765 26827 285831 26830
rect 293902 26828 293908 26830
rect 293972 26828 293978 26892
rect 208158 24108 208164 24172
rect 208228 24170 208234 24172
rect 345013 24170 345079 24173
rect 208228 24168 345079 24170
rect 208228 24112 345018 24168
rect 345074 24112 345079 24168
rect 208228 24110 345079 24112
rect 208228 24108 208234 24110
rect 345013 24107 345079 24110
rect 583520 19818 584960 19908
rect 583342 19758 584960 19818
rect 583342 19682 583402 19758
rect 583520 19682 584960 19758
rect 583342 19668 584960 19682
rect 583342 19622 583586 19668
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 388294 19348 388300 19412
rect 388364 19410 388370 19412
rect 583526 19410 583586 19622
rect 388364 19350 583586 19410
rect 388364 19348 388370 19350
rect 77385 17234 77451 17237
rect 306966 17234 306972 17236
rect 77385 17232 306972 17234
rect 77385 17176 77390 17232
rect 77446 17176 306972 17232
rect 77385 17174 306972 17176
rect 77385 17171 77451 17174
rect 306966 17172 306972 17174
rect 307036 17172 307042 17236
rect 173750 15812 173756 15876
rect 173820 15874 173826 15876
rect 579613 15874 579679 15877
rect 173820 15872 579679 15874
rect 173820 15816 579618 15872
rect 579674 15816 579679 15872
rect 173820 15814 579679 15816
rect 173820 15812 173826 15814
rect 579613 15811 579679 15814
rect 580257 6626 580323 6629
rect 583520 6626 584960 6716
rect 580257 6624 584960 6626
rect -960 6490 480 6580
rect 580257 6568 580262 6624
rect 580318 6568 584960 6624
rect 580257 6566 584960 6568
rect 580257 6563 580323 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 259453 6354 259519 6357
rect 288934 6354 288940 6356
rect 259453 6352 288940 6354
rect 259453 6296 259458 6352
rect 259514 6296 288940 6352
rect 259453 6294 288940 6296
rect 259453 6291 259519 6294
rect 288934 6292 288940 6294
rect 289004 6292 289010 6356
rect 176510 6156 176516 6220
rect 176580 6218 176586 6220
rect 304349 6218 304415 6221
rect 176580 6216 304415 6218
rect 176580 6160 304354 6216
rect 304410 6160 304415 6216
rect 176580 6158 304415 6160
rect 176580 6156 176586 6158
rect 304349 6155 304415 6158
rect 32397 4858 32463 4861
rect 301446 4858 301452 4860
rect 32397 4856 301452 4858
rect 32397 4800 32402 4856
rect 32458 4800 301452 4856
rect 32397 4798 301452 4800
rect 32397 4795 32463 4798
rect 301446 4796 301452 4798
rect 301516 4796 301522 4860
rect 255865 3500 255931 3501
rect 255814 3436 255820 3500
rect 255884 3498 255931 3500
rect 257061 3498 257127 3501
rect 257838 3498 257844 3500
rect 255884 3496 255976 3498
rect 255926 3440 255976 3496
rect 255884 3438 255976 3440
rect 257061 3496 257844 3498
rect 257061 3440 257066 3496
rect 257122 3440 257844 3496
rect 257061 3438 257844 3440
rect 255884 3436 255931 3438
rect 255865 3435 255931 3436
rect 257061 3435 257127 3438
rect 257838 3436 257844 3438
rect 257908 3436 257914 3500
rect 271229 3498 271295 3501
rect 275134 3498 275140 3500
rect 271229 3496 275140 3498
rect 271229 3440 271234 3496
rect 271290 3440 275140 3496
rect 271229 3438 275140 3440
rect 271229 3435 271295 3438
rect 275134 3436 275140 3438
rect 275204 3436 275210 3500
rect 337326 3436 337332 3500
rect 337396 3498 337402 3500
rect 338665 3498 338731 3501
rect 337396 3496 338731 3498
rect 337396 3440 338670 3496
rect 338726 3440 338731 3496
rect 337396 3438 338731 3440
rect 337396 3436 337402 3438
rect 338665 3435 338731 3438
rect 219198 3300 219204 3364
rect 219268 3362 219274 3364
rect 219268 3302 238770 3362
rect 219268 3300 219274 3302
rect 238710 3226 238770 3302
rect 264094 3300 264100 3364
rect 264164 3362 264170 3364
rect 278313 3362 278379 3365
rect 264164 3360 278379 3362
rect 264164 3304 278318 3360
rect 278374 3304 278379 3360
rect 264164 3302 278379 3304
rect 264164 3300 264170 3302
rect 278313 3299 278379 3302
rect 296069 3362 296135 3365
rect 327022 3362 327028 3364
rect 296069 3360 327028 3362
rect 296069 3304 296074 3360
rect 296130 3304 327028 3360
rect 296069 3302 327028 3304
rect 296069 3299 296135 3302
rect 327022 3300 327028 3302
rect 327092 3300 327098 3364
rect 242893 3226 242959 3229
rect 238710 3224 242959 3226
rect 238710 3168 242898 3224
rect 242954 3168 242959 3224
rect 238710 3166 242959 3168
rect 242893 3163 242959 3166
<< obsm3 >>
rect 68800 171594 164756 174600
rect 68800 171534 164694 171594
rect 68800 129304 164756 171534
rect 68816 129244 164756 129304
rect 68800 128080 164756 129244
rect 68816 128020 164756 128080
rect 68800 126312 164756 128020
rect 68816 126252 164756 126312
rect 68800 125224 164756 126252
rect 68816 125164 164756 125224
rect 68800 123592 164756 125164
rect 68816 123532 164756 123592
rect 68800 122640 164756 123532
rect 68816 122580 164756 122640
rect 68800 120872 164756 122580
rect 68816 120812 164756 120872
rect 68800 111754 164756 120812
rect 68800 111694 164694 111754
rect 68800 110122 164756 111694
rect 68800 110062 164694 110122
rect 68800 108762 164756 110062
rect 68800 108702 164694 108762
rect 68800 102376 164756 108702
rect 68816 102316 164756 102376
rect 68800 100744 164756 102316
rect 68816 100684 164756 100744
rect 68800 95100 164756 100684
<< via3 >>
rect 295932 702476 295996 702540
rect 121500 579668 121564 579732
rect 579660 511260 579724 511324
rect 579660 510580 579724 510644
rect 295932 365740 295996 365804
rect 570092 364380 570156 364444
rect 69060 363020 69124 363084
rect 294092 358804 294156 358868
rect 292436 356220 292500 356284
rect 335860 356084 335924 356148
rect 167500 354860 167564 354924
rect 293172 354860 293236 354924
rect 171732 354724 171796 354788
rect 292620 352956 292684 353020
rect 295380 352276 295444 352340
rect 177068 350100 177132 350164
rect 293908 347516 293972 347580
rect 295748 343436 295812 343500
rect 295748 341396 295812 341460
rect 173756 339220 173820 339284
rect 179276 334460 179340 334524
rect 175044 330380 175108 330444
rect 176332 323580 176396 323644
rect 176516 316780 176580 316844
rect 161244 311884 161308 311948
rect 292620 311884 292684 311948
rect 388484 311068 388548 311132
rect 387012 301412 387076 301476
rect 149652 299432 149716 299436
rect 149652 299376 149702 299432
rect 149702 299376 149716 299432
rect 149652 299372 149716 299376
rect 293172 298692 293236 298756
rect 167684 298284 167748 298348
rect 149652 298148 149716 298212
rect 66116 297332 66180 297396
rect 166212 296924 166276 296988
rect 158484 296848 158548 296852
rect 158484 296792 158498 296848
rect 158498 296792 158548 296848
rect 158484 296788 158548 296792
rect 574692 294476 574756 294540
rect 170260 294068 170324 294132
rect 126100 292980 126164 293044
rect 146892 292844 146956 292908
rect 64644 292572 64708 292636
rect 568620 285636 568684 285700
rect 571564 284820 571628 284884
rect 178540 283188 178604 283252
rect 390692 280468 390756 280532
rect 569540 278700 569604 278764
rect 385540 276252 385604 276316
rect 389772 276116 389836 276180
rect 293172 275980 293236 276044
rect 390508 275632 390572 275636
rect 390508 275576 390522 275632
rect 390522 275576 390572 275632
rect 390508 275572 390572 275576
rect 502012 275572 502076 275636
rect 502012 274620 502076 274684
rect 568620 274484 568684 274548
rect 390508 274212 390572 274276
rect 121500 272716 121564 272780
rect 390508 272444 390572 272508
rect 171916 267820 171980 267884
rect 161980 266324 162044 266388
rect 169156 265100 169220 265164
rect 59124 263664 59188 263668
rect 59124 263608 59174 263664
rect 59174 263608 59188 263664
rect 59124 263604 59188 263608
rect 120028 257212 120092 257276
rect 156460 257272 156524 257276
rect 156460 257216 156510 257272
rect 156510 257216 156524 257272
rect 156460 257212 156524 257216
rect 124812 255036 124876 255100
rect 61884 254084 61948 254148
rect 120580 254220 120644 254284
rect 142660 248372 142724 248436
rect 296668 248372 296732 248436
rect 171732 247012 171796 247076
rect 63356 245788 63420 245852
rect 67404 246196 67468 246260
rect 167500 244836 167564 244900
rect 571380 244292 571444 244356
rect 69060 242932 69124 242996
rect 179828 242932 179892 242996
rect 292620 242932 292684 242996
rect 120028 242524 120092 242588
rect 63172 241708 63236 241772
rect 126100 242116 126164 242180
rect 66116 241436 66180 241500
rect 70532 240212 70596 240276
rect 61884 240136 61948 240140
rect 61884 240080 61898 240136
rect 61898 240080 61948 240136
rect 61884 240076 61948 240080
rect 288940 240076 289004 240140
rect 294092 240076 294156 240140
rect 120580 239668 120644 239732
rect 161980 239396 162044 239460
rect 178540 239396 178604 239460
rect 149652 238716 149716 238780
rect 389772 238716 389836 238780
rect 119844 238580 119908 238644
rect 293172 238444 293236 238508
rect 119660 238308 119724 238372
rect 208164 237356 208228 237420
rect 167684 235860 167748 235924
rect 146892 235180 146956 235244
rect 161244 234500 161308 234564
rect 296484 234364 296548 234428
rect 166212 233140 166276 233204
rect 158484 232596 158548 232660
rect 322060 232460 322124 232524
rect 292620 230420 292684 230484
rect 59124 229740 59188 229804
rect 63172 228924 63236 228988
rect 161980 228788 162044 228852
rect 265572 227760 265636 227764
rect 265572 227704 265622 227760
rect 265622 227704 265636 227760
rect 265572 227700 265636 227704
rect 291700 226204 291764 226268
rect 70900 224844 70964 224908
rect 63356 224708 63420 224772
rect 387012 224572 387076 224636
rect 64644 222804 64708 222868
rect 388300 222124 388364 222188
rect 255268 218588 255332 218652
rect 142660 216548 142724 216612
rect 388484 213888 388548 213892
rect 388484 213832 388498 213888
rect 388498 213832 388548 213888
rect 388484 213828 388548 213832
rect 171916 211788 171980 211852
rect 67404 207572 67468 207636
rect 263548 204852 263612 204916
rect 256740 203492 256804 203556
rect 156460 200772 156524 200836
rect 571564 200772 571628 200836
rect 124812 200636 124876 200700
rect 269068 195196 269132 195260
rect 337332 195196 337396 195260
rect 275140 193836 275204 193900
rect 571564 193836 571628 193900
rect 266308 191116 266372 191180
rect 256924 190980 256988 191044
rect 264100 189756 264164 189820
rect 254532 189620 254596 189684
rect 324268 189076 324332 189140
rect 252508 188396 252572 188460
rect 259500 188260 259564 188324
rect 326660 187172 326724 187236
rect 265020 187036 265084 187100
rect 320220 186900 320284 186964
rect 328500 184996 328564 185060
rect 331812 184180 331876 184244
rect 171180 182956 171244 183020
rect 261156 182956 261220 183020
rect 327580 182820 327644 182884
rect 167500 181596 167564 181660
rect 260788 181596 260852 181660
rect 251220 181460 251284 181524
rect 262260 181324 262324 181388
rect 332548 179964 332612 180028
rect 249012 179148 249076 179212
rect 166396 178060 166460 178124
rect 273852 178060 273916 178124
rect 97028 177924 97092 177988
rect 100708 177652 100772 177716
rect 99420 177516 99484 177580
rect 103284 177516 103348 177580
rect 110644 177576 110708 177580
rect 110644 177520 110694 177576
rect 110694 177520 110708 177576
rect 110644 177516 110708 177520
rect 112116 177516 112180 177580
rect 115796 177576 115860 177580
rect 115796 177520 115846 177576
rect 115846 177520 115860 177576
rect 115796 177516 115860 177520
rect 119660 177516 119724 177580
rect 120764 177516 120828 177580
rect 125732 177516 125796 177580
rect 127020 177516 127084 177580
rect 130700 177576 130764 177580
rect 130700 177520 130750 177576
rect 130750 177520 130764 177576
rect 130700 177516 130764 177520
rect 249196 177516 249260 177580
rect 259684 177380 259748 177444
rect 327028 177244 327092 177308
rect 109540 176972 109604 177036
rect 113220 176972 113284 177036
rect 131988 177032 132052 177036
rect 131988 176976 132038 177032
rect 132038 176976 132052 177032
rect 131988 176972 132052 176976
rect 101996 176836 102060 176900
rect 104572 176760 104636 176764
rect 104572 176704 104622 176760
rect 104622 176704 104636 176760
rect 104572 176700 104636 176704
rect 106964 176760 107028 176764
rect 106964 176704 107014 176760
rect 107014 176704 107028 176760
rect 106964 176700 107028 176704
rect 108068 176760 108132 176764
rect 108068 176704 108118 176760
rect 108118 176704 108132 176760
rect 108068 176700 108132 176704
rect 118372 176760 118436 176764
rect 118372 176704 118422 176760
rect 118422 176704 118436 176760
rect 118372 176700 118436 176704
rect 121868 176700 121932 176764
rect 122972 176760 123036 176764
rect 122972 176704 123022 176760
rect 123022 176704 123036 176760
rect 122972 176700 123036 176704
rect 129412 176760 129476 176764
rect 129412 176704 129462 176760
rect 129462 176704 129476 176760
rect 129412 176700 129476 176704
rect 133092 176760 133156 176764
rect 133092 176704 133142 176760
rect 133142 176704 133156 176760
rect 133092 176700 133156 176704
rect 135668 176760 135732 176764
rect 135668 176704 135718 176760
rect 135718 176704 135732 176760
rect 135668 176700 135732 176704
rect 148180 176760 148244 176764
rect 148180 176704 148230 176760
rect 148230 176704 148244 176760
rect 148180 176700 148244 176704
rect 158852 176700 158916 176764
rect 321324 176700 321388 176764
rect 128124 176428 128188 176492
rect 255452 176428 255516 176492
rect 387012 176292 387076 176356
rect 252692 176020 252756 176084
rect 328684 176020 328748 176084
rect 257844 175884 257908 175948
rect 271092 175884 271156 175948
rect 116900 175672 116964 175676
rect 116900 175616 116950 175672
rect 116950 175616 116964 175672
rect 116900 175612 116964 175616
rect 124444 175672 124508 175676
rect 124444 175616 124494 175672
rect 124494 175616 124508 175672
rect 124444 175612 124508 175616
rect 134380 175672 134444 175676
rect 134380 175616 134430 175672
rect 134430 175616 134444 175672
rect 134380 175612 134444 175616
rect 342300 175884 342364 175948
rect 387564 175884 387628 175948
rect 114324 175476 114388 175540
rect 166212 175476 166276 175540
rect 98316 175400 98380 175404
rect 98316 175344 98366 175400
rect 98366 175344 98380 175400
rect 98316 175340 98380 175344
rect 105676 175340 105740 175404
rect 167684 175340 167748 175404
rect 306972 175204 307036 175268
rect 249380 174660 249444 174724
rect 254532 174252 254596 174316
rect 249196 173708 249260 173772
rect 326660 173844 326724 173908
rect 569540 173844 569604 173908
rect 321324 172076 321388 172140
rect 170260 171668 170324 171732
rect 321324 170308 321388 170372
rect 252508 170036 252572 170100
rect 257844 168540 257908 168604
rect 166212 164324 166276 164388
rect 269068 163100 269132 163164
rect 261156 162964 261220 163028
rect 328684 162692 328748 162756
rect 331812 161196 331876 161260
rect 256924 161060 256988 161124
rect 171180 160108 171244 160172
rect 265020 159564 265084 159628
rect 167684 158748 167748 158812
rect 262260 157932 262324 157996
rect 307340 157388 307404 157452
rect 252692 157252 252756 157316
rect 324268 155484 324332 155548
rect 166396 154532 166460 154596
rect 255452 150180 255516 150244
rect 307156 150180 307220 150244
rect 306972 149636 307036 149700
rect 322060 148684 322124 148748
rect 251956 148140 252020 148204
rect 321508 148004 321572 148068
rect 251220 147868 251284 147932
rect 251772 146236 251836 146300
rect 255820 146236 255884 146300
rect 266308 145556 266372 145620
rect 307340 145556 307404 145620
rect 328500 145556 328564 145620
rect 259684 142564 259748 142628
rect 307708 142020 307772 142084
rect 256740 141748 256804 141812
rect 255268 140796 255332 140860
rect 307708 139980 307772 140044
rect 305500 139708 305564 139772
rect 253244 138348 253308 138412
rect 332548 138620 332612 138684
rect 259500 138212 259564 138276
rect 263548 137940 263612 138004
rect 171916 136852 171980 136916
rect 260972 136580 261036 136644
rect 307156 134404 307220 134468
rect 306972 133996 307036 134060
rect 166396 133860 166460 133924
rect 214420 132636 214484 132700
rect 299980 132636 300044 132700
rect 166212 131412 166276 131476
rect 170260 130052 170324 130116
rect 171732 129916 171796 129980
rect 257844 128964 257908 129028
rect 342300 128964 342364 129028
rect 301452 128420 301516 128484
rect 251956 127604 252020 127668
rect 167684 127196 167748 127260
rect 287652 125836 287716 125900
rect 327580 121408 327644 121412
rect 327580 121352 327594 121408
rect 327594 121352 327644 121408
rect 327580 121348 327644 121352
rect 385540 121348 385604 121412
rect 304212 117812 304276 117876
rect 387196 116452 387260 116516
rect 389772 115092 389836 115156
rect 301636 113596 301700 113660
rect 283420 112100 283484 112164
rect 387564 112372 387628 112436
rect 251772 111148 251836 111212
rect 387012 109652 387076 109716
rect 570092 109652 570156 109716
rect 305684 105844 305748 105908
rect 324268 104756 324332 104820
rect 295380 104076 295444 104140
rect 335860 102172 335924 102236
rect 214604 101492 214668 101556
rect 271092 101356 271156 101420
rect 302740 99588 302804 99652
rect 273852 97820 273916 97884
rect 167316 97140 167380 97204
rect 579660 97140 579724 97204
rect 307156 97004 307220 97068
rect 324452 96596 324516 96660
rect 322060 96460 322124 96524
rect 324452 96324 324516 96388
rect 387196 96324 387260 96388
rect 571564 96324 571628 96388
rect 219204 95916 219268 95980
rect 389772 96188 389836 96252
rect 112326 94752 112390 94756
rect 112326 94696 112350 94752
rect 112350 94696 112390 94752
rect 112326 94692 112390 94696
rect 113142 94752 113206 94756
rect 113142 94696 113178 94752
rect 113178 94696 113206 94752
rect 113142 94692 113206 94696
rect 119398 94692 119462 94756
rect 119844 94692 119908 94756
rect 123206 94752 123270 94756
rect 123206 94696 123262 94752
rect 123262 94696 123270 94752
rect 123206 94692 123270 94696
rect 151308 94692 151372 94756
rect 151630 94692 151694 94756
rect 151902 94752 151966 94756
rect 151902 94696 151910 94752
rect 151910 94696 151966 94752
rect 151902 94692 151966 94696
rect 167500 94420 167564 94484
rect 116716 93740 116780 93804
rect 121684 93664 121748 93668
rect 121684 93608 121734 93664
rect 121734 93608 121748 93664
rect 121684 93604 121748 93608
rect 169156 93740 169220 93804
rect 171916 93604 171980 93668
rect 574692 93604 574756 93668
rect 93900 93528 93964 93532
rect 93900 93472 93950 93528
rect 93950 93472 93964 93528
rect 93900 93468 93964 93472
rect 107700 93528 107764 93532
rect 107700 93472 107750 93528
rect 107750 93472 107764 93528
rect 107700 93468 107764 93472
rect 151492 93528 151556 93532
rect 151492 93472 151542 93528
rect 151542 93472 151556 93528
rect 151492 93468 151556 93472
rect 110092 93256 110156 93260
rect 110092 93200 110142 93256
rect 110142 93200 110156 93256
rect 110092 93196 110156 93200
rect 128124 93256 128188 93260
rect 128124 93200 128174 93256
rect 128174 93200 128188 93256
rect 128124 93196 128188 93200
rect 324268 93256 324332 93260
rect 324268 93200 324318 93256
rect 324318 93200 324332 93256
rect 324268 93196 324332 93200
rect 214420 93060 214484 93124
rect 85620 92380 85684 92444
rect 87092 92380 87156 92444
rect 88932 92440 88996 92444
rect 88932 92384 88982 92440
rect 88982 92384 88996 92440
rect 88932 92380 88996 92384
rect 99604 92380 99668 92444
rect 106780 92380 106844 92444
rect 109172 92380 109236 92444
rect 111196 92380 111260 92444
rect 114140 92440 114204 92444
rect 114140 92384 114190 92440
rect 114190 92384 114204 92440
rect 114140 92380 114204 92384
rect 118004 92440 118068 92444
rect 118004 92384 118054 92440
rect 118054 92384 118068 92440
rect 118004 92380 118068 92384
rect 124444 92440 124508 92444
rect 124444 92384 124494 92440
rect 124494 92384 124508 92440
rect 124444 92380 124508 92384
rect 125364 92440 125428 92444
rect 125364 92384 125414 92440
rect 125414 92384 125428 92440
rect 125364 92380 125428 92384
rect 125732 92440 125796 92444
rect 125732 92384 125782 92440
rect 125782 92384 125796 92440
rect 125732 92380 125796 92384
rect 129412 92440 129476 92444
rect 129412 92384 129462 92440
rect 129462 92384 129476 92440
rect 129412 92380 129476 92384
rect 135668 92440 135732 92444
rect 135668 92384 135718 92440
rect 135718 92384 135732 92440
rect 135668 92380 135732 92384
rect 115428 92244 115492 92308
rect 167316 92244 167380 92308
rect 151676 92168 151740 92172
rect 151676 92112 151726 92168
rect 151726 92112 151740 92168
rect 151676 92108 151740 92112
rect 115060 91700 115124 91764
rect 104204 91624 104268 91628
rect 104204 91568 104254 91624
rect 104254 91568 104268 91624
rect 104204 91564 104268 91568
rect 131988 91564 132052 91628
rect 151308 91624 151372 91628
rect 151308 91568 151358 91624
rect 151358 91568 151372 91624
rect 151308 91564 151372 91568
rect 98500 91428 98564 91492
rect 101812 91488 101876 91492
rect 101812 91432 101862 91488
rect 101862 91432 101876 91488
rect 101812 91428 101876 91432
rect 122788 91428 122852 91492
rect 98132 91292 98196 91356
rect 101628 91292 101692 91356
rect 102916 91292 102980 91356
rect 105124 91292 105188 91356
rect 119844 91352 119908 91356
rect 119844 91296 119894 91352
rect 119894 91296 119908 91352
rect 119844 91292 119908 91296
rect 120580 91292 120644 91356
rect 126652 91292 126716 91356
rect 74764 91156 74828 91220
rect 84332 91156 84396 91220
rect 86724 91156 86788 91220
rect 90220 91156 90284 91220
rect 91324 91156 91388 91220
rect 92612 91156 92676 91220
rect 95004 91156 95068 91220
rect 96108 91156 96172 91220
rect 97028 91216 97092 91220
rect 97028 91160 97078 91216
rect 97078 91160 97092 91216
rect 97028 91156 97092 91160
rect 97212 91156 97276 91220
rect 99236 91216 99300 91220
rect 99236 91160 99250 91216
rect 99250 91160 99300 91216
rect 99236 91156 99300 91160
rect 100524 91216 100588 91220
rect 100524 91160 100574 91216
rect 100574 91160 100588 91216
rect 100524 91156 100588 91160
rect 101996 91216 102060 91220
rect 101996 91160 102010 91216
rect 102010 91160 102060 91216
rect 101996 91156 102060 91160
rect 103284 91156 103348 91220
rect 104572 91156 104636 91220
rect 106044 91216 106108 91220
rect 106044 91160 106094 91216
rect 106094 91160 106108 91216
rect 106044 91156 106108 91160
rect 106412 91156 106476 91220
rect 108068 91156 108132 91220
rect 109540 91156 109604 91220
rect 110644 91156 110708 91220
rect 111932 91156 111996 91220
rect 113772 91156 113836 91220
rect 115796 91216 115860 91220
rect 115796 91160 115846 91216
rect 115846 91160 115860 91216
rect 115796 91156 115860 91160
rect 117084 91216 117148 91220
rect 117084 91160 117134 91216
rect 117134 91160 117148 91216
rect 117084 91156 117148 91160
rect 118188 91216 118252 91220
rect 118188 91160 118238 91216
rect 118238 91160 118252 91216
rect 118188 91156 118252 91160
rect 119660 91156 119724 91220
rect 120212 91156 120276 91220
rect 122052 91156 122116 91220
rect 124076 91216 124140 91220
rect 124076 91160 124090 91216
rect 124090 91160 124140 91216
rect 124076 91156 124140 91160
rect 126468 91156 126532 91220
rect 130700 91216 130764 91220
rect 130700 91160 130750 91216
rect 130750 91160 130764 91216
rect 130700 91156 130764 91160
rect 133092 91216 133156 91220
rect 133092 91160 133142 91216
rect 133142 91160 133156 91216
rect 133092 91156 133156 91160
rect 134380 91156 134444 91220
rect 179276 91020 179340 91084
rect 214604 90884 214668 90948
rect 166396 88164 166460 88228
rect 167684 86804 167748 86868
rect 265572 86804 265636 86868
rect 307156 84764 307220 84828
rect 166212 84084 166276 84148
rect 387012 84084 387076 84148
rect 571380 84084 571444 84148
rect 171732 82724 171796 82788
rect 170260 81364 170324 81428
rect 301636 75108 301700 75172
rect 287652 66812 287716 66876
rect 305500 64092 305564 64156
rect 299980 59876 300044 59940
rect 305684 54436 305748 54500
rect 177068 51716 177132 51780
rect 176332 50220 176396 50284
rect 302740 46140 302804 46204
rect 175044 42060 175108 42124
rect 283420 40564 283484 40628
rect 304212 36484 304276 36548
rect 179828 26964 179892 27028
rect 253060 26828 253124 26892
rect 293908 26828 293972 26892
rect 208164 24108 208228 24172
rect 388300 19348 388364 19412
rect 306972 17172 307036 17236
rect 173756 15812 173820 15876
rect 288940 6292 289004 6356
rect 176516 6156 176580 6220
rect 301452 4796 301516 4860
rect 255820 3496 255884 3500
rect 255820 3440 255870 3496
rect 255870 3440 255884 3496
rect 255820 3436 255884 3440
rect 257844 3436 257908 3500
rect 275140 3436 275204 3500
rect 337332 3436 337396 3500
rect 219204 3300 219268 3364
rect 264100 3300 264164 3364
rect 327028 3300 327092 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69059 363084 69125 363085
rect 69059 363020 69060 363084
rect 69124 363020 69125 363084
rect 69059 363019 69125 363020
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64643 292636 64709 292637
rect 64643 292572 64644 292636
rect 64708 292572 64709 292636
rect 64643 292571 64709 292572
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 59123 263668 59189 263669
rect 59123 263604 59124 263668
rect 59188 263604 59189 263668
rect 59123 263603 59189 263604
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 59126 229805 59186 263603
rect 60294 241954 60914 277398
rect 61883 254148 61949 254149
rect 61883 254084 61884 254148
rect 61948 254084 61949 254148
rect 61883 254083 61949 254084
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 59123 229804 59189 229805
rect 59123 229740 59124 229804
rect 59188 229740 59189 229804
rect 59123 229739 59189 229740
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 205954 60914 241398
rect 61886 240141 61946 254083
rect 63355 245852 63421 245853
rect 63355 245788 63356 245852
rect 63420 245788 63421 245852
rect 63355 245787 63421 245788
rect 63171 241772 63237 241773
rect 63171 241708 63172 241772
rect 63236 241708 63237 241772
rect 63171 241707 63237 241708
rect 61883 240140 61949 240141
rect 61883 240076 61884 240140
rect 61948 240076 61949 240140
rect 61883 240075 61949 240076
rect 63174 228989 63234 241707
rect 63171 228988 63237 228989
rect 63171 228924 63172 228988
rect 63236 228924 63237 228988
rect 63171 228923 63237 228924
rect 63358 224773 63418 245787
rect 63355 224772 63421 224773
rect 63355 224708 63356 224772
rect 63420 224708 63421 224772
rect 63355 224707 63421 224708
rect 64646 222869 64706 292571
rect 64794 282454 65414 317898
rect 66115 297396 66181 297397
rect 66115 297332 66116 297396
rect 66180 297332 66181 297396
rect 66115 297331 66181 297332
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64643 222868 64709 222869
rect 64643 222804 64644 222868
rect 64708 222804 64709 222868
rect 64643 222803 64709 222804
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 210454 65414 245898
rect 66118 241501 66178 297331
rect 67403 246260 67469 246261
rect 67403 246196 67404 246260
rect 67468 246196 67469 246260
rect 67403 246195 67469 246196
rect 66115 241500 66181 241501
rect 66115 241436 66116 241500
rect 66180 241436 66181 241500
rect 66115 241435 66181 241436
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 67406 207637 67466 246195
rect 69062 242997 69122 363019
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 294000 69914 322398
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 294000 74414 326898
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 294000 78914 295398
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 294000 83414 299898
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 294000 87914 304398
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 294000 92414 308898
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 294000 96914 313398
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 294000 101414 317898
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 294000 105914 322398
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 294000 110414 326898
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 294000 114914 295398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 121499 579732 121565 579733
rect 121499 579668 121500 579732
rect 121564 579668 121565 579732
rect 121499 579667 121565 579668
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 294000 119414 299898
rect 121502 272781 121562 579667
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 121499 272780 121565 272781
rect 121499 272716 121500 272780
rect 121564 272716 121565 272780
rect 121499 272715 121565 272716
rect 123294 268954 123914 304398
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 126099 293044 126165 293045
rect 126099 292980 126100 293044
rect 126164 292980 126165 293044
rect 126099 292979 126165 292980
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 89568 259954 89888 259986
rect 89568 259718 89610 259954
rect 89846 259718 89888 259954
rect 89568 259634 89888 259718
rect 89568 259398 89610 259634
rect 89846 259398 89888 259634
rect 89568 259366 89888 259398
rect 120027 257276 120093 257277
rect 120027 257212 120028 257276
rect 120092 257212 120093 257276
rect 120027 257211 120093 257212
rect 74208 255454 74528 255486
rect 74208 255218 74250 255454
rect 74486 255218 74528 255454
rect 74208 255134 74528 255218
rect 74208 254898 74250 255134
rect 74486 254898 74528 255134
rect 74208 254866 74528 254898
rect 104928 255454 105248 255486
rect 104928 255218 104970 255454
rect 105206 255218 105248 255454
rect 104928 255134 105248 255218
rect 104928 254898 104970 255134
rect 105206 254898 105248 255134
rect 104928 254866 105248 254898
rect 120030 248430 120090 257211
rect 120579 254284 120645 254285
rect 120579 254220 120580 254284
rect 120644 254220 120645 254284
rect 120579 254219 120645 254220
rect 119662 248370 120090 248430
rect 69059 242996 69125 242997
rect 69059 242932 69060 242996
rect 69124 242932 69125 242996
rect 69059 242931 69125 242932
rect 70531 240276 70597 240277
rect 70531 240212 70532 240276
rect 70596 240212 70597 240276
rect 70531 240211 70597 240212
rect 70534 238770 70594 240211
rect 70534 238710 70962 238770
rect 69294 214954 69914 238000
rect 70902 224909 70962 238710
rect 119662 238373 119722 248370
rect 120027 242588 120093 242589
rect 120027 242524 120028 242588
rect 120092 242524 120093 242588
rect 120027 242523 120093 242524
rect 120030 238770 120090 242523
rect 120582 239733 120642 254219
rect 120579 239732 120645 239733
rect 120579 239668 120580 239732
rect 120644 239668 120645 239732
rect 120579 239667 120645 239668
rect 119846 238710 120090 238770
rect 119846 238645 119906 238710
rect 119843 238644 119909 238645
rect 119843 238580 119844 238644
rect 119908 238580 119909 238644
rect 119843 238579 119909 238580
rect 119659 238372 119725 238373
rect 119659 238308 119660 238372
rect 119724 238308 119725 238372
rect 119659 238307 119725 238308
rect 70899 224908 70965 224909
rect 70899 224844 70900 224908
rect 70964 224844 70965 224908
rect 70899 224843 70965 224844
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 67403 207636 67469 207637
rect 67403 207572 67404 207636
rect 67468 207572 67469 207636
rect 67403 207571 67469 207572
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 176600 69914 178398
rect 73794 219454 74414 238000
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 176600 74414 182898
rect 78294 223954 78914 238000
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 176600 78914 187398
rect 82794 228454 83414 238000
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 176600 83414 191898
rect 87294 232954 87914 238000
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 176600 87914 196398
rect 91794 237454 92414 238000
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 176600 92414 200898
rect 105294 214954 105914 238000
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 97027 177988 97093 177989
rect 97027 177924 97028 177988
rect 97092 177924 97093 177988
rect 97027 177923 97093 177924
rect 97030 175130 97090 177923
rect 100707 177716 100773 177717
rect 100707 177652 100708 177716
rect 100772 177652 100773 177716
rect 100707 177651 100773 177652
rect 99419 177580 99485 177581
rect 99419 177516 99420 177580
rect 99484 177516 99485 177580
rect 99419 177515 99485 177516
rect 98315 175404 98381 175405
rect 98315 175340 98316 175404
rect 98380 175340 98381 175404
rect 98315 175339 98381 175340
rect 96960 175070 97090 175130
rect 98318 175130 98378 175339
rect 99422 175130 99482 177515
rect 98318 175070 98380 175130
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 96960 174494 97020 175070
rect 98320 174494 98380 175070
rect 99408 175070 99482 175130
rect 100710 175130 100770 177651
rect 103283 177580 103349 177581
rect 103283 177516 103284 177580
rect 103348 177516 103349 177580
rect 103283 177515 103349 177516
rect 101995 176900 102061 176901
rect 101995 176836 101996 176900
rect 102060 176836 102061 176900
rect 101995 176835 102061 176836
rect 101998 175130 102058 176835
rect 100710 175070 100828 175130
rect 99408 174494 99468 175070
rect 100768 174494 100828 175070
rect 101992 175070 102058 175130
rect 103286 175130 103346 177515
rect 104571 176764 104637 176765
rect 104571 176700 104572 176764
rect 104636 176700 104637 176764
rect 104571 176699 104637 176700
rect 104574 175130 104634 176699
rect 105294 176600 105914 178398
rect 109794 219454 110414 238000
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109539 177036 109605 177037
rect 109539 176972 109540 177036
rect 109604 176972 109605 177036
rect 109539 176971 109605 176972
rect 106963 176764 107029 176765
rect 106963 176700 106964 176764
rect 107028 176700 107029 176764
rect 106963 176699 107029 176700
rect 108067 176764 108133 176765
rect 108067 176700 108068 176764
rect 108132 176700 108133 176764
rect 108067 176699 108133 176700
rect 105675 175404 105741 175405
rect 105675 175340 105676 175404
rect 105740 175340 105741 175404
rect 105675 175339 105741 175340
rect 105678 175130 105738 175339
rect 103286 175070 103412 175130
rect 104574 175070 104636 175130
rect 101992 174494 102052 175070
rect 103352 174494 103412 175070
rect 104576 174494 104636 175070
rect 105664 175070 105738 175130
rect 106966 175130 107026 176699
rect 108070 175130 108130 176699
rect 109542 175130 109602 176971
rect 109794 176600 110414 182898
rect 114294 223954 114914 238000
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 110643 177580 110709 177581
rect 110643 177516 110644 177580
rect 110708 177516 110709 177580
rect 110643 177515 110709 177516
rect 112115 177580 112181 177581
rect 112115 177516 112116 177580
rect 112180 177516 112181 177580
rect 112115 177515 112181 177516
rect 106966 175070 107084 175130
rect 108070 175070 108172 175130
rect 105664 174494 105724 175070
rect 107024 174494 107084 175070
rect 108112 174494 108172 175070
rect 109472 175070 109602 175130
rect 110646 175130 110706 177515
rect 112118 175130 112178 177515
rect 113219 177036 113285 177037
rect 113219 176972 113220 177036
rect 113284 176972 113285 177036
rect 113219 176971 113285 176972
rect 113222 175130 113282 176971
rect 114294 176600 114914 187398
rect 118794 228454 119414 238000
rect 118794 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 119414 228454
rect 118794 228134 119414 228218
rect 118794 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 119414 228134
rect 118794 192454 119414 227898
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 115795 177580 115861 177581
rect 115795 177516 115796 177580
rect 115860 177516 115861 177580
rect 115795 177515 115861 177516
rect 114323 175540 114389 175541
rect 114323 175476 114324 175540
rect 114388 175476 114389 175540
rect 114323 175475 114389 175476
rect 110646 175070 110756 175130
rect 109472 174494 109532 175070
rect 110696 174494 110756 175070
rect 112056 175070 112178 175130
rect 113144 175070 113282 175130
rect 114326 175130 114386 175475
rect 115798 175130 115858 177515
rect 118371 176764 118437 176765
rect 118371 176700 118372 176764
rect 118436 176700 118437 176764
rect 118371 176699 118437 176700
rect 116899 175676 116965 175677
rect 116899 175612 116900 175676
rect 116964 175612 116965 175676
rect 116899 175611 116965 175612
rect 114326 175070 114428 175130
rect 112056 174494 112116 175070
rect 113144 174494 113204 175070
rect 114368 174494 114428 175070
rect 115728 175070 115858 175130
rect 116902 175130 116962 175611
rect 118374 175130 118434 176699
rect 118794 176600 119414 191898
rect 123294 232954 123914 268398
rect 124811 255100 124877 255101
rect 124811 255036 124812 255100
rect 124876 255036 124877 255100
rect 124811 255035 124877 255036
rect 123294 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 123914 232954
rect 123294 232634 123914 232718
rect 123294 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 123914 232634
rect 123294 196954 123914 232398
rect 124814 200701 124874 255035
rect 126102 242181 126162 292979
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 126099 242180 126165 242181
rect 126099 242116 126100 242180
rect 126164 242116 126165 242180
rect 126099 242115 126165 242116
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 124811 200700 124877 200701
rect 124811 200636 124812 200700
rect 124876 200636 124877 200700
rect 124811 200635 124877 200636
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 119659 177580 119725 177581
rect 119659 177516 119660 177580
rect 119724 177516 119725 177580
rect 119659 177515 119725 177516
rect 120763 177580 120829 177581
rect 120763 177516 120764 177580
rect 120828 177516 120829 177580
rect 120763 177515 120829 177516
rect 119662 175130 119722 177515
rect 120766 175130 120826 177515
rect 121867 176764 121933 176765
rect 121867 176700 121868 176764
rect 121932 176700 121933 176764
rect 121867 176699 121933 176700
rect 122971 176764 123037 176765
rect 122971 176700 122972 176764
rect 123036 176700 123037 176764
rect 122971 176699 123037 176700
rect 121870 175130 121930 176699
rect 116902 175070 117012 175130
rect 115728 174494 115788 175070
rect 116952 174494 117012 175070
rect 118312 175070 118434 175130
rect 119400 175070 119722 175130
rect 120760 175070 120826 175130
rect 121848 175070 121930 175130
rect 122974 175130 123034 176699
rect 123294 176600 123914 196398
rect 125731 177580 125797 177581
rect 125731 177516 125732 177580
rect 125796 177516 125797 177580
rect 125731 177515 125797 177516
rect 127019 177580 127085 177581
rect 127019 177516 127020 177580
rect 127084 177516 127085 177580
rect 127019 177515 127085 177516
rect 124443 175676 124509 175677
rect 124443 175612 124444 175676
rect 124508 175612 124509 175676
rect 124443 175611 124509 175612
rect 124446 175130 124506 175611
rect 125734 175130 125794 177515
rect 127022 175130 127082 177515
rect 127794 176600 128414 200898
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 241954 132914 277398
rect 132294 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 132914 241954
rect 132294 241634 132914 241718
rect 132294 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 132914 241634
rect 132294 205954 132914 241398
rect 132294 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 132914 205954
rect 132294 205634 132914 205718
rect 132294 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 132914 205634
rect 130699 177580 130765 177581
rect 130699 177516 130700 177580
rect 130764 177516 130765 177580
rect 130699 177515 130765 177516
rect 129411 176764 129477 176765
rect 129411 176700 129412 176764
rect 129476 176700 129477 176764
rect 129411 176699 129477 176700
rect 128123 176492 128189 176493
rect 128123 176428 128124 176492
rect 128188 176428 128189 176492
rect 128123 176427 128189 176428
rect 128126 175130 128186 176427
rect 122974 175070 123132 175130
rect 118312 174494 118372 175070
rect 119400 174494 119460 175070
rect 120760 174494 120820 175070
rect 121848 174494 121908 175070
rect 123072 174494 123132 175070
rect 124432 175070 124506 175130
rect 125656 175070 125794 175130
rect 127016 175070 127082 175130
rect 128104 175070 128186 175130
rect 129414 175130 129474 176699
rect 130702 175130 130762 177515
rect 131987 177036 132053 177037
rect 131987 176972 131988 177036
rect 132052 176972 132053 177036
rect 131987 176971 132053 176972
rect 129414 175070 129524 175130
rect 124432 174494 124492 175070
rect 125656 174494 125716 175070
rect 127016 174494 127076 175070
rect 128104 174494 128164 175070
rect 129464 174494 129524 175070
rect 130688 175070 130762 175130
rect 131990 175130 132050 176971
rect 132294 176600 132914 205398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 246454 137414 281898
rect 136794 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 137414 246454
rect 136794 246134 137414 246218
rect 136794 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 137414 246134
rect 136794 210454 137414 245898
rect 136794 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 137414 210454
rect 136794 210134 137414 210218
rect 136794 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 137414 210134
rect 133091 176764 133157 176765
rect 133091 176700 133092 176764
rect 133156 176700 133157 176764
rect 133091 176699 133157 176700
rect 135667 176764 135733 176765
rect 135667 176700 135668 176764
rect 135732 176700 135733 176764
rect 135667 176699 135733 176700
rect 133094 175130 133154 176699
rect 134379 175676 134445 175677
rect 134379 175612 134380 175676
rect 134444 175612 134445 175676
rect 134379 175611 134445 175612
rect 134382 175130 134442 175611
rect 131990 175070 132108 175130
rect 133094 175070 133196 175130
rect 130688 174494 130748 175070
rect 132048 174494 132108 175070
rect 133136 174494 133196 175070
rect 134360 175070 134442 175130
rect 135670 175130 135730 176699
rect 136794 176600 137414 209898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 214954 141914 250398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 149651 299436 149717 299437
rect 149651 299372 149652 299436
rect 149716 299372 149717 299436
rect 149651 299371 149717 299372
rect 149654 298213 149714 299371
rect 149651 298212 149717 298213
rect 149651 298148 149652 298212
rect 149716 298148 149717 298212
rect 149651 298147 149717 298148
rect 146891 292908 146957 292909
rect 146891 292844 146892 292908
rect 146956 292844 146957 292908
rect 146891 292843 146957 292844
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 142659 248436 142725 248437
rect 142659 248372 142660 248436
rect 142724 248372 142725 248436
rect 142659 248371 142725 248372
rect 142662 216613 142722 248371
rect 145794 219454 146414 254898
rect 146894 235245 146954 292843
rect 149654 238781 149714 298147
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 149651 238780 149717 238781
rect 149651 238716 149652 238780
rect 149716 238716 149717 238780
rect 149651 238715 149717 238716
rect 146891 235244 146957 235245
rect 146891 235180 146892 235244
rect 146956 235180 146957 235244
rect 146891 235179 146957 235180
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 142659 216612 142725 216613
rect 142659 216548 142660 216612
rect 142724 216548 142725 216612
rect 142659 216547 142725 216548
rect 141294 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 141914 214954
rect 141294 214634 141914 214718
rect 141294 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 141914 214634
rect 141294 178954 141914 214398
rect 141294 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 141914 178954
rect 141294 178634 141914 178718
rect 141294 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 141914 178634
rect 141294 176600 141914 178398
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 176600 146414 182898
rect 150294 223954 150914 259398
rect 150294 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 150914 223954
rect 150294 223634 150914 223718
rect 150294 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 150914 223634
rect 150294 187954 150914 223398
rect 150294 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 150914 187954
rect 150294 187634 150914 187718
rect 150294 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 150914 187634
rect 148179 176764 148245 176765
rect 148179 176700 148180 176764
rect 148244 176700 148245 176764
rect 148179 176699 148245 176700
rect 148182 175130 148242 176699
rect 150294 176600 150914 187398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 167499 354924 167565 354925
rect 167499 354860 167500 354924
rect 167564 354860 167565 354924
rect 167499 354859 167565 354860
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 161243 311948 161309 311949
rect 161243 311884 161244 311948
rect 161308 311884 161309 311948
rect 161243 311883 161309 311884
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 158483 296852 158549 296853
rect 158483 296788 158484 296852
rect 158548 296788 158549 296852
rect 158483 296787 158549 296788
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 228454 155414 263898
rect 156459 257276 156525 257277
rect 156459 257212 156460 257276
rect 156524 257212 156525 257276
rect 156459 257211 156525 257212
rect 154794 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 155414 228454
rect 154794 228134 155414 228218
rect 154794 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 155414 228134
rect 154794 192454 155414 227898
rect 156462 200837 156522 257211
rect 158486 232661 158546 296787
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 232954 159914 268398
rect 161246 234565 161306 311883
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 166211 296988 166277 296989
rect 166211 296924 166212 296988
rect 166276 296924 166277 296988
rect 166211 296923 166277 296924
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 161979 266388 162045 266389
rect 161979 266324 161980 266388
rect 162044 266324 162045 266388
rect 161979 266323 162045 266324
rect 161982 239461 162042 266323
rect 161979 239460 162045 239461
rect 161979 239396 161980 239460
rect 162044 239396 162045 239460
rect 161979 239395 162045 239396
rect 161243 234564 161309 234565
rect 161243 234500 161244 234564
rect 161308 234500 161309 234564
rect 161243 234499 161309 234500
rect 159294 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 159914 232954
rect 158483 232660 158549 232661
rect 158483 232596 158484 232660
rect 158548 232596 158549 232660
rect 158483 232595 158549 232596
rect 159294 232634 159914 232718
rect 159294 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 159914 232634
rect 156459 200836 156525 200837
rect 156459 200772 156460 200836
rect 156524 200772 156525 200836
rect 156459 200771 156525 200772
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 154794 176600 155414 191898
rect 159294 196954 159914 232398
rect 161982 228853 162042 239395
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 161979 228852 162045 228853
rect 161979 228788 161980 228852
rect 162044 228788 162045 228852
rect 161979 228787 162045 228788
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 159294 196634 159914 196718
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 158851 176764 158917 176765
rect 158851 176700 158852 176764
rect 158916 176700 158917 176764
rect 158851 176699 158917 176700
rect 158854 175130 158914 176699
rect 159294 176600 159914 196398
rect 163794 201454 164414 236898
rect 166214 233205 166274 296923
rect 167502 244901 167562 354859
rect 168294 349954 168914 385398
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 171731 354788 171797 354789
rect 171731 354724 171732 354788
rect 171796 354724 171797 354788
rect 171731 354723 171797 354724
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 167683 298348 167749 298349
rect 167683 298284 167684 298348
rect 167748 298284 167749 298348
rect 167683 298283 167749 298284
rect 167499 244900 167565 244901
rect 167499 244836 167500 244900
rect 167564 244836 167565 244900
rect 167499 244835 167565 244836
rect 167686 235925 167746 298283
rect 168294 277954 168914 313398
rect 170259 294132 170325 294133
rect 170259 294068 170260 294132
rect 170324 294068 170325 294132
rect 170259 294067 170325 294068
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 241954 168914 277398
rect 169155 265164 169221 265165
rect 169155 265100 169156 265164
rect 169220 265100 169221 265164
rect 169155 265099 169221 265100
rect 168294 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 168914 241954
rect 168294 241634 168914 241718
rect 168294 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 168914 241634
rect 167683 235924 167749 235925
rect 167683 235860 167684 235924
rect 167748 235860 167749 235924
rect 167683 235859 167749 235860
rect 166211 233204 166277 233205
rect 166211 233140 166212 233204
rect 166276 233140 166277 233204
rect 166211 233139 166277 233140
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 176600 164414 200898
rect 168294 205954 168914 241398
rect 168294 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 168914 205954
rect 168294 205634 168914 205718
rect 168294 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 168914 205634
rect 167499 181660 167565 181661
rect 167499 181596 167500 181660
rect 167564 181596 167565 181660
rect 167499 181595 167565 181596
rect 166395 178124 166461 178125
rect 166395 178060 166396 178124
rect 166460 178060 166461 178124
rect 166395 178059 166461 178060
rect 166211 175540 166277 175541
rect 166211 175476 166212 175540
rect 166276 175476 166277 175540
rect 166211 175475 166277 175476
rect 135670 175070 135780 175130
rect 148182 175070 148292 175130
rect 134360 174494 134420 175070
rect 135720 174494 135780 175070
rect 148232 174494 148292 175070
rect 158840 175070 158914 175130
rect 158840 174494 158900 175070
rect 166214 164389 166274 175475
rect 166211 164388 166277 164389
rect 166211 164324 166212 164388
rect 166276 164324 166277 164388
rect 166211 164323 166277 164324
rect 166398 154597 166458 178059
rect 166395 154596 166461 154597
rect 166395 154532 166396 154596
rect 166460 154532 166461 154596
rect 166395 154531 166461 154532
rect 69072 151954 69420 151986
rect 69072 151718 69128 151954
rect 69364 151718 69420 151954
rect 69072 151634 69420 151718
rect 69072 151398 69128 151634
rect 69364 151398 69420 151634
rect 69072 151366 69420 151398
rect 164136 151954 164484 151986
rect 164136 151718 164192 151954
rect 164428 151718 164484 151954
rect 164136 151634 164484 151718
rect 164136 151398 164192 151634
rect 164428 151398 164484 151634
rect 164136 151366 164484 151398
rect 69752 147454 70100 147486
rect 69752 147218 69808 147454
rect 70044 147218 70100 147454
rect 69752 147134 70100 147218
rect 69752 146898 69808 147134
rect 70044 146898 70100 147134
rect 69752 146866 70100 146898
rect 163456 147454 163804 147486
rect 163456 147218 163512 147454
rect 163748 147218 163804 147454
rect 163456 147134 163804 147218
rect 163456 146898 163512 147134
rect 163748 146898 163804 147134
rect 163456 146866 163804 146898
rect 166395 133924 166461 133925
rect 166395 133860 166396 133924
rect 166460 133860 166461 133924
rect 166395 133859 166461 133860
rect 166211 131476 166277 131477
rect 166211 131412 166212 131476
rect 166276 131412 166277 131476
rect 166211 131411 166277 131412
rect 69072 115954 69420 115986
rect 69072 115718 69128 115954
rect 69364 115718 69420 115954
rect 69072 115634 69420 115718
rect 69072 115398 69128 115634
rect 69364 115398 69420 115634
rect 69072 115366 69420 115398
rect 164136 115954 164484 115986
rect 164136 115718 164192 115954
rect 164428 115718 164484 115954
rect 164136 115634 164484 115718
rect 164136 115398 164192 115634
rect 164428 115398 164484 115634
rect 164136 115366 164484 115398
rect 69752 111454 70100 111486
rect 69752 111218 69808 111454
rect 70044 111218 70100 111454
rect 69752 111134 70100 111218
rect 69752 110898 69808 111134
rect 70044 110898 70100 111134
rect 69752 110866 70100 110898
rect 163456 111454 163804 111486
rect 163456 111218 163512 111454
rect 163748 111218 163804 111454
rect 163456 111134 163804 111218
rect 163456 110898 163512 111134
rect 163748 110898 163804 111134
rect 163456 110866 163804 110898
rect 74656 94890 74716 95200
rect 84312 94890 84372 95200
rect 85536 94890 85596 95200
rect 86624 94890 86684 95200
rect 87984 94890 88044 95200
rect 88936 94890 88996 95200
rect 74656 94830 74826 94890
rect 84312 94830 84394 94890
rect 85536 94830 85682 94890
rect 86624 94830 86786 94890
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 70954 69914 93100
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 75454 74414 93100
rect 74766 91221 74826 94830
rect 74763 91220 74829 91221
rect 74763 91156 74764 91220
rect 74828 91156 74829 91220
rect 74763 91155 74829 91156
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 79954 78914 93100
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 84454 83414 93100
rect 84334 91221 84394 94830
rect 85622 92445 85682 94830
rect 85619 92444 85685 92445
rect 85619 92380 85620 92444
rect 85684 92380 85685 92444
rect 85619 92379 85685 92380
rect 86726 91221 86786 94830
rect 87094 94830 88044 94890
rect 88934 94830 88996 94890
rect 90160 94890 90220 95200
rect 91384 94890 91444 95200
rect 90160 94830 90282 94890
rect 87094 92445 87154 94830
rect 87091 92444 87157 92445
rect 87091 92380 87092 92444
rect 87156 92380 87157 92444
rect 87091 92379 87157 92380
rect 84331 91220 84397 91221
rect 84331 91156 84332 91220
rect 84396 91156 84397 91220
rect 84331 91155 84397 91156
rect 86723 91220 86789 91221
rect 86723 91156 86724 91220
rect 86788 91156 86789 91220
rect 86723 91155 86789 91156
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 88954 87914 93100
rect 88934 92445 88994 94830
rect 88931 92444 88997 92445
rect 88931 92380 88932 92444
rect 88996 92380 88997 92444
rect 88931 92379 88997 92380
rect 90222 91221 90282 94830
rect 91326 94830 91444 94890
rect 92472 94890 92532 95200
rect 93832 94890 93892 95200
rect 94920 94890 94980 95200
rect 96008 94890 96068 95200
rect 96688 94890 96748 95200
rect 97096 94890 97156 95200
rect 98048 94890 98108 95200
rect 98456 94890 98516 95200
rect 99136 94890 99196 95200
rect 99544 94890 99604 95200
rect 100632 94890 100692 95200
rect 92472 94830 92674 94890
rect 93832 94830 93962 94890
rect 94920 94830 95066 94890
rect 96008 94830 96170 94890
rect 96688 94830 96906 94890
rect 97096 94830 97274 94890
rect 98048 94830 98194 94890
rect 98456 94830 98562 94890
rect 99136 94830 99298 94890
rect 99544 94830 99666 94890
rect 91326 91221 91386 94830
rect 90219 91220 90285 91221
rect 90219 91156 90220 91220
rect 90284 91156 90285 91220
rect 90219 91155 90285 91156
rect 91323 91220 91389 91221
rect 91323 91156 91324 91220
rect 91388 91156 91389 91220
rect 91323 91155 91389 91156
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 57454 92414 93100
rect 92614 91221 92674 94830
rect 93902 93533 93962 94830
rect 93899 93532 93965 93533
rect 93899 93468 93900 93532
rect 93964 93468 93965 93532
rect 93899 93467 93965 93468
rect 95006 91221 95066 94830
rect 96110 91221 96170 94830
rect 96846 93870 96906 94830
rect 96846 93810 97090 93870
rect 92611 91220 92677 91221
rect 92611 91156 92612 91220
rect 92676 91156 92677 91220
rect 92611 91155 92677 91156
rect 95003 91220 95069 91221
rect 95003 91156 95004 91220
rect 95068 91156 95069 91220
rect 95003 91155 95069 91156
rect 96107 91220 96173 91221
rect 96107 91156 96108 91220
rect 96172 91156 96173 91220
rect 96107 91155 96173 91156
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 61954 96914 93100
rect 97030 91221 97090 93810
rect 97214 91221 97274 94830
rect 98134 91357 98194 94830
rect 98502 91493 98562 94830
rect 98499 91492 98565 91493
rect 98499 91428 98500 91492
rect 98564 91428 98565 91492
rect 98499 91427 98565 91428
rect 98131 91356 98197 91357
rect 98131 91292 98132 91356
rect 98196 91292 98197 91356
rect 98131 91291 98197 91292
rect 99238 91221 99298 94830
rect 99606 92445 99666 94830
rect 100526 94830 100692 94890
rect 100768 94890 100828 95200
rect 101856 94890 101916 95200
rect 100768 94830 101690 94890
rect 99603 92444 99669 92445
rect 99603 92380 99604 92444
rect 99668 92380 99669 92444
rect 99603 92379 99669 92380
rect 100526 91221 100586 94830
rect 97027 91220 97093 91221
rect 97027 91156 97028 91220
rect 97092 91156 97093 91220
rect 97027 91155 97093 91156
rect 97211 91220 97277 91221
rect 97211 91156 97212 91220
rect 97276 91156 97277 91220
rect 97211 91155 97277 91156
rect 99235 91220 99301 91221
rect 99235 91156 99236 91220
rect 99300 91156 99301 91220
rect 99235 91155 99301 91156
rect 100523 91220 100589 91221
rect 100523 91156 100524 91220
rect 100588 91156 100589 91220
rect 100523 91155 100589 91156
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 66454 101414 93100
rect 101630 91357 101690 94830
rect 101814 94830 101916 94890
rect 101992 94890 102052 95200
rect 102944 94890 103004 95200
rect 101992 94830 102058 94890
rect 101814 91493 101874 94830
rect 101811 91492 101877 91493
rect 101811 91428 101812 91492
rect 101876 91428 101877 91492
rect 101811 91427 101877 91428
rect 101627 91356 101693 91357
rect 101627 91292 101628 91356
rect 101692 91292 101693 91356
rect 101627 91291 101693 91292
rect 101998 91221 102058 94830
rect 102918 94830 103004 94890
rect 103216 94890 103276 95200
rect 103216 94830 103346 94890
rect 102918 91357 102978 94830
rect 102915 91356 102981 91357
rect 102915 91292 102916 91356
rect 102980 91292 102981 91356
rect 102915 91291 102981 91292
rect 103286 91221 103346 94830
rect 104304 94754 104364 95200
rect 104206 94694 104364 94754
rect 104440 94754 104500 95200
rect 105392 94754 105452 95200
rect 104440 94694 104634 94754
rect 104206 91629 104266 94694
rect 104203 91628 104269 91629
rect 104203 91564 104204 91628
rect 104268 91564 104269 91628
rect 104203 91563 104269 91564
rect 104574 91221 104634 94694
rect 105126 94694 105452 94754
rect 105664 94754 105724 95200
rect 106480 94754 106540 95200
rect 105664 94694 106106 94754
rect 105126 91357 105186 94694
rect 105123 91356 105189 91357
rect 105123 91292 105124 91356
rect 105188 91292 105189 91356
rect 105123 91291 105189 91292
rect 101995 91220 102061 91221
rect 101995 91156 101996 91220
rect 102060 91156 102061 91220
rect 101995 91155 102061 91156
rect 103283 91220 103349 91221
rect 103283 91156 103284 91220
rect 103348 91156 103349 91220
rect 103283 91155 103349 91156
rect 104571 91220 104637 91221
rect 104571 91156 104572 91220
rect 104636 91156 104637 91220
rect 104571 91155 104637 91156
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 70954 105914 93100
rect 106046 91221 106106 94694
rect 106414 94694 106540 94754
rect 106616 94754 106676 95200
rect 107704 94754 107764 95200
rect 108112 94754 108172 95200
rect 106616 94694 106842 94754
rect 106414 91221 106474 94694
rect 106782 92445 106842 94694
rect 107702 94694 107764 94754
rect 108070 94694 108172 94754
rect 109064 94754 109124 95200
rect 109472 94754 109532 95200
rect 110152 94754 110212 95200
rect 110696 94754 110756 95200
rect 111240 94754 111300 95200
rect 109064 94694 109234 94754
rect 109472 94694 109602 94754
rect 107702 93533 107762 94694
rect 107699 93532 107765 93533
rect 107699 93468 107700 93532
rect 107764 93468 107765 93532
rect 107699 93467 107765 93468
rect 106779 92444 106845 92445
rect 106779 92380 106780 92444
rect 106844 92380 106845 92444
rect 106779 92379 106845 92380
rect 108070 91221 108130 94694
rect 109174 92445 109234 94694
rect 109171 92444 109237 92445
rect 109171 92380 109172 92444
rect 109236 92380 109237 92444
rect 109171 92379 109237 92380
rect 109542 91221 109602 94694
rect 110094 94694 110212 94754
rect 110646 94694 110756 94754
rect 111198 94694 111300 94754
rect 111920 94754 111980 95200
rect 112328 94757 112388 95200
rect 113144 94757 113204 95200
rect 112325 94756 112391 94757
rect 111920 94694 111994 94754
rect 110094 93261 110154 94694
rect 110091 93260 110157 93261
rect 110091 93196 110092 93260
rect 110156 93196 110157 93260
rect 110091 93195 110157 93196
rect 106043 91220 106109 91221
rect 106043 91156 106044 91220
rect 106108 91156 106109 91220
rect 106043 91155 106109 91156
rect 106411 91220 106477 91221
rect 106411 91156 106412 91220
rect 106476 91156 106477 91220
rect 106411 91155 106477 91156
rect 108067 91220 108133 91221
rect 108067 91156 108068 91220
rect 108132 91156 108133 91220
rect 108067 91155 108133 91156
rect 109539 91220 109605 91221
rect 109539 91156 109540 91220
rect 109604 91156 109605 91220
rect 109539 91155 109605 91156
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 75454 110414 93100
rect 110646 91221 110706 94694
rect 111198 92445 111258 94694
rect 111195 92444 111261 92445
rect 111195 92380 111196 92444
rect 111260 92380 111261 92444
rect 111195 92379 111261 92380
rect 111934 91221 111994 94694
rect 112325 94692 112326 94756
rect 112390 94692 112391 94756
rect 112325 94691 112391 94692
rect 113141 94756 113207 94757
rect 113141 94692 113142 94756
rect 113206 94692 113207 94756
rect 113688 94754 113748 95200
rect 114368 94754 114428 95200
rect 113688 94694 113834 94754
rect 113141 94691 113207 94692
rect 113774 91221 113834 94694
rect 114142 94694 114428 94754
rect 114776 94754 114836 95200
rect 115456 94754 115516 95200
rect 115864 94754 115924 95200
rect 114776 94694 115122 94754
rect 114142 92445 114202 94694
rect 114139 92444 114205 92445
rect 114139 92380 114140 92444
rect 114204 92380 114205 92444
rect 114139 92379 114205 92380
rect 110643 91220 110709 91221
rect 110643 91156 110644 91220
rect 110708 91156 110709 91220
rect 110643 91155 110709 91156
rect 111931 91220 111997 91221
rect 111931 91156 111932 91220
rect 111996 91156 111997 91220
rect 111931 91155 111997 91156
rect 113771 91220 113837 91221
rect 113771 91156 113772 91220
rect 113836 91156 113837 91220
rect 113771 91155 113837 91156
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 79954 114914 93100
rect 115062 91765 115122 94694
rect 115430 94694 115516 94754
rect 115798 94694 115924 94754
rect 116680 94754 116740 95200
rect 117088 94754 117148 95200
rect 116680 94694 116778 94754
rect 115430 92309 115490 94694
rect 115427 92308 115493 92309
rect 115427 92244 115428 92308
rect 115492 92244 115493 92308
rect 115427 92243 115493 92244
rect 115059 91764 115125 91765
rect 115059 91700 115060 91764
rect 115124 91700 115125 91764
rect 115059 91699 115125 91700
rect 115798 91221 115858 94694
rect 116718 93805 116778 94694
rect 117086 94694 117148 94754
rect 117904 94754 117964 95200
rect 118176 94754 118236 95200
rect 119400 94757 119460 95200
rect 119397 94756 119463 94757
rect 117904 94694 118066 94754
rect 118176 94694 118250 94754
rect 116715 93804 116781 93805
rect 116715 93740 116716 93804
rect 116780 93740 116781 93804
rect 116715 93739 116781 93740
rect 117086 91221 117146 94694
rect 118006 92445 118066 94694
rect 118003 92444 118069 92445
rect 118003 92380 118004 92444
rect 118068 92380 118069 92444
rect 118003 92379 118069 92380
rect 118190 91221 118250 94694
rect 119397 94692 119398 94756
rect 119462 94692 119463 94756
rect 119536 94754 119596 95200
rect 119843 94756 119909 94757
rect 119536 94694 119722 94754
rect 119397 94691 119463 94692
rect 115795 91220 115861 91221
rect 115795 91156 115796 91220
rect 115860 91156 115861 91220
rect 115795 91155 115861 91156
rect 117083 91220 117149 91221
rect 117083 91156 117084 91220
rect 117148 91156 117149 91220
rect 117083 91155 117149 91156
rect 118187 91220 118253 91221
rect 118187 91156 118188 91220
rect 118252 91156 118253 91220
rect 118187 91155 118253 91156
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114294 43954 114914 79398
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 84454 119414 93100
rect 119662 91221 119722 94694
rect 119843 94692 119844 94756
rect 119908 94692 119909 94756
rect 120216 94754 120276 95200
rect 120624 94754 120684 95200
rect 121712 94754 121772 95200
rect 119843 94691 119909 94692
rect 120214 94694 120276 94754
rect 120582 94694 120684 94754
rect 121686 94694 121772 94754
rect 121984 94754 122044 95200
rect 122800 94890 122860 95200
rect 122800 94830 123034 94890
rect 121984 94694 122114 94754
rect 119846 91357 119906 94691
rect 119843 91356 119909 91357
rect 119843 91292 119844 91356
rect 119908 91292 119909 91356
rect 119843 91291 119909 91292
rect 120214 91221 120274 94694
rect 120582 91357 120642 94694
rect 121686 93669 121746 94694
rect 121683 93668 121749 93669
rect 121683 93604 121684 93668
rect 121748 93604 121749 93668
rect 121683 93603 121749 93604
rect 120579 91356 120645 91357
rect 120579 91292 120580 91356
rect 120644 91292 120645 91356
rect 120579 91291 120645 91292
rect 122054 91221 122114 94694
rect 122974 93870 123034 94830
rect 123208 94757 123268 95200
rect 124024 94890 124084 95200
rect 124432 94890 124492 95200
rect 125384 94890 125444 95200
rect 124024 94830 124138 94890
rect 124432 94830 124506 94890
rect 123205 94756 123271 94757
rect 123205 94692 123206 94756
rect 123270 94692 123271 94756
rect 123205 94691 123271 94692
rect 122606 93810 123034 93870
rect 122606 91490 122666 93810
rect 122787 91492 122853 91493
rect 122787 91490 122788 91492
rect 122606 91430 122788 91490
rect 122787 91428 122788 91430
rect 122852 91428 122853 91492
rect 122787 91427 122853 91428
rect 119659 91220 119725 91221
rect 119659 91156 119660 91220
rect 119724 91156 119725 91220
rect 119659 91155 119725 91156
rect 120211 91220 120277 91221
rect 120211 91156 120212 91220
rect 120276 91156 120277 91220
rect 120211 91155 120277 91156
rect 122051 91220 122117 91221
rect 122051 91156 122052 91220
rect 122116 91156 122117 91220
rect 122051 91155 122117 91156
rect 118794 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 119414 84454
rect 118794 84134 119414 84218
rect 118794 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 119414 84134
rect 118794 48454 119414 83898
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 88954 123914 93100
rect 124078 91221 124138 94830
rect 124446 92445 124506 94830
rect 125366 94830 125444 94890
rect 125656 94890 125716 95200
rect 126472 94890 126532 95200
rect 125656 94830 125794 94890
rect 125366 92445 125426 94830
rect 125734 92445 125794 94830
rect 126470 94830 126532 94890
rect 126608 94890 126668 95200
rect 128104 94890 128164 95200
rect 129328 94890 129388 95200
rect 130688 94890 130748 95200
rect 131912 94890 131972 95200
rect 133136 94890 133196 95200
rect 126608 94830 126714 94890
rect 128104 94830 128186 94890
rect 129328 94830 129474 94890
rect 130688 94830 130762 94890
rect 131912 94830 132050 94890
rect 124443 92444 124509 92445
rect 124443 92380 124444 92444
rect 124508 92380 124509 92444
rect 124443 92379 124509 92380
rect 125363 92444 125429 92445
rect 125363 92380 125364 92444
rect 125428 92380 125429 92444
rect 125363 92379 125429 92380
rect 125731 92444 125797 92445
rect 125731 92380 125732 92444
rect 125796 92380 125797 92444
rect 125731 92379 125797 92380
rect 126470 91221 126530 94830
rect 126654 91357 126714 94830
rect 128126 93261 128186 94830
rect 128123 93260 128189 93261
rect 128123 93196 128124 93260
rect 128188 93196 128189 93260
rect 128123 93195 128189 93196
rect 126651 91356 126717 91357
rect 126651 91292 126652 91356
rect 126716 91292 126717 91356
rect 126651 91291 126717 91292
rect 124075 91220 124141 91221
rect 124075 91156 124076 91220
rect 124140 91156 124141 91220
rect 124075 91155 124141 91156
rect 126467 91220 126533 91221
rect 126467 91156 126468 91220
rect 126532 91156 126533 91220
rect 126467 91155 126533 91156
rect 123294 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 123914 88954
rect 123294 88634 123914 88718
rect 123294 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 123914 88634
rect 123294 52954 123914 88398
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 57454 128414 93100
rect 129414 92445 129474 94830
rect 129411 92444 129477 92445
rect 129411 92380 129412 92444
rect 129476 92380 129477 92444
rect 129411 92379 129477 92380
rect 130702 91221 130762 94830
rect 131990 91629 132050 94830
rect 133094 94830 133196 94890
rect 134360 94890 134420 95200
rect 135584 94890 135644 95200
rect 134360 94830 134442 94890
rect 135584 94830 135730 94890
rect 131987 91628 132053 91629
rect 131987 91564 131988 91628
rect 132052 91564 132053 91628
rect 131987 91563 132053 91564
rect 130699 91220 130765 91221
rect 130699 91156 130700 91220
rect 130764 91156 130765 91220
rect 130699 91155 130765 91156
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 61954 132914 93100
rect 133094 91221 133154 94830
rect 134382 91221 134442 94830
rect 135670 92445 135730 94830
rect 151307 94756 151373 94757
rect 151307 94692 151308 94756
rect 151372 94692 151373 94756
rect 151496 94754 151556 95200
rect 151632 94757 151692 95200
rect 151307 94691 151373 94692
rect 151494 94694 151556 94754
rect 151629 94756 151695 94757
rect 135667 92444 135733 92445
rect 135667 92380 135668 92444
rect 135732 92380 135733 92444
rect 135667 92379 135733 92380
rect 133091 91220 133157 91221
rect 133091 91156 133092 91220
rect 133156 91156 133157 91220
rect 133091 91155 133157 91156
rect 134379 91220 134445 91221
rect 134379 91156 134380 91220
rect 134444 91156 134445 91220
rect 134379 91155 134445 91156
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5146 132914 25398
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 66454 137414 93100
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6106 137414 29898
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 70954 141914 93100
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7066 141914 34398
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 75454 146414 93100
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 79954 150914 93100
rect 151310 91629 151370 94691
rect 151494 93533 151554 94694
rect 151629 94692 151630 94756
rect 151694 94692 151695 94756
rect 151629 94691 151695 94692
rect 151768 94210 151828 95200
rect 151904 94757 151964 95200
rect 151901 94756 151967 94757
rect 151901 94692 151902 94756
rect 151966 94692 151967 94756
rect 151901 94691 151967 94692
rect 151678 94150 151828 94210
rect 151491 93532 151557 93533
rect 151491 93468 151492 93532
rect 151556 93468 151557 93532
rect 151491 93467 151557 93468
rect 151678 92173 151738 94150
rect 151675 92172 151741 92173
rect 151675 92108 151676 92172
rect 151740 92108 151741 92172
rect 151675 92107 151741 92108
rect 151307 91628 151373 91629
rect 151307 91564 151308 91628
rect 151372 91564 151373 91628
rect 151307 91563 151373 91564
rect 150294 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 150914 79954
rect 150294 79634 150914 79718
rect 150294 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 150914 79634
rect 150294 43954 150914 79398
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 84454 155414 93100
rect 154794 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 155414 84454
rect 154794 84134 155414 84218
rect 154794 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 155414 84134
rect 154794 48454 155414 83898
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 88954 159914 93100
rect 159294 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 159914 88954
rect 159294 88634 159914 88718
rect 159294 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 159914 88634
rect 159294 52954 159914 88398
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 57454 164414 93100
rect 166214 84149 166274 131411
rect 166398 88229 166458 133859
rect 167315 97204 167381 97205
rect 167315 97140 167316 97204
rect 167380 97140 167381 97204
rect 167315 97139 167381 97140
rect 167318 92309 167378 97139
rect 167502 94485 167562 181595
rect 167683 175404 167749 175405
rect 167683 175340 167684 175404
rect 167748 175340 167749 175404
rect 167683 175339 167749 175340
rect 167686 158813 167746 175339
rect 168294 169954 168914 205398
rect 168294 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 168914 169954
rect 168294 169634 168914 169718
rect 168294 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 168914 169634
rect 167683 158812 167749 158813
rect 167683 158748 167684 158812
rect 167748 158748 167749 158812
rect 167683 158747 167749 158748
rect 168294 133954 168914 169398
rect 168294 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 168914 133954
rect 168294 133634 168914 133718
rect 168294 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 168914 133634
rect 167683 127260 167749 127261
rect 167683 127196 167684 127260
rect 167748 127196 167749 127260
rect 167683 127195 167749 127196
rect 167499 94484 167565 94485
rect 167499 94420 167500 94484
rect 167564 94420 167565 94484
rect 167499 94419 167565 94420
rect 167315 92308 167381 92309
rect 167315 92244 167316 92308
rect 167380 92244 167381 92308
rect 167315 92243 167381 92244
rect 166395 88228 166461 88229
rect 166395 88164 166396 88228
rect 166460 88164 166461 88228
rect 166395 88163 166461 88164
rect 167686 86869 167746 127195
rect 168294 97954 168914 133398
rect 168294 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 168914 97954
rect 168294 97634 168914 97718
rect 168294 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 168914 97634
rect 167683 86868 167749 86869
rect 167683 86804 167684 86868
rect 167748 86804 167749 86868
rect 167683 86803 167749 86804
rect 166211 84148 166277 84149
rect 166211 84084 166212 84148
rect 166276 84084 166277 84148
rect 166211 84083 166277 84084
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 61954 168914 97398
rect 169158 93805 169218 265099
rect 170262 171733 170322 294067
rect 171734 247077 171794 354723
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177067 350164 177133 350165
rect 177067 350100 177068 350164
rect 177132 350100 177133 350164
rect 177067 350099 177133 350100
rect 173755 339284 173821 339285
rect 173755 339220 173756 339284
rect 173820 339220 173821 339284
rect 173755 339219 173821 339220
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 171915 267884 171981 267885
rect 171915 267820 171916 267884
rect 171980 267820 171981 267884
rect 171915 267819 171981 267820
rect 171731 247076 171797 247077
rect 171731 247012 171732 247076
rect 171796 247012 171797 247076
rect 171731 247011 171797 247012
rect 171918 211853 171978 267819
rect 172794 246454 173414 281898
rect 172794 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 173414 246454
rect 172794 246134 173414 246218
rect 172794 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 173414 246134
rect 171915 211852 171981 211853
rect 171915 211788 171916 211852
rect 171980 211788 171981 211852
rect 171915 211787 171981 211788
rect 172794 210454 173414 245898
rect 172794 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 173414 210454
rect 172794 210134 173414 210218
rect 172794 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 173414 210134
rect 171179 183020 171245 183021
rect 171179 182956 171180 183020
rect 171244 182956 171245 183020
rect 171179 182955 171245 182956
rect 170259 171732 170325 171733
rect 170259 171668 170260 171732
rect 170324 171668 170325 171732
rect 170259 171667 170325 171668
rect 171182 160173 171242 182955
rect 172794 174454 173414 209898
rect 172794 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 173414 174454
rect 172794 174134 173414 174218
rect 172794 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 173414 174134
rect 171179 160172 171245 160173
rect 171179 160108 171180 160172
rect 171244 160108 171245 160172
rect 171179 160107 171245 160108
rect 172794 138454 173414 173898
rect 172794 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 173414 138454
rect 172794 138134 173414 138218
rect 172794 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 173414 138134
rect 171915 136916 171981 136917
rect 171915 136852 171916 136916
rect 171980 136852 171981 136916
rect 171915 136851 171981 136852
rect 170259 130116 170325 130117
rect 170259 130052 170260 130116
rect 170324 130052 170325 130116
rect 170259 130051 170325 130052
rect 169155 93804 169221 93805
rect 169155 93740 169156 93804
rect 169220 93740 169221 93804
rect 169155 93739 169221 93740
rect 170262 81429 170322 130051
rect 171731 129980 171797 129981
rect 171731 129916 171732 129980
rect 171796 129916 171797 129980
rect 171731 129915 171797 129916
rect 171734 82789 171794 129915
rect 171918 93669 171978 136851
rect 172794 102454 173414 137898
rect 172794 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 173414 102454
rect 172794 102134 173414 102218
rect 172794 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 173414 102134
rect 171915 93668 171981 93669
rect 171915 93604 171916 93668
rect 171980 93604 171981 93668
rect 171915 93603 171981 93604
rect 171731 82788 171797 82789
rect 171731 82724 171732 82788
rect 171796 82724 171797 82788
rect 171731 82723 171797 82724
rect 170259 81428 170325 81429
rect 170259 81364 170260 81428
rect 170324 81364 170325 81428
rect 170259 81363 170325 81364
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5146 168914 25398
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 66454 173414 101898
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6106 173414 29898
rect 173758 15877 173818 339219
rect 175043 330444 175109 330445
rect 175043 330380 175044 330444
rect 175108 330380 175109 330444
rect 175043 330379 175109 330380
rect 175046 42125 175106 330379
rect 176331 323644 176397 323645
rect 176331 323580 176332 323644
rect 176396 323580 176397 323644
rect 176331 323579 176397 323580
rect 176334 50285 176394 323579
rect 176515 316844 176581 316845
rect 176515 316780 176516 316844
rect 176580 316780 176581 316844
rect 176515 316779 176581 316780
rect 176331 50284 176397 50285
rect 176331 50220 176332 50284
rect 176396 50220 176397 50284
rect 176331 50219 176397 50220
rect 175043 42124 175109 42125
rect 175043 42060 175044 42124
rect 175108 42060 175109 42124
rect 175043 42059 175109 42060
rect 173755 15876 173821 15877
rect 173755 15812 173756 15876
rect 173820 15812 173821 15876
rect 173755 15811 173821 15812
rect 176518 6221 176578 316779
rect 177070 51781 177130 350099
rect 177294 322954 177914 358398
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 357154 182414 362898
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 357154 186914 367398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 357154 191414 371898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 357154 195914 376398
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 357154 200414 380898
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 357154 204914 385398
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 357154 209414 389898
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 357154 213914 358398
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 357154 218414 362898
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 547954 222914 583398
rect 222294 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 222914 547954
rect 222294 547634 222914 547718
rect 222294 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 222914 547634
rect 222294 511954 222914 547398
rect 222294 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 222914 511954
rect 222294 511634 222914 511718
rect 222294 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 222914 511634
rect 222294 475954 222914 511398
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 357154 222914 367398
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 552454 227414 587898
rect 226794 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 227414 552454
rect 226794 552134 227414 552218
rect 226794 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 227414 552134
rect 226794 516454 227414 551898
rect 226794 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 227414 516454
rect 226794 516134 227414 516218
rect 226794 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 227414 516134
rect 226794 480454 227414 515898
rect 226794 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 227414 480454
rect 226794 480134 227414 480218
rect 226794 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 227414 480134
rect 226794 444454 227414 479898
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 357154 227414 371898
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 556954 231914 592398
rect 231294 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 231914 556954
rect 231294 556634 231914 556718
rect 231294 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 231914 556634
rect 231294 520954 231914 556398
rect 231294 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 231914 520954
rect 231294 520634 231914 520718
rect 231294 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 231914 520634
rect 231294 484954 231914 520398
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 231294 412954 231914 448398
rect 231294 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 231914 412954
rect 231294 412634 231914 412718
rect 231294 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 231914 412634
rect 231294 376954 231914 412398
rect 231294 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 231914 376954
rect 231294 376634 231914 376718
rect 231294 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 231914 376634
rect 231294 357154 231914 376398
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 357154 236414 380898
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 529954 240914 565398
rect 240294 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 240914 529954
rect 240294 529634 240914 529718
rect 240294 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 240914 529634
rect 240294 493954 240914 529398
rect 240294 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 240914 493954
rect 240294 493634 240914 493718
rect 240294 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 240914 493634
rect 240294 457954 240914 493398
rect 240294 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 240914 457954
rect 240294 457634 240914 457718
rect 240294 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 240914 457634
rect 240294 421954 240914 457398
rect 240294 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 240914 421954
rect 240294 421634 240914 421718
rect 240294 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 240914 421634
rect 240294 385954 240914 421398
rect 240294 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 240914 385954
rect 240294 385634 240914 385718
rect 240294 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 240914 385634
rect 240294 357154 240914 385398
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 534454 245414 569898
rect 244794 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 245414 534454
rect 244794 534134 245414 534218
rect 244794 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 245414 534134
rect 244794 498454 245414 533898
rect 244794 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 245414 498454
rect 244794 498134 245414 498218
rect 244794 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 245414 498134
rect 244794 462454 245414 497898
rect 244794 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 245414 462454
rect 244794 462134 245414 462218
rect 244794 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 245414 462134
rect 244794 426454 245414 461898
rect 244794 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 245414 426454
rect 244794 426134 245414 426218
rect 244794 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 245414 426134
rect 244794 390454 245414 425898
rect 244794 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 245414 390454
rect 244794 390134 245414 390218
rect 244794 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 245414 390134
rect 244794 357154 245414 389898
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 538954 249914 574398
rect 249294 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 249914 538954
rect 249294 538634 249914 538718
rect 249294 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 249914 538634
rect 249294 502954 249914 538398
rect 249294 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 249914 502954
rect 249294 502634 249914 502718
rect 249294 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 249914 502634
rect 249294 466954 249914 502398
rect 249294 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 249914 466954
rect 249294 466634 249914 466718
rect 249294 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 249914 466634
rect 249294 430954 249914 466398
rect 249294 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 249914 430954
rect 249294 430634 249914 430718
rect 249294 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 249914 430634
rect 249294 394954 249914 430398
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 249294 358954 249914 394398
rect 249294 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 249914 358954
rect 249294 358634 249914 358718
rect 249294 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 249914 358634
rect 249294 357154 249914 358398
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 357154 254414 362898
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 258294 367954 258914 403398
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 258294 357154 258914 367398
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 372454 263414 407898
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 357154 263414 371898
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 376954 267914 412398
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 357154 267914 376398
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 357154 272414 380898
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 529954 276914 565398
rect 276294 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 276914 529954
rect 276294 529634 276914 529718
rect 276294 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 276914 529634
rect 276294 493954 276914 529398
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 357154 276914 385398
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 534454 281414 569898
rect 280794 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 281414 534454
rect 280794 534134 281414 534218
rect 280794 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 281414 534134
rect 280794 498454 281414 533898
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 462454 281414 497898
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 357154 281414 389898
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 357154 285914 358398
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 357154 290414 362898
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 295931 702540 295997 702541
rect 295931 702476 295932 702540
rect 295996 702476 295997 702540
rect 295931 702475 295997 702476
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294091 358868 294157 358869
rect 294091 358804 294092 358868
rect 294156 358804 294157 358868
rect 294091 358803 294157 358804
rect 292435 356284 292501 356285
rect 292435 356220 292436 356284
rect 292500 356220 292501 356284
rect 292435 356219 292501 356220
rect 292438 353290 292498 356219
rect 293171 354924 293237 354925
rect 293171 354860 293172 354924
rect 293236 354860 293237 354924
rect 293171 354859 293237 354860
rect 292438 353230 292682 353290
rect 292622 353021 292682 353230
rect 292619 353020 292685 353021
rect 292619 352956 292620 353020
rect 292684 352956 292685 353020
rect 292619 352955 292685 352956
rect 179275 334524 179341 334525
rect 179275 334460 179276 334524
rect 179340 334460 179341 334524
rect 179275 334459 179341 334460
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 250954 177914 286398
rect 178539 283252 178605 283253
rect 178539 283188 178540 283252
rect 178604 283188 178605 283252
rect 178539 283187 178605 283188
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 214954 177914 250398
rect 178542 239461 178602 283187
rect 178539 239460 178605 239461
rect 178539 239396 178540 239460
rect 178604 239396 178605 239460
rect 178539 239395 178605 239396
rect 177294 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 177914 214954
rect 177294 214634 177914 214718
rect 177294 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 177914 214634
rect 177294 178954 177914 214398
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 106954 177914 142398
rect 177294 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 177914 106954
rect 177294 106634 177914 106718
rect 177294 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 177914 106634
rect 177294 70954 177914 106398
rect 179278 91085 179338 334459
rect 199568 331954 199888 331986
rect 199568 331718 199610 331954
rect 199846 331718 199888 331954
rect 199568 331634 199888 331718
rect 199568 331398 199610 331634
rect 199846 331398 199888 331634
rect 199568 331366 199888 331398
rect 230288 331954 230608 331986
rect 230288 331718 230330 331954
rect 230566 331718 230608 331954
rect 230288 331634 230608 331718
rect 230288 331398 230330 331634
rect 230566 331398 230608 331634
rect 230288 331366 230608 331398
rect 261008 331954 261328 331986
rect 261008 331718 261050 331954
rect 261286 331718 261328 331954
rect 261008 331634 261328 331718
rect 261008 331398 261050 331634
rect 261286 331398 261328 331634
rect 261008 331366 261328 331398
rect 184208 327454 184528 327486
rect 184208 327218 184250 327454
rect 184486 327218 184528 327454
rect 184208 327134 184528 327218
rect 184208 326898 184250 327134
rect 184486 326898 184528 327134
rect 184208 326866 184528 326898
rect 214928 327454 215248 327486
rect 214928 327218 214970 327454
rect 215206 327218 215248 327454
rect 214928 327134 215248 327218
rect 214928 326898 214970 327134
rect 215206 326898 215248 327134
rect 214928 326866 215248 326898
rect 245648 327454 245968 327486
rect 245648 327218 245690 327454
rect 245926 327218 245968 327454
rect 245648 327134 245968 327218
rect 245648 326898 245690 327134
rect 245926 326898 245968 327134
rect 245648 326866 245968 326898
rect 276368 327454 276688 327486
rect 276368 327218 276410 327454
rect 276646 327218 276688 327454
rect 276368 327134 276688 327218
rect 276368 326898 276410 327134
rect 276646 326898 276688 327134
rect 276368 326866 276688 326898
rect 292619 311948 292685 311949
rect 292619 311884 292620 311948
rect 292684 311884 292685 311948
rect 292619 311883 292685 311884
rect 199568 295954 199888 295986
rect 199568 295718 199610 295954
rect 199846 295718 199888 295954
rect 199568 295634 199888 295718
rect 199568 295398 199610 295634
rect 199846 295398 199888 295634
rect 199568 295366 199888 295398
rect 230288 295954 230608 295986
rect 230288 295718 230330 295954
rect 230566 295718 230608 295954
rect 230288 295634 230608 295718
rect 230288 295398 230330 295634
rect 230566 295398 230608 295634
rect 230288 295366 230608 295398
rect 261008 295954 261328 295986
rect 261008 295718 261050 295954
rect 261286 295718 261328 295954
rect 261008 295634 261328 295718
rect 261008 295398 261050 295634
rect 261286 295398 261328 295634
rect 261008 295366 261328 295398
rect 184208 291454 184528 291486
rect 184208 291218 184250 291454
rect 184486 291218 184528 291454
rect 184208 291134 184528 291218
rect 184208 290898 184250 291134
rect 184486 290898 184528 291134
rect 184208 290866 184528 290898
rect 214928 291454 215248 291486
rect 214928 291218 214970 291454
rect 215206 291218 215248 291454
rect 214928 291134 215248 291218
rect 214928 290898 214970 291134
rect 215206 290898 215248 291134
rect 214928 290866 215248 290898
rect 245648 291454 245968 291486
rect 245648 291218 245690 291454
rect 245926 291218 245968 291454
rect 245648 291134 245968 291218
rect 245648 290898 245690 291134
rect 245926 290898 245968 291134
rect 245648 290866 245968 290898
rect 276368 291454 276688 291486
rect 276368 291218 276410 291454
rect 276646 291218 276688 291454
rect 276368 291134 276688 291218
rect 276368 290898 276410 291134
rect 276646 290898 276688 291134
rect 276368 290866 276688 290898
rect 199568 259954 199888 259986
rect 199568 259718 199610 259954
rect 199846 259718 199888 259954
rect 199568 259634 199888 259718
rect 199568 259398 199610 259634
rect 199846 259398 199888 259634
rect 199568 259366 199888 259398
rect 230288 259954 230608 259986
rect 230288 259718 230330 259954
rect 230566 259718 230608 259954
rect 230288 259634 230608 259718
rect 230288 259398 230330 259634
rect 230566 259398 230608 259634
rect 230288 259366 230608 259398
rect 261008 259954 261328 259986
rect 261008 259718 261050 259954
rect 261286 259718 261328 259954
rect 261008 259634 261328 259718
rect 261008 259398 261050 259634
rect 261286 259398 261328 259634
rect 261008 259366 261328 259398
rect 184208 255454 184528 255486
rect 184208 255218 184250 255454
rect 184486 255218 184528 255454
rect 184208 255134 184528 255218
rect 184208 254898 184250 255134
rect 184486 254898 184528 255134
rect 184208 254866 184528 254898
rect 214928 255454 215248 255486
rect 214928 255218 214970 255454
rect 215206 255218 215248 255454
rect 214928 255134 215248 255218
rect 214928 254898 214970 255134
rect 215206 254898 215248 255134
rect 214928 254866 215248 254898
rect 245648 255454 245968 255486
rect 245648 255218 245690 255454
rect 245926 255218 245968 255454
rect 245648 255134 245968 255218
rect 245648 254898 245690 255134
rect 245926 254898 245968 255134
rect 245648 254866 245968 254898
rect 276368 255454 276688 255486
rect 276368 255218 276410 255454
rect 276646 255218 276688 255454
rect 276368 255134 276688 255218
rect 276368 254898 276410 255134
rect 276646 254898 276688 255134
rect 276368 254866 276688 254898
rect 292622 248430 292682 311883
rect 293174 298757 293234 354859
rect 293907 347580 293973 347581
rect 293907 347516 293908 347580
rect 293972 347516 293973 347580
rect 293907 347515 293973 347516
rect 293171 298756 293237 298757
rect 293171 298692 293172 298756
rect 293236 298692 293237 298756
rect 293171 298691 293237 298692
rect 293171 276044 293237 276045
rect 293171 275980 293172 276044
rect 293236 275980 293237 276044
rect 293171 275979 293237 275980
rect 292622 248370 293050 248430
rect 179827 242996 179893 242997
rect 179827 242932 179828 242996
rect 179892 242932 179893 242996
rect 179827 242931 179893 242932
rect 292619 242996 292685 242997
rect 292619 242932 292620 242996
rect 292684 242932 292685 242996
rect 292619 242931 292685 242932
rect 179275 91084 179341 91085
rect 179275 91020 179276 91084
rect 179340 91020 179341 91084
rect 179275 91019 179341 91020
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177067 51780 177133 51781
rect 177067 51716 177068 51780
rect 177132 51716 177133 51780
rect 177067 51715 177133 51716
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 176515 6220 176581 6221
rect 176515 6156 176516 6220
rect 176580 6156 176581 6220
rect 176515 6155 176581 6156
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 -7066 177914 34398
rect 179830 27029 179890 242931
rect 292622 242450 292682 242931
rect 292438 242390 292682 242450
rect 288939 240140 289005 240141
rect 288939 240076 288940 240140
rect 289004 240076 289005 240140
rect 288939 240075 289005 240076
rect 181794 219454 182414 238000
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 179827 27028 179893 27029
rect 179827 26964 179828 27028
rect 179892 26964 179893 27028
rect 179827 26963 179893 26964
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 223954 186914 238000
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 187954 186914 223398
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 115954 186914 151398
rect 186294 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 186914 115954
rect 186294 115634 186914 115718
rect 186294 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 186914 115634
rect 186294 79954 186914 115398
rect 186294 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 186914 79954
rect 186294 79634 186914 79718
rect 186294 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 186914 79634
rect 186294 43954 186914 79398
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 228454 191414 238000
rect 190794 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 191414 228454
rect 190794 228134 191414 228218
rect 190794 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 191414 228134
rect 190794 192454 191414 227898
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 120454 191414 155898
rect 190794 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 191414 120454
rect 190794 120134 191414 120218
rect 190794 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 191414 120134
rect 190794 84454 191414 119898
rect 190794 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 191414 84454
rect 190794 84134 191414 84218
rect 190794 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 191414 84134
rect 190794 48454 191414 83898
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 232954 195914 238000
rect 195294 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 195914 232954
rect 195294 232634 195914 232718
rect 195294 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 195914 232634
rect 195294 196954 195914 232398
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 237454 200414 238000
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 205954 204914 238000
rect 208163 237420 208229 237421
rect 208163 237356 208164 237420
rect 208228 237356 208229 237420
rect 208163 237355 208229 237356
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 208166 24173 208226 237355
rect 208794 210454 209414 238000
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208163 24172 208229 24173
rect 208163 24108 208164 24172
rect 208228 24108 208229 24172
rect 208163 24107 208229 24108
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 214954 213914 238000
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 217794 219454 218414 238000
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 178000 218414 182898
rect 222294 223954 222914 238000
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 178000 222914 187398
rect 226794 228454 227414 238000
rect 226794 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 227414 228454
rect 226794 228134 227414 228218
rect 226794 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 227414 228134
rect 226794 192454 227414 227898
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 178000 227414 191898
rect 231294 232954 231914 238000
rect 231294 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 231914 232954
rect 231294 232634 231914 232718
rect 231294 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 231914 232634
rect 231294 196954 231914 232398
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 178000 231914 196398
rect 235794 237454 236414 238000
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 178000 236414 200898
rect 249294 214954 249914 238000
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249011 179212 249077 179213
rect 249011 179148 249012 179212
rect 249076 179148 249077 179212
rect 249011 179147 249077 179148
rect 249014 177850 249074 179147
rect 249294 178954 249914 214398
rect 253794 219454 254414 238000
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 252507 188460 252573 188461
rect 252507 188396 252508 188460
rect 252572 188396 252573 188460
rect 252507 188395 252573 188396
rect 251219 181524 251285 181525
rect 251219 181460 251220 181524
rect 251284 181460 251285 181524
rect 251219 181459 251285 181460
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 178000 249914 178398
rect 249014 177790 249442 177850
rect 249195 177580 249261 177581
rect 249195 177516 249196 177580
rect 249260 177516 249261 177580
rect 249195 177515 249261 177516
rect 249198 173773 249258 177515
rect 249382 174725 249442 177790
rect 249379 174724 249445 174725
rect 249379 174660 249380 174724
rect 249444 174660 249445 174724
rect 249379 174659 249445 174660
rect 249195 173772 249261 173773
rect 249195 173708 249196 173772
rect 249260 173708 249261 173772
rect 249195 173707 249261 173708
rect 227874 151954 228194 151986
rect 227874 151718 227916 151954
rect 228152 151718 228194 151954
rect 227874 151634 228194 151718
rect 227874 151398 227916 151634
rect 228152 151398 228194 151634
rect 227874 151366 228194 151398
rect 237805 151954 238125 151986
rect 237805 151718 237847 151954
rect 238083 151718 238125 151954
rect 237805 151634 238125 151718
rect 237805 151398 237847 151634
rect 238083 151398 238125 151634
rect 237805 151366 238125 151398
rect 251222 147933 251282 181459
rect 252510 170101 252570 188395
rect 253794 183454 254414 218898
rect 258294 223954 258914 238000
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 255267 218652 255333 218653
rect 255267 218588 255268 218652
rect 255332 218588 255333 218652
rect 255267 218587 255333 218588
rect 254531 189684 254597 189685
rect 254531 189620 254532 189684
rect 254596 189620 254597 189684
rect 254531 189619 254597 189620
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 252691 176084 252757 176085
rect 252691 176020 252692 176084
rect 252756 176020 252757 176084
rect 252691 176019 252757 176020
rect 252507 170100 252573 170101
rect 252507 170036 252508 170100
rect 252572 170036 252573 170100
rect 252507 170035 252573 170036
rect 252694 157317 252754 176019
rect 252691 157316 252757 157317
rect 252691 157252 252692 157316
rect 252756 157252 252757 157316
rect 252691 157251 252757 157252
rect 251955 148204 252021 148205
rect 251955 148140 251956 148204
rect 252020 148140 252021 148204
rect 251955 148139 252021 148140
rect 251219 147932 251285 147933
rect 251219 147868 251220 147932
rect 251284 147868 251285 147932
rect 251219 147867 251285 147868
rect 222910 147454 223230 147486
rect 222910 147218 222952 147454
rect 223188 147218 223230 147454
rect 222910 147134 223230 147218
rect 222910 146898 222952 147134
rect 223188 146898 223230 147134
rect 222910 146866 223230 146898
rect 232840 147454 233160 147486
rect 232840 147218 232882 147454
rect 233118 147218 233160 147454
rect 232840 147134 233160 147218
rect 232840 146898 232882 147134
rect 233118 146898 233160 147134
rect 232840 146866 233160 146898
rect 242771 147454 243091 147486
rect 242771 147218 242813 147454
rect 243049 147218 243091 147454
rect 242771 147134 243091 147218
rect 242771 146898 242813 147134
rect 243049 146898 243091 147134
rect 242771 146866 243091 146898
rect 251771 146300 251837 146301
rect 251771 146236 251772 146300
rect 251836 146236 251837 146300
rect 251771 146235 251837 146236
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 214419 132700 214485 132701
rect 214419 132636 214420 132700
rect 214484 132636 214485 132700
rect 214419 132635 214485 132636
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 214422 93125 214482 132635
rect 227874 115954 228194 115986
rect 227874 115718 227916 115954
rect 228152 115718 228194 115954
rect 227874 115634 228194 115718
rect 227874 115398 227916 115634
rect 228152 115398 228194 115634
rect 227874 115366 228194 115398
rect 237805 115954 238125 115986
rect 237805 115718 237847 115954
rect 238083 115718 238125 115954
rect 237805 115634 238125 115718
rect 237805 115398 237847 115634
rect 238083 115398 238125 115634
rect 237805 115366 238125 115398
rect 222910 111454 223230 111486
rect 222910 111218 222952 111454
rect 223188 111218 223230 111454
rect 222910 111134 223230 111218
rect 222910 110898 222952 111134
rect 223188 110898 223230 111134
rect 222910 110866 223230 110898
rect 232840 111454 233160 111486
rect 232840 111218 232882 111454
rect 233118 111218 233160 111454
rect 232840 111134 233160 111218
rect 232840 110898 232882 111134
rect 233118 110898 233160 111134
rect 232840 110866 233160 110898
rect 242771 111454 243091 111486
rect 242771 111218 242813 111454
rect 243049 111218 243091 111454
rect 242771 111134 243091 111218
rect 251774 111213 251834 146235
rect 251958 127669 252018 148139
rect 253794 147454 254414 182898
rect 254534 174317 254594 189619
rect 254531 174316 254597 174317
rect 254531 174252 254532 174316
rect 254596 174252 254597 174316
rect 254531 174251 254597 174252
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253243 138412 253309 138413
rect 253243 138348 253244 138412
rect 253308 138348 253309 138412
rect 253243 138347 253309 138348
rect 251955 127668 252021 127669
rect 251955 127604 251956 127668
rect 252020 127604 252021 127668
rect 251955 127603 252021 127604
rect 253246 122850 253306 138347
rect 253062 122790 253306 122850
rect 251771 111212 251837 111213
rect 251771 111148 251772 111212
rect 251836 111148 251837 111212
rect 251771 111147 251837 111148
rect 242771 110898 242813 111134
rect 243049 110898 243091 111134
rect 242771 110866 243091 110898
rect 214603 101556 214669 101557
rect 214603 101492 214604 101556
rect 214668 101492 214669 101556
rect 214603 101491 214669 101492
rect 214419 93124 214485 93125
rect 214419 93060 214420 93124
rect 214484 93060 214485 93124
rect 214419 93059 214485 93060
rect 214606 90949 214666 101491
rect 219203 95980 219269 95981
rect 219203 95916 219204 95980
rect 219268 95916 219269 95980
rect 219203 95915 219269 95916
rect 214603 90948 214669 90949
rect 214603 90884 214604 90948
rect 214668 90884 214669 90948
rect 214603 90883 214669 90884
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 75454 218414 94000
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 219206 3365 219266 95915
rect 222294 79954 222914 94000
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 219203 3364 219269 3365
rect 219203 3300 219204 3364
rect 219268 3300 219269 3364
rect 219203 3299 219269 3300
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 84454 227414 94000
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 88954 231914 94000
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 93454 236414 94000
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 61954 240914 94000
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 66454 245414 94000
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 70954 249914 94000
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 253062 26893 253122 122790
rect 253794 111454 254414 146898
rect 255270 140861 255330 218587
rect 256739 203556 256805 203557
rect 256739 203492 256740 203556
rect 256804 203492 256805 203556
rect 256739 203491 256805 203492
rect 255451 176492 255517 176493
rect 255451 176428 255452 176492
rect 255516 176428 255517 176492
rect 255451 176427 255517 176428
rect 255454 150245 255514 176427
rect 255451 150244 255517 150245
rect 255451 150180 255452 150244
rect 255516 150180 255517 150244
rect 255451 150179 255517 150180
rect 255819 146300 255885 146301
rect 255819 146236 255820 146300
rect 255884 146236 255885 146300
rect 255819 146235 255885 146236
rect 255267 140860 255333 140861
rect 255267 140796 255268 140860
rect 255332 140796 255333 140860
rect 255267 140795 255333 140796
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253059 26892 253125 26893
rect 253059 26828 253060 26892
rect 253124 26828 253125 26892
rect 253059 26827 253125 26828
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 3454 254414 38898
rect 255822 3501 255882 146235
rect 256742 141813 256802 203491
rect 256923 191044 256989 191045
rect 256923 190980 256924 191044
rect 256988 190980 256989 191044
rect 256923 190979 256989 190980
rect 256926 161125 256986 190979
rect 258294 187954 258914 223398
rect 262794 228454 263414 238000
rect 262794 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 263414 228454
rect 262794 228134 263414 228218
rect 262794 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 263414 228134
rect 262794 192454 263414 227898
rect 267294 232954 267914 238000
rect 267294 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 267914 232954
rect 267294 232634 267914 232718
rect 267294 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 267914 232634
rect 265571 227764 265637 227765
rect 265571 227700 265572 227764
rect 265636 227700 265637 227764
rect 265571 227699 265637 227700
rect 263547 204916 263613 204917
rect 263547 204852 263548 204916
rect 263612 204852 263613 204916
rect 263547 204851 263613 204852
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 259499 188324 259565 188325
rect 259499 188260 259500 188324
rect 259564 188260 259565 188324
rect 259499 188259 259565 188260
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 257843 175948 257909 175949
rect 257843 175884 257844 175948
rect 257908 175884 257909 175948
rect 257843 175883 257909 175884
rect 257846 168605 257906 175883
rect 257843 168604 257909 168605
rect 257843 168540 257844 168604
rect 257908 168540 257909 168604
rect 257843 168539 257909 168540
rect 256923 161124 256989 161125
rect 256923 161060 256924 161124
rect 256988 161060 256989 161124
rect 256923 161059 256989 161060
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 256739 141812 256805 141813
rect 256739 141748 256740 141812
rect 256804 141748 256805 141812
rect 256739 141747 256805 141748
rect 257843 129028 257909 129029
rect 257843 128964 257844 129028
rect 257908 128964 257909 129028
rect 257843 128963 257909 128964
rect 257846 3501 257906 128963
rect 258294 115954 258914 151398
rect 259502 138277 259562 188259
rect 261155 183020 261221 183021
rect 261155 182956 261156 183020
rect 261220 182956 261221 183020
rect 261155 182955 261221 182956
rect 260787 181660 260853 181661
rect 260787 181596 260788 181660
rect 260852 181596 260853 181660
rect 260787 181595 260853 181596
rect 259683 177444 259749 177445
rect 259683 177380 259684 177444
rect 259748 177380 259749 177444
rect 259683 177379 259749 177380
rect 259686 142629 259746 177379
rect 260790 171150 260850 181595
rect 260790 171090 261034 171150
rect 259683 142628 259749 142629
rect 259683 142564 259684 142628
rect 259748 142564 259749 142628
rect 259683 142563 259749 142564
rect 259499 138276 259565 138277
rect 259499 138212 259500 138276
rect 259564 138212 259565 138276
rect 259499 138211 259565 138212
rect 260974 136645 261034 171090
rect 261158 163029 261218 182955
rect 262259 181388 262325 181389
rect 262259 181324 262260 181388
rect 262324 181324 262325 181388
rect 262259 181323 262325 181324
rect 261155 163028 261221 163029
rect 261155 162964 261156 163028
rect 261220 162964 261221 163028
rect 261155 162963 261221 162964
rect 262262 157997 262322 181323
rect 262259 157996 262325 157997
rect 262259 157932 262260 157996
rect 262324 157932 262325 157996
rect 262259 157931 262325 157932
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 260971 136644 261037 136645
rect 260971 136580 260972 136644
rect 261036 136580 261037 136644
rect 260971 136579 261037 136580
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 255819 3500 255885 3501
rect 255819 3436 255820 3500
rect 255884 3436 255885 3500
rect 255819 3435 255885 3436
rect 257843 3500 257909 3501
rect 257843 3436 257844 3500
rect 257908 3436 257909 3500
rect 257843 3435 257909 3436
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 120454 263414 155898
rect 263550 138005 263610 204851
rect 264099 189820 264165 189821
rect 264099 189756 264100 189820
rect 264164 189756 264165 189820
rect 264099 189755 264165 189756
rect 263547 138004 263613 138005
rect 263547 137940 263548 138004
rect 263612 137940 263613 138004
rect 263547 137939 263613 137940
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 264102 3365 264162 189755
rect 265019 187100 265085 187101
rect 265019 187036 265020 187100
rect 265084 187036 265085 187100
rect 265019 187035 265085 187036
rect 265022 159629 265082 187035
rect 265019 159628 265085 159629
rect 265019 159564 265020 159628
rect 265084 159564 265085 159628
rect 265019 159563 265085 159564
rect 265574 86869 265634 227699
rect 267294 196954 267914 232398
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 266307 191180 266373 191181
rect 266307 191116 266308 191180
rect 266372 191116 266373 191180
rect 266307 191115 266373 191116
rect 266310 145621 266370 191115
rect 267294 160954 267914 196398
rect 271794 237454 272414 238000
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 269067 195260 269133 195261
rect 269067 195196 269068 195260
rect 269132 195196 269133 195260
rect 269067 195195 269133 195196
rect 269070 163165 269130 195195
rect 271091 175948 271157 175949
rect 271091 175884 271092 175948
rect 271156 175884 271157 175948
rect 271091 175883 271157 175884
rect 269067 163164 269133 163165
rect 269067 163100 269068 163164
rect 269132 163100 269133 163164
rect 269067 163099 269133 163100
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 266307 145620 266373 145621
rect 266307 145556 266308 145620
rect 266372 145556 266373 145620
rect 266307 145555 266373 145556
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 271094 101421 271154 175883
rect 271794 165454 272414 200898
rect 276294 205954 276914 238000
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 275139 193900 275205 193901
rect 275139 193836 275140 193900
rect 275204 193836 275205 193900
rect 275139 193835 275205 193836
rect 273851 178124 273917 178125
rect 273851 178060 273852 178124
rect 273916 178060 273917 178124
rect 273851 178059 273917 178060
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271091 101420 271157 101421
rect 271091 101356 271092 101420
rect 271156 101356 271157 101420
rect 271091 101355 271157 101356
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 265571 86868 265637 86869
rect 265571 86804 265572 86868
rect 265636 86804 265637 86868
rect 265571 86803 265637 86804
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 264099 3364 264165 3365
rect 264099 3300 264100 3364
rect 264164 3300 264165 3364
rect 264099 3299 264165 3300
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 93454 272414 128898
rect 273854 97885 273914 178059
rect 273851 97884 273917 97885
rect 273851 97820 273852 97884
rect 273916 97820 273917 97884
rect 273851 97819 273917 97820
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 275142 3501 275202 193835
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 275139 3500 275205 3501
rect 275139 3436 275140 3500
rect 275204 3436 275205 3500
rect 275139 3435 275205 3436
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 210454 281414 238000
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 285294 214954 285914 238000
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 283419 112164 283485 112165
rect 283419 112100 283420 112164
rect 283484 112100 283485 112164
rect 283419 112099 283485 112100
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 283422 40629 283482 112099
rect 285294 106954 285914 142398
rect 287651 125900 287717 125901
rect 287651 125836 287652 125900
rect 287716 125836 287717 125900
rect 287651 125835 287717 125836
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 283419 40628 283485 40629
rect 283419 40564 283420 40628
rect 283484 40564 283485 40628
rect 283419 40563 283485 40564
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 34954 285914 70398
rect 287654 66877 287714 125835
rect 287651 66876 287717 66877
rect 287651 66812 287652 66876
rect 287716 66812 287717 66876
rect 287651 66811 287717 66812
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 288942 6357 289002 240075
rect 292438 238770 292498 242390
rect 292990 238770 293050 248370
rect 291702 238710 292498 238770
rect 292622 238710 293050 238770
rect 289794 219454 290414 238000
rect 291702 226269 291762 238710
rect 292622 230485 292682 238710
rect 293174 238509 293234 275979
rect 293171 238508 293237 238509
rect 293171 238444 293172 238508
rect 293236 238444 293237 238508
rect 293171 238443 293237 238444
rect 292619 230484 292685 230485
rect 292619 230420 292620 230484
rect 292684 230420 292685 230484
rect 292619 230419 292685 230420
rect 291699 226268 291765 226269
rect 291699 226204 291700 226268
rect 291764 226204 291765 226268
rect 291699 226203 291765 226204
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 288939 6356 289005 6357
rect 288939 6292 288940 6356
rect 289004 6292 289005 6356
rect 288939 6291 289005 6292
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 3454 290414 38898
rect 293910 26893 293970 347515
rect 294094 240141 294154 358803
rect 294294 357154 294914 367398
rect 295934 365805 295994 702475
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 552454 299414 587898
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 298794 516454 299414 551898
rect 298794 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 299414 516454
rect 298794 516134 299414 516218
rect 298794 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 299414 516134
rect 298794 480454 299414 515898
rect 298794 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 299414 480454
rect 298794 480134 299414 480218
rect 298794 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 299414 480134
rect 298794 444454 299414 479898
rect 298794 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 299414 444454
rect 298794 444134 299414 444218
rect 298794 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 299414 444134
rect 298794 408454 299414 443898
rect 298794 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 299414 408454
rect 298794 408134 299414 408218
rect 298794 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 299414 408134
rect 298794 372454 299414 407898
rect 298794 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 299414 372454
rect 298794 372134 299414 372218
rect 298794 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 299414 372134
rect 295931 365804 295997 365805
rect 295931 365740 295932 365804
rect 295996 365740 295997 365804
rect 295931 365739 295997 365740
rect 295934 354690 295994 365739
rect 295750 354630 295994 354690
rect 295379 352340 295445 352341
rect 295379 352276 295380 352340
rect 295444 352276 295445 352340
rect 295379 352275 295445 352276
rect 294091 240140 294157 240141
rect 294091 240076 294092 240140
rect 294156 240076 294157 240140
rect 294091 240075 294157 240076
rect 294294 223954 294914 238000
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 295382 104141 295442 352275
rect 295750 343501 295810 354630
rect 295747 343500 295813 343501
rect 295747 343436 295748 343500
rect 295812 343436 295813 343500
rect 295747 343435 295813 343436
rect 295750 341461 295810 343435
rect 295747 341460 295813 341461
rect 295747 341396 295748 341460
rect 295812 341396 295813 341460
rect 295747 341395 295813 341396
rect 298794 336454 299414 371898
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 298794 300454 299414 335898
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 296667 248436 296733 248437
rect 296667 248430 296668 248436
rect 296486 248372 296668 248430
rect 296732 248372 296733 248436
rect 296486 248371 296733 248372
rect 296486 248370 296730 248371
rect 296486 234429 296546 248370
rect 296483 234428 296549 234429
rect 296483 234364 296484 234428
rect 296548 234364 296549 234428
rect 296483 234363 296549 234364
rect 298794 228454 299414 263898
rect 298794 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 299414 228454
rect 298794 228134 299414 228218
rect 298794 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 299414 228134
rect 298794 192454 299414 227898
rect 298794 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 299414 192454
rect 298794 192134 299414 192218
rect 298794 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 299414 192134
rect 298794 156454 299414 191898
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 556954 303914 592398
rect 303294 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 303914 556954
rect 303294 556634 303914 556718
rect 303294 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 303914 556634
rect 303294 520954 303914 556398
rect 303294 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 303914 520954
rect 303294 520634 303914 520718
rect 303294 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 303914 520634
rect 303294 484954 303914 520398
rect 303294 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 303914 484954
rect 303294 484634 303914 484718
rect 303294 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 303914 484634
rect 303294 448954 303914 484398
rect 303294 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 303914 448954
rect 303294 448634 303914 448718
rect 303294 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 303914 448634
rect 303294 412954 303914 448398
rect 303294 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 303914 412954
rect 303294 412634 303914 412718
rect 303294 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 303914 412634
rect 303294 376954 303914 412398
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 303294 340954 303914 376398
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 303294 304954 303914 340398
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 232954 303914 268398
rect 303294 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 303914 232954
rect 303294 232634 303914 232718
rect 303294 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 303914 232634
rect 303294 196954 303914 232398
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 178000 308414 200898
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 529954 312914 565398
rect 312294 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 312914 529954
rect 312294 529634 312914 529718
rect 312294 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 312914 529634
rect 312294 493954 312914 529398
rect 312294 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 312914 493954
rect 312294 493634 312914 493718
rect 312294 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 312914 493634
rect 312294 457954 312914 493398
rect 312294 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 312914 457954
rect 312294 457634 312914 457718
rect 312294 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 312914 457634
rect 312294 421954 312914 457398
rect 312294 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 312914 421954
rect 312294 421634 312914 421718
rect 312294 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 312914 421634
rect 312294 385954 312914 421398
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 313954 312914 349398
rect 312294 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 312914 313954
rect 312294 313634 312914 313718
rect 312294 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 312914 313634
rect 312294 277954 312914 313398
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 241954 312914 277398
rect 312294 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 312914 241954
rect 312294 241634 312914 241718
rect 312294 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 312914 241634
rect 312294 205954 312914 241398
rect 312294 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 312914 205954
rect 312294 205634 312914 205718
rect 312294 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 312914 205634
rect 312294 178000 312914 205398
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 534454 317414 569898
rect 316794 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 317414 534454
rect 316794 534134 317414 534218
rect 316794 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 317414 534134
rect 316794 498454 317414 533898
rect 316794 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 317414 498454
rect 316794 498134 317414 498218
rect 316794 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 317414 498134
rect 316794 462454 317414 497898
rect 316794 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 317414 462454
rect 316794 462134 317414 462218
rect 316794 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 317414 462134
rect 316794 426454 317414 461898
rect 316794 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 317414 426454
rect 316794 426134 317414 426218
rect 316794 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 317414 426134
rect 316794 390454 317414 425898
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 318454 317414 353898
rect 316794 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 317414 318454
rect 316794 318134 317414 318218
rect 316794 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 317414 318134
rect 316794 282454 317414 317898
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 246454 317414 281898
rect 316794 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 317414 246454
rect 316794 246134 317414 246218
rect 316794 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 317414 246134
rect 316794 210454 317414 245898
rect 316794 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 317414 210454
rect 316794 210134 317414 210218
rect 316794 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 317414 210134
rect 316794 178000 317414 209898
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 538954 321914 574398
rect 321294 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 321914 538954
rect 321294 538634 321914 538718
rect 321294 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 321914 538634
rect 321294 502954 321914 538398
rect 321294 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 321914 502954
rect 321294 502634 321914 502718
rect 321294 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 321914 502634
rect 321294 466954 321914 502398
rect 321294 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 321914 466954
rect 321294 466634 321914 466718
rect 321294 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 321914 466634
rect 321294 430954 321914 466398
rect 321294 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 321914 430954
rect 321294 430634 321914 430718
rect 321294 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 321914 430634
rect 321294 394954 321914 430398
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 322954 321914 358398
rect 321294 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 321914 322954
rect 321294 322634 321914 322718
rect 321294 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 321914 322634
rect 321294 286954 321914 322398
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 214954 321914 250398
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 322059 232524 322125 232525
rect 322059 232460 322060 232524
rect 322124 232460 322125 232524
rect 322059 232459 322125 232460
rect 321294 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 321914 214954
rect 321294 214634 321914 214718
rect 321294 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 321914 214634
rect 320219 186964 320285 186965
rect 320219 186900 320220 186964
rect 320284 186900 320285 186964
rect 320219 186899 320285 186900
rect 306971 175268 307037 175269
rect 306971 175204 306972 175268
rect 307036 175204 307037 175268
rect 306971 175203 307037 175204
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 299979 132700 300045 132701
rect 299979 132636 299980 132700
rect 300044 132636 300045 132700
rect 299979 132635 300045 132636
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 295379 104140 295445 104141
rect 295379 104076 295380 104140
rect 295444 104076 295445 104140
rect 295379 104075 295445 104076
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 293907 26892 293973 26893
rect 293907 26828 293908 26892
rect 293972 26828 293973 26892
rect 293907 26827 293973 26828
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 299982 59941 300042 132635
rect 301451 128484 301517 128485
rect 301451 128420 301452 128484
rect 301516 128420 301517 128484
rect 301451 128419 301517 128420
rect 299979 59940 300045 59941
rect 299979 59876 299980 59940
rect 300044 59876 300045 59940
rect 299979 59875 300045 59876
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 301454 4861 301514 128419
rect 303294 124954 303914 160398
rect 306974 149701 307034 175203
rect 320222 171150 320282 186899
rect 321294 178954 321914 214398
rect 321294 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 321914 178954
rect 321294 178634 321914 178718
rect 321294 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 321914 178634
rect 321294 178000 321914 178398
rect 321323 176764 321389 176765
rect 321323 176700 321324 176764
rect 321388 176700 321389 176764
rect 321323 176699 321389 176700
rect 321326 172141 321386 176699
rect 321323 172140 321389 172141
rect 321323 172076 321324 172140
rect 321388 172076 321389 172140
rect 321323 172075 321389 172076
rect 320222 171090 321386 171150
rect 321326 170373 321386 171090
rect 321323 170372 321389 170373
rect 321323 170308 321324 170372
rect 321388 170308 321389 170372
rect 321323 170307 321389 170308
rect 307339 157452 307405 157453
rect 307339 157388 307340 157452
rect 307404 157388 307405 157452
rect 307339 157387 307405 157388
rect 307155 150244 307221 150245
rect 307155 150180 307156 150244
rect 307220 150180 307221 150244
rect 307155 150179 307221 150180
rect 306971 149700 307037 149701
rect 306971 149636 306972 149700
rect 307036 149636 307037 149700
rect 306971 149635 307037 149636
rect 305499 139772 305565 139773
rect 305499 139708 305500 139772
rect 305564 139708 305565 139772
rect 305499 139707 305565 139708
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 301635 113660 301701 113661
rect 301635 113596 301636 113660
rect 301700 113596 301701 113660
rect 301635 113595 301701 113596
rect 301638 75173 301698 113595
rect 302739 99652 302805 99653
rect 302739 99588 302740 99652
rect 302804 99588 302805 99652
rect 302739 99587 302805 99588
rect 301635 75172 301701 75173
rect 301635 75108 301636 75172
rect 301700 75108 301701 75172
rect 301635 75107 301701 75108
rect 302742 46205 302802 99587
rect 303294 88954 303914 124398
rect 304211 117876 304277 117877
rect 304211 117812 304212 117876
rect 304276 117812 304277 117876
rect 304211 117811 304277 117812
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 302739 46204 302805 46205
rect 302739 46140 302740 46204
rect 302804 46140 302805 46204
rect 302739 46139 302805 46140
rect 303294 16954 303914 52398
rect 304214 36549 304274 117811
rect 305502 64157 305562 139707
rect 307158 134469 307218 150179
rect 307342 145621 307402 157387
rect 314208 151954 314528 151986
rect 314208 151718 314250 151954
rect 314486 151718 314528 151954
rect 314208 151634 314528 151718
rect 314208 151398 314250 151634
rect 314486 151398 314528 151634
rect 314208 151366 314528 151398
rect 317472 151954 317792 151986
rect 317472 151718 317514 151954
rect 317750 151718 317792 151954
rect 317472 151634 317792 151718
rect 317472 151398 317514 151634
rect 317750 151398 317792 151634
rect 317472 151366 317792 151398
rect 322062 148749 322122 232459
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 324267 189140 324333 189141
rect 324267 189076 324268 189140
rect 324332 189076 324333 189140
rect 324267 189075 324333 189076
rect 324270 155549 324330 189075
rect 325794 183454 326414 218898
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 511954 330914 547398
rect 330294 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 330914 511954
rect 330294 511634 330914 511718
rect 330294 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 330914 511634
rect 330294 475954 330914 511398
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 330294 439954 330914 475398
rect 330294 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 330914 439954
rect 330294 439634 330914 439718
rect 330294 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 330914 439634
rect 330294 403954 330914 439398
rect 330294 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 330914 403954
rect 330294 403634 330914 403718
rect 330294 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 330914 403634
rect 330294 367954 330914 403398
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 331954 330914 367398
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 223954 330914 259398
rect 330294 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 330914 223954
rect 330294 223634 330914 223718
rect 330294 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 330914 223634
rect 330294 187954 330914 223398
rect 330294 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 330914 187954
rect 330294 187634 330914 187718
rect 330294 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 330914 187634
rect 326659 187236 326725 187237
rect 326659 187172 326660 187236
rect 326724 187172 326725 187236
rect 326659 187171 326725 187172
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 324267 155548 324333 155549
rect 324267 155484 324268 155548
rect 324332 155484 324333 155548
rect 324267 155483 324333 155484
rect 322059 148748 322125 148749
rect 322059 148684 322060 148748
rect 322124 148684 322125 148748
rect 322059 148683 322125 148684
rect 321507 148068 321573 148069
rect 321507 148004 321508 148068
rect 321572 148004 321573 148068
rect 321507 148003 321573 148004
rect 312576 147454 312896 147486
rect 312576 147218 312618 147454
rect 312854 147218 312896 147454
rect 312576 147134 312896 147218
rect 312576 146898 312618 147134
rect 312854 146898 312896 147134
rect 312576 146866 312896 146898
rect 315840 147454 316160 147486
rect 315840 147218 315882 147454
rect 316118 147218 316160 147454
rect 315840 147134 316160 147218
rect 315840 146898 315882 147134
rect 316118 146898 316160 147134
rect 315840 146866 316160 146898
rect 319104 147454 319424 147486
rect 319104 147218 319146 147454
rect 319382 147218 319424 147454
rect 319104 147134 319424 147218
rect 319104 146898 319146 147134
rect 319382 146898 319424 147134
rect 319104 146866 319424 146898
rect 307339 145620 307405 145621
rect 307339 145556 307340 145620
rect 307404 145556 307405 145620
rect 307339 145555 307405 145556
rect 307707 142084 307773 142085
rect 307707 142020 307708 142084
rect 307772 142020 307773 142084
rect 307707 142019 307773 142020
rect 307710 140045 307770 142019
rect 307707 140044 307773 140045
rect 307707 139980 307708 140044
rect 307772 139980 307773 140044
rect 307707 139979 307773 139980
rect 307155 134468 307221 134469
rect 307155 134404 307156 134468
rect 307220 134404 307221 134468
rect 307155 134403 307221 134404
rect 306971 134060 307037 134061
rect 306971 133996 306972 134060
rect 307036 133996 307037 134060
rect 306971 133995 307037 133996
rect 305683 105908 305749 105909
rect 305683 105844 305684 105908
rect 305748 105844 305749 105908
rect 305683 105843 305749 105844
rect 305499 64156 305565 64157
rect 305499 64092 305500 64156
rect 305564 64092 305565 64156
rect 305499 64091 305565 64092
rect 305686 54501 305746 105843
rect 305683 54500 305749 54501
rect 305683 54436 305684 54500
rect 305748 54436 305749 54500
rect 305683 54435 305749 54436
rect 304211 36548 304277 36549
rect 304211 36484 304212 36548
rect 304276 36484 304277 36548
rect 304211 36483 304277 36484
rect 306974 17237 307034 133995
rect 314208 115954 314528 115986
rect 314208 115718 314250 115954
rect 314486 115718 314528 115954
rect 314208 115634 314528 115718
rect 314208 115398 314250 115634
rect 314486 115398 314528 115634
rect 314208 115366 314528 115398
rect 317472 115954 317792 115986
rect 317472 115718 317514 115954
rect 317750 115718 317792 115954
rect 317472 115634 317792 115718
rect 317472 115398 317514 115634
rect 317750 115398 317792 115634
rect 317472 115366 317792 115398
rect 321510 113190 321570 148003
rect 325794 147454 326414 182898
rect 326662 173909 326722 187171
rect 328499 185060 328565 185061
rect 328499 184996 328500 185060
rect 328564 184996 328565 185060
rect 328499 184995 328565 184996
rect 327579 182884 327645 182885
rect 327579 182820 327580 182884
rect 327644 182820 327645 182884
rect 327579 182819 327645 182820
rect 327027 177308 327093 177309
rect 327027 177244 327028 177308
rect 327092 177244 327093 177308
rect 327027 177243 327093 177244
rect 326659 173908 326725 173909
rect 326659 173844 326660 173908
rect 326724 173844 326725 173908
rect 326659 173843 326725 173844
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 321510 113130 322122 113190
rect 312576 111454 312896 111486
rect 312576 111218 312618 111454
rect 312854 111218 312896 111454
rect 312576 111134 312896 111218
rect 312576 110898 312618 111134
rect 312854 110898 312896 111134
rect 312576 110866 312896 110898
rect 315840 111454 316160 111486
rect 315840 111218 315882 111454
rect 316118 111218 316160 111454
rect 315840 111134 316160 111218
rect 315840 110898 315882 111134
rect 316118 110898 316160 111134
rect 315840 110866 316160 110898
rect 319104 111454 319424 111486
rect 319104 111218 319146 111454
rect 319382 111218 319424 111454
rect 319104 111134 319424 111218
rect 319104 110898 319146 111134
rect 319382 110898 319424 111134
rect 319104 110866 319424 110898
rect 307155 97068 307221 97069
rect 307155 97004 307156 97068
rect 307220 97004 307221 97068
rect 307155 97003 307221 97004
rect 307158 84829 307218 97003
rect 322062 96525 322122 113130
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 324267 104820 324333 104821
rect 324267 104756 324268 104820
rect 324332 104756 324333 104820
rect 324267 104755 324333 104756
rect 322059 96524 322125 96525
rect 322059 96460 322060 96524
rect 322124 96460 322125 96524
rect 322059 96459 322125 96460
rect 307794 93454 308414 94000
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307155 84828 307221 84829
rect 307155 84764 307156 84828
rect 307220 84764 307221 84828
rect 307155 84763 307221 84764
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 306971 17236 307037 17237
rect 306971 17172 306972 17236
rect 307036 17172 307037 17236
rect 306971 17171 307037 17172
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 301451 4860 301517 4861
rect 301451 4796 301452 4860
rect 301516 4796 301517 4860
rect 301451 4795 301517 4796
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 61954 312914 94000
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 66454 317414 94000
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 70954 321914 94000
rect 324270 93261 324330 104755
rect 324451 96660 324517 96661
rect 324451 96596 324452 96660
rect 324516 96596 324517 96660
rect 324451 96595 324517 96596
rect 324454 96389 324514 96595
rect 324451 96388 324517 96389
rect 324451 96324 324452 96388
rect 324516 96324 324517 96388
rect 324451 96323 324517 96324
rect 324267 93260 324333 93261
rect 324267 93196 324268 93260
rect 324332 93196 324333 93260
rect 324267 93195 324333 93196
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 327030 3365 327090 177243
rect 327582 121413 327642 182819
rect 328502 145621 328562 184995
rect 328683 176084 328749 176085
rect 328683 176020 328684 176084
rect 328748 176020 328749 176084
rect 328683 176019 328749 176020
rect 328686 162757 328746 176019
rect 328683 162756 328749 162757
rect 328683 162692 328684 162756
rect 328748 162692 328749 162756
rect 328683 162691 328749 162692
rect 330294 151954 330914 187398
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 552454 335414 587898
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 516454 335414 551898
rect 334794 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 335414 516454
rect 334794 516134 335414 516218
rect 334794 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 335414 516134
rect 334794 480454 335414 515898
rect 334794 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 335414 480454
rect 334794 480134 335414 480218
rect 334794 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 335414 480134
rect 334794 444454 335414 479898
rect 334794 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 335414 444454
rect 334794 444134 335414 444218
rect 334794 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 335414 444134
rect 334794 408454 335414 443898
rect 334794 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 335414 408454
rect 334794 408134 335414 408218
rect 334794 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 335414 408134
rect 334794 372454 335414 407898
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 334794 336454 335414 371898
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 556954 339914 592398
rect 339294 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 339914 556954
rect 339294 556634 339914 556718
rect 339294 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 339914 556634
rect 339294 520954 339914 556398
rect 339294 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 339914 520954
rect 339294 520634 339914 520718
rect 339294 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 339914 520634
rect 339294 484954 339914 520398
rect 339294 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 339914 484954
rect 339294 484634 339914 484718
rect 339294 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 339914 484634
rect 339294 448954 339914 484398
rect 339294 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 339914 448954
rect 339294 448634 339914 448718
rect 339294 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 339914 448634
rect 339294 412954 339914 448398
rect 339294 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 339914 412954
rect 339294 412634 339914 412718
rect 339294 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 339914 412634
rect 339294 376954 339914 412398
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 335859 356148 335925 356149
rect 335859 356084 335860 356148
rect 335924 356084 335925 356148
rect 335859 356083 335925 356084
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 300454 335414 335898
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 228454 335414 263898
rect 334794 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 335414 228454
rect 334794 228134 335414 228218
rect 334794 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 335414 228134
rect 334794 192454 335414 227898
rect 334794 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 335414 192454
rect 334794 192134 335414 192218
rect 334794 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 335414 192134
rect 331811 184244 331877 184245
rect 331811 184180 331812 184244
rect 331876 184180 331877 184244
rect 331811 184179 331877 184180
rect 331814 161261 331874 184179
rect 332547 180028 332613 180029
rect 332547 179964 332548 180028
rect 332612 179964 332613 180028
rect 332547 179963 332613 179964
rect 331811 161260 331877 161261
rect 331811 161196 331812 161260
rect 331876 161196 331877 161260
rect 331811 161195 331877 161196
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 328499 145620 328565 145621
rect 328499 145556 328500 145620
rect 328564 145556 328565 145620
rect 328499 145555 328565 145556
rect 327579 121412 327645 121413
rect 327579 121348 327580 121412
rect 327644 121348 327645 121412
rect 327579 121347 327645 121348
rect 330294 115954 330914 151398
rect 332550 138685 332610 179963
rect 334794 156454 335414 191898
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 332547 138684 332613 138685
rect 332547 138620 332548 138684
rect 332612 138620 332613 138684
rect 332547 138619 332613 138620
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 327027 3364 327093 3365
rect 327027 3300 327028 3364
rect 327092 3300 327093 3364
rect 327027 3299 327093 3300
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 335862 102237 335922 356083
rect 339294 340954 339914 376398
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 304954 339914 340398
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 232954 339914 268398
rect 339294 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 339914 232954
rect 339294 232634 339914 232718
rect 339294 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 339914 232634
rect 339294 196954 339914 232398
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 337331 195260 337397 195261
rect 337331 195196 337332 195260
rect 337396 195196 337397 195260
rect 337331 195195 337397 195196
rect 335859 102236 335925 102237
rect 335859 102172 335860 102236
rect 335924 102172 335925 102236
rect 335859 102171 335925 102172
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 337334 3501 337394 195195
rect 339294 160954 339914 196398
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 342299 175948 342365 175949
rect 342299 175884 342300 175948
rect 342364 175884 342365 175948
rect 342299 175883 342365 175884
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 339294 124954 339914 160398
rect 342302 129029 342362 175883
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 342299 129028 342365 129029
rect 342299 128964 342300 129028
rect 342364 128964 342365 129028
rect 342299 128963 342365 128964
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 337331 3500 337397 3501
rect 337331 3436 337332 3500
rect 337396 3436 337397 3500
rect 337331 3435 337397 3436
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 529954 348914 565398
rect 348294 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 348914 529954
rect 348294 529634 348914 529718
rect 348294 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 348914 529634
rect 348294 493954 348914 529398
rect 348294 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 348914 493954
rect 348294 493634 348914 493718
rect 348294 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 348914 493634
rect 348294 457954 348914 493398
rect 348294 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 348914 457954
rect 348294 457634 348914 457718
rect 348294 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 348914 457634
rect 348294 421954 348914 457398
rect 348294 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 348914 421954
rect 348294 421634 348914 421718
rect 348294 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 348914 421634
rect 348294 385954 348914 421398
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 313954 348914 349398
rect 348294 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 348914 313954
rect 348294 313634 348914 313718
rect 348294 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 348914 313634
rect 348294 277954 348914 313398
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 241954 348914 277398
rect 348294 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 348914 241954
rect 348294 241634 348914 241718
rect 348294 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 348914 241634
rect 348294 205954 348914 241398
rect 348294 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 348914 205954
rect 348294 205634 348914 205718
rect 348294 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 348914 205634
rect 348294 169954 348914 205398
rect 348294 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 348914 169954
rect 348294 169634 348914 169718
rect 348294 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 348914 169634
rect 348294 133954 348914 169398
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 534454 353414 569898
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 352794 498454 353414 533898
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 426454 353414 461898
rect 352794 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 353414 426454
rect 352794 426134 353414 426218
rect 352794 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 353414 426134
rect 352794 390454 353414 425898
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 210454 353414 245898
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 138454 353414 173898
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 538954 357914 574398
rect 357294 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 357914 538954
rect 357294 538634 357914 538718
rect 357294 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 357914 538634
rect 357294 502954 357914 538398
rect 357294 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 357914 502954
rect 357294 502634 357914 502718
rect 357294 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 357914 502634
rect 357294 466954 357914 502398
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 430954 357914 466398
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 357294 430634 357914 430718
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 214954 357914 250398
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388483 311132 388549 311133
rect 388483 311068 388484 311132
rect 388548 311068 388549 311132
rect 388483 311067 388549 311068
rect 387011 301476 387077 301477
rect 387011 301412 387012 301476
rect 387076 301412 387077 301476
rect 387011 301411 387077 301412
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 241954 384914 277398
rect 385539 276316 385605 276317
rect 385539 276252 385540 276316
rect 385604 276252 385605 276316
rect 385539 276251 385605 276252
rect 384294 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 384914 241954
rect 384294 241634 384914 241718
rect 384294 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 384914 241634
rect 384294 205954 384914 241398
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 385542 121413 385602 276251
rect 387014 224637 387074 301411
rect 387011 224636 387077 224637
rect 387011 224572 387012 224636
rect 387076 224572 387077 224636
rect 387011 224571 387077 224572
rect 387014 176357 387074 224571
rect 388299 222188 388365 222189
rect 388299 222124 388300 222188
rect 388364 222124 388365 222188
rect 388299 222123 388365 222124
rect 387011 176356 387077 176357
rect 387011 176292 387012 176356
rect 387076 176292 387077 176356
rect 387011 176291 387077 176292
rect 387563 175948 387629 175949
rect 387563 175884 387564 175948
rect 387628 175884 387629 175948
rect 387563 175883 387629 175884
rect 385539 121412 385605 121413
rect 385539 121348 385540 121412
rect 385604 121348 385605 121412
rect 385539 121347 385605 121348
rect 387195 116516 387261 116517
rect 387195 116452 387196 116516
rect 387260 116452 387261 116516
rect 387195 116451 387261 116452
rect 387011 109716 387077 109717
rect 387011 109652 387012 109716
rect 387076 109652 387077 109716
rect 387011 109651 387077 109652
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 387014 84149 387074 109651
rect 387198 96389 387258 116451
rect 387566 112437 387626 175883
rect 387563 112436 387629 112437
rect 387563 112372 387564 112436
rect 387628 112372 387629 112436
rect 387563 112371 387629 112372
rect 387195 96388 387261 96389
rect 387195 96324 387196 96388
rect 387260 96324 387261 96388
rect 387195 96323 387261 96324
rect 387011 84148 387077 84149
rect 387011 84084 387012 84148
rect 387076 84084 387077 84148
rect 387011 84083 387077 84084
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 388302 19413 388362 222123
rect 388486 213893 388546 311067
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 278000 389414 281898
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 390691 280532 390757 280533
rect 390691 280468 390692 280532
rect 390756 280468 390757 280532
rect 390691 280467 390757 280468
rect 389771 276180 389837 276181
rect 389771 276116 389772 276180
rect 389836 276116 389837 276180
rect 389771 276115 389837 276116
rect 389774 238781 389834 276115
rect 390507 275636 390573 275637
rect 390507 275572 390508 275636
rect 390572 275572 390573 275636
rect 390507 275571 390573 275572
rect 390510 274277 390570 275571
rect 390507 274276 390573 274277
rect 390507 274212 390508 274276
rect 390572 274212 390573 274276
rect 390507 274211 390573 274212
rect 390694 273050 390754 280467
rect 393294 278000 393914 286398
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 278000 398414 290898
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 278000 402914 295398
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 278000 407414 299898
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 278000 411914 304398
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 278000 416414 308898
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 278000 420914 313398
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 278000 425414 281898
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 278000 429914 286398
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 278000 434414 290898
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 278000 438914 295398
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 278000 443414 299898
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 278000 447914 304398
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 278000 452414 308898
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 278000 456914 313398
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 278000 461414 281898
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 278000 465914 286398
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 278000 470414 290898
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 278000 474914 295398
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 278000 479414 299898
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 278000 483914 304398
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 278000 488414 308898
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 278000 492914 313398
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 278000 497414 281898
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 278000 501914 286398
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 278000 506414 290898
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 278000 510914 295398
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 278000 515414 299898
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 278000 519914 304398
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 278000 524414 308898
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 278000 528914 313398
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 278000 533414 281898
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 278000 537914 286398
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 278000 542414 290898
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 278000 546914 295398
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 278000 551414 299898
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 278000 555914 304398
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 278000 560414 308898
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 278000 564914 313398
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 570091 364444 570157 364445
rect 570091 364380 570092 364444
rect 570156 364380 570157 364444
rect 570091 364379 570157 364380
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568619 285700 568685 285701
rect 568619 285636 568620 285700
rect 568684 285636 568685 285700
rect 568619 285635 568685 285636
rect 502011 275636 502077 275637
rect 502011 275572 502012 275636
rect 502076 275572 502077 275636
rect 502011 275571 502077 275572
rect 502014 274685 502074 275571
rect 502011 274684 502077 274685
rect 502011 274620 502012 274684
rect 502076 274620 502077 274684
rect 502011 274619 502077 274620
rect 568622 274549 568682 285635
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 278000 569414 281898
rect 569539 278764 569605 278765
rect 569539 278700 569540 278764
rect 569604 278700 569605 278764
rect 569539 278699 569605 278700
rect 568619 274548 568685 274549
rect 568619 274484 568620 274548
rect 568684 274484 568685 274548
rect 568619 274483 568685 274484
rect 390510 272990 390754 273050
rect 390510 272509 390570 272990
rect 390507 272508 390573 272509
rect 390507 272444 390508 272508
rect 390572 272444 390573 272508
rect 390507 272443 390573 272444
rect 409568 259954 409888 259986
rect 409568 259718 409610 259954
rect 409846 259718 409888 259954
rect 409568 259634 409888 259718
rect 409568 259398 409610 259634
rect 409846 259398 409888 259634
rect 409568 259366 409888 259398
rect 440288 259954 440608 259986
rect 440288 259718 440330 259954
rect 440566 259718 440608 259954
rect 440288 259634 440608 259718
rect 440288 259398 440330 259634
rect 440566 259398 440608 259634
rect 440288 259366 440608 259398
rect 471008 259954 471328 259986
rect 471008 259718 471050 259954
rect 471286 259718 471328 259954
rect 471008 259634 471328 259718
rect 471008 259398 471050 259634
rect 471286 259398 471328 259634
rect 471008 259366 471328 259398
rect 501728 259954 502048 259986
rect 501728 259718 501770 259954
rect 502006 259718 502048 259954
rect 501728 259634 502048 259718
rect 501728 259398 501770 259634
rect 502006 259398 502048 259634
rect 501728 259366 502048 259398
rect 532448 259954 532768 259986
rect 532448 259718 532490 259954
rect 532726 259718 532768 259954
rect 532448 259634 532768 259718
rect 532448 259398 532490 259634
rect 532726 259398 532768 259634
rect 532448 259366 532768 259398
rect 563168 259954 563488 259986
rect 563168 259718 563210 259954
rect 563446 259718 563488 259954
rect 563168 259634 563488 259718
rect 563168 259398 563210 259634
rect 563446 259398 563488 259634
rect 563168 259366 563488 259398
rect 394208 255454 394528 255486
rect 394208 255218 394250 255454
rect 394486 255218 394528 255454
rect 394208 255134 394528 255218
rect 394208 254898 394250 255134
rect 394486 254898 394528 255134
rect 394208 254866 394528 254898
rect 424928 255454 425248 255486
rect 424928 255218 424970 255454
rect 425206 255218 425248 255454
rect 424928 255134 425248 255218
rect 424928 254898 424970 255134
rect 425206 254898 425248 255134
rect 424928 254866 425248 254898
rect 455648 255454 455968 255486
rect 455648 255218 455690 255454
rect 455926 255218 455968 255454
rect 455648 255134 455968 255218
rect 455648 254898 455690 255134
rect 455926 254898 455968 255134
rect 455648 254866 455968 254898
rect 486368 255454 486688 255486
rect 486368 255218 486410 255454
rect 486646 255218 486688 255454
rect 486368 255134 486688 255218
rect 486368 254898 486410 255134
rect 486646 254898 486688 255134
rect 486368 254866 486688 254898
rect 517088 255454 517408 255486
rect 517088 255218 517130 255454
rect 517366 255218 517408 255454
rect 517088 255134 517408 255218
rect 517088 254898 517130 255134
rect 517366 254898 517408 255134
rect 517088 254866 517408 254898
rect 547808 255454 548128 255486
rect 547808 255218 547850 255454
rect 548086 255218 548128 255454
rect 547808 255134 548128 255218
rect 547808 254898 547850 255134
rect 548086 254898 548128 255134
rect 547808 254866 548128 254898
rect 389771 238780 389837 238781
rect 389771 238716 389772 238780
rect 389836 238716 389837 238780
rect 389771 238715 389837 238716
rect 409568 223954 409888 223986
rect 409568 223718 409610 223954
rect 409846 223718 409888 223954
rect 409568 223634 409888 223718
rect 409568 223398 409610 223634
rect 409846 223398 409888 223634
rect 409568 223366 409888 223398
rect 440288 223954 440608 223986
rect 440288 223718 440330 223954
rect 440566 223718 440608 223954
rect 440288 223634 440608 223718
rect 440288 223398 440330 223634
rect 440566 223398 440608 223634
rect 440288 223366 440608 223398
rect 471008 223954 471328 223986
rect 471008 223718 471050 223954
rect 471286 223718 471328 223954
rect 471008 223634 471328 223718
rect 471008 223398 471050 223634
rect 471286 223398 471328 223634
rect 471008 223366 471328 223398
rect 501728 223954 502048 223986
rect 501728 223718 501770 223954
rect 502006 223718 502048 223954
rect 501728 223634 502048 223718
rect 501728 223398 501770 223634
rect 502006 223398 502048 223634
rect 501728 223366 502048 223398
rect 532448 223954 532768 223986
rect 532448 223718 532490 223954
rect 532726 223718 532768 223954
rect 532448 223634 532768 223718
rect 532448 223398 532490 223634
rect 532726 223398 532768 223634
rect 532448 223366 532768 223398
rect 563168 223954 563488 223986
rect 563168 223718 563210 223954
rect 563446 223718 563488 223954
rect 563168 223634 563488 223718
rect 563168 223398 563210 223634
rect 563446 223398 563488 223634
rect 563168 223366 563488 223398
rect 394208 219454 394528 219486
rect 394208 219218 394250 219454
rect 394486 219218 394528 219454
rect 394208 219134 394528 219218
rect 394208 218898 394250 219134
rect 394486 218898 394528 219134
rect 394208 218866 394528 218898
rect 424928 219454 425248 219486
rect 424928 219218 424970 219454
rect 425206 219218 425248 219454
rect 424928 219134 425248 219218
rect 424928 218898 424970 219134
rect 425206 218898 425248 219134
rect 424928 218866 425248 218898
rect 455648 219454 455968 219486
rect 455648 219218 455690 219454
rect 455926 219218 455968 219454
rect 455648 219134 455968 219218
rect 455648 218898 455690 219134
rect 455926 218898 455968 219134
rect 455648 218866 455968 218898
rect 486368 219454 486688 219486
rect 486368 219218 486410 219454
rect 486646 219218 486688 219454
rect 486368 219134 486688 219218
rect 486368 218898 486410 219134
rect 486646 218898 486688 219134
rect 486368 218866 486688 218898
rect 517088 219454 517408 219486
rect 517088 219218 517130 219454
rect 517366 219218 517408 219454
rect 517088 219134 517408 219218
rect 517088 218898 517130 219134
rect 517366 218898 517408 219134
rect 517088 218866 517408 218898
rect 547808 219454 548128 219486
rect 547808 219218 547850 219454
rect 548086 219218 548128 219454
rect 547808 219134 548128 219218
rect 547808 218898 547850 219134
rect 548086 218898 548128 219134
rect 547808 218866 548128 218898
rect 388483 213892 388549 213893
rect 388483 213828 388484 213892
rect 388548 213828 388549 213892
rect 388483 213827 388549 213828
rect 409568 187954 409888 187986
rect 409568 187718 409610 187954
rect 409846 187718 409888 187954
rect 409568 187634 409888 187718
rect 409568 187398 409610 187634
rect 409846 187398 409888 187634
rect 409568 187366 409888 187398
rect 440288 187954 440608 187986
rect 440288 187718 440330 187954
rect 440566 187718 440608 187954
rect 440288 187634 440608 187718
rect 440288 187398 440330 187634
rect 440566 187398 440608 187634
rect 440288 187366 440608 187398
rect 471008 187954 471328 187986
rect 471008 187718 471050 187954
rect 471286 187718 471328 187954
rect 471008 187634 471328 187718
rect 471008 187398 471050 187634
rect 471286 187398 471328 187634
rect 471008 187366 471328 187398
rect 501728 187954 502048 187986
rect 501728 187718 501770 187954
rect 502006 187718 502048 187954
rect 501728 187634 502048 187718
rect 501728 187398 501770 187634
rect 502006 187398 502048 187634
rect 501728 187366 502048 187398
rect 532448 187954 532768 187986
rect 532448 187718 532490 187954
rect 532726 187718 532768 187954
rect 532448 187634 532768 187718
rect 532448 187398 532490 187634
rect 532726 187398 532768 187634
rect 532448 187366 532768 187398
rect 563168 187954 563488 187986
rect 563168 187718 563210 187954
rect 563446 187718 563488 187954
rect 563168 187634 563488 187718
rect 563168 187398 563210 187634
rect 563446 187398 563488 187634
rect 563168 187366 563488 187398
rect 394208 183454 394528 183486
rect 394208 183218 394250 183454
rect 394486 183218 394528 183454
rect 394208 183134 394528 183218
rect 394208 182898 394250 183134
rect 394486 182898 394528 183134
rect 394208 182866 394528 182898
rect 424928 183454 425248 183486
rect 424928 183218 424970 183454
rect 425206 183218 425248 183454
rect 424928 183134 425248 183218
rect 424928 182898 424970 183134
rect 425206 182898 425248 183134
rect 424928 182866 425248 182898
rect 455648 183454 455968 183486
rect 455648 183218 455690 183454
rect 455926 183218 455968 183454
rect 455648 183134 455968 183218
rect 455648 182898 455690 183134
rect 455926 182898 455968 183134
rect 455648 182866 455968 182898
rect 486368 183454 486688 183486
rect 486368 183218 486410 183454
rect 486646 183218 486688 183454
rect 486368 183134 486688 183218
rect 486368 182898 486410 183134
rect 486646 182898 486688 183134
rect 486368 182866 486688 182898
rect 517088 183454 517408 183486
rect 517088 183218 517130 183454
rect 517366 183218 517408 183454
rect 517088 183134 517408 183218
rect 517088 182898 517130 183134
rect 517366 182898 517408 183134
rect 517088 182866 517408 182898
rect 547808 183454 548128 183486
rect 547808 183218 547850 183454
rect 548086 183218 548128 183454
rect 547808 183134 548128 183218
rect 547808 182898 547850 183134
rect 548086 182898 548128 183134
rect 547808 182866 548128 182898
rect 569542 173909 569602 278699
rect 569539 173908 569605 173909
rect 569539 173844 569540 173908
rect 569604 173844 569605 173908
rect 569539 173843 569605 173844
rect 409568 151954 409888 151986
rect 409568 151718 409610 151954
rect 409846 151718 409888 151954
rect 409568 151634 409888 151718
rect 409568 151398 409610 151634
rect 409846 151398 409888 151634
rect 409568 151366 409888 151398
rect 440288 151954 440608 151986
rect 440288 151718 440330 151954
rect 440566 151718 440608 151954
rect 440288 151634 440608 151718
rect 440288 151398 440330 151634
rect 440566 151398 440608 151634
rect 440288 151366 440608 151398
rect 471008 151954 471328 151986
rect 471008 151718 471050 151954
rect 471286 151718 471328 151954
rect 471008 151634 471328 151718
rect 471008 151398 471050 151634
rect 471286 151398 471328 151634
rect 471008 151366 471328 151398
rect 501728 151954 502048 151986
rect 501728 151718 501770 151954
rect 502006 151718 502048 151954
rect 501728 151634 502048 151718
rect 501728 151398 501770 151634
rect 502006 151398 502048 151634
rect 501728 151366 502048 151398
rect 532448 151954 532768 151986
rect 532448 151718 532490 151954
rect 532726 151718 532768 151954
rect 532448 151634 532768 151718
rect 532448 151398 532490 151634
rect 532726 151398 532768 151634
rect 532448 151366 532768 151398
rect 563168 151954 563488 151986
rect 563168 151718 563210 151954
rect 563446 151718 563488 151954
rect 563168 151634 563488 151718
rect 563168 151398 563210 151634
rect 563446 151398 563488 151634
rect 563168 151366 563488 151398
rect 394208 147454 394528 147486
rect 394208 147218 394250 147454
rect 394486 147218 394528 147454
rect 394208 147134 394528 147218
rect 394208 146898 394250 147134
rect 394486 146898 394528 147134
rect 394208 146866 394528 146898
rect 424928 147454 425248 147486
rect 424928 147218 424970 147454
rect 425206 147218 425248 147454
rect 424928 147134 425248 147218
rect 424928 146898 424970 147134
rect 425206 146898 425248 147134
rect 424928 146866 425248 146898
rect 455648 147454 455968 147486
rect 455648 147218 455690 147454
rect 455926 147218 455968 147454
rect 455648 147134 455968 147218
rect 455648 146898 455690 147134
rect 455926 146898 455968 147134
rect 455648 146866 455968 146898
rect 486368 147454 486688 147486
rect 486368 147218 486410 147454
rect 486646 147218 486688 147454
rect 486368 147134 486688 147218
rect 486368 146898 486410 147134
rect 486646 146898 486688 147134
rect 486368 146866 486688 146898
rect 517088 147454 517408 147486
rect 517088 147218 517130 147454
rect 517366 147218 517408 147454
rect 517088 147134 517408 147218
rect 517088 146898 517130 147134
rect 517366 146898 517408 147134
rect 517088 146866 517408 146898
rect 547808 147454 548128 147486
rect 547808 147218 547850 147454
rect 548086 147218 548128 147454
rect 547808 147134 548128 147218
rect 547808 146898 547850 147134
rect 548086 146898 548128 147134
rect 547808 146866 548128 146898
rect 409568 115954 409888 115986
rect 409568 115718 409610 115954
rect 409846 115718 409888 115954
rect 409568 115634 409888 115718
rect 409568 115398 409610 115634
rect 409846 115398 409888 115634
rect 409568 115366 409888 115398
rect 440288 115954 440608 115986
rect 440288 115718 440330 115954
rect 440566 115718 440608 115954
rect 440288 115634 440608 115718
rect 440288 115398 440330 115634
rect 440566 115398 440608 115634
rect 440288 115366 440608 115398
rect 471008 115954 471328 115986
rect 471008 115718 471050 115954
rect 471286 115718 471328 115954
rect 471008 115634 471328 115718
rect 471008 115398 471050 115634
rect 471286 115398 471328 115634
rect 471008 115366 471328 115398
rect 501728 115954 502048 115986
rect 501728 115718 501770 115954
rect 502006 115718 502048 115954
rect 501728 115634 502048 115718
rect 501728 115398 501770 115634
rect 502006 115398 502048 115634
rect 501728 115366 502048 115398
rect 532448 115954 532768 115986
rect 532448 115718 532490 115954
rect 532726 115718 532768 115954
rect 532448 115634 532768 115718
rect 532448 115398 532490 115634
rect 532726 115398 532768 115634
rect 532448 115366 532768 115398
rect 563168 115954 563488 115986
rect 563168 115718 563210 115954
rect 563446 115718 563488 115954
rect 563168 115634 563488 115718
rect 563168 115398 563210 115634
rect 563446 115398 563488 115634
rect 563168 115366 563488 115398
rect 389771 115156 389837 115157
rect 389771 115092 389772 115156
rect 389836 115092 389837 115156
rect 389771 115091 389837 115092
rect 389774 96253 389834 115091
rect 394208 111454 394528 111486
rect 394208 111218 394250 111454
rect 394486 111218 394528 111454
rect 394208 111134 394528 111218
rect 394208 110898 394250 111134
rect 394486 110898 394528 111134
rect 394208 110866 394528 110898
rect 424928 111454 425248 111486
rect 424928 111218 424970 111454
rect 425206 111218 425248 111454
rect 424928 111134 425248 111218
rect 424928 110898 424970 111134
rect 425206 110898 425248 111134
rect 424928 110866 425248 110898
rect 455648 111454 455968 111486
rect 455648 111218 455690 111454
rect 455926 111218 455968 111454
rect 455648 111134 455968 111218
rect 455648 110898 455690 111134
rect 455926 110898 455968 111134
rect 455648 110866 455968 110898
rect 486368 111454 486688 111486
rect 486368 111218 486410 111454
rect 486646 111218 486688 111454
rect 486368 111134 486688 111218
rect 486368 110898 486410 111134
rect 486646 110898 486688 111134
rect 486368 110866 486688 110898
rect 517088 111454 517408 111486
rect 517088 111218 517130 111454
rect 517366 111218 517408 111454
rect 517088 111134 517408 111218
rect 517088 110898 517130 111134
rect 517366 110898 517408 111134
rect 517088 110866 517408 110898
rect 547808 111454 548128 111486
rect 547808 111218 547850 111454
rect 548086 111218 548128 111454
rect 547808 111134 548128 111218
rect 547808 110898 547850 111134
rect 548086 110898 548128 111134
rect 547808 110866 548128 110898
rect 570094 109717 570154 364379
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 579659 511324 579725 511325
rect 579659 511260 579660 511324
rect 579724 511260 579725 511324
rect 579659 511259 579725 511260
rect 579662 510645 579722 511259
rect 579659 510644 579725 510645
rect 579659 510580 579660 510644
rect 579724 510580 579725 510644
rect 579659 510579 579725 510580
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 574691 294540 574757 294541
rect 574691 294476 574692 294540
rect 574756 294476 574757 294540
rect 574691 294475 574757 294476
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 571563 284884 571629 284885
rect 571563 284820 571564 284884
rect 571628 284820 571629 284884
rect 571563 284819 571629 284820
rect 571379 244356 571445 244357
rect 571379 244292 571380 244356
rect 571444 244292 571445 244356
rect 571379 244291 571445 244292
rect 570091 109716 570157 109717
rect 570091 109652 570092 109716
rect 570156 109652 570157 109716
rect 570091 109651 570157 109652
rect 389771 96252 389837 96253
rect 389771 96188 389772 96252
rect 389836 96188 389837 96252
rect 389771 96187 389837 96188
rect 388794 66454 389414 94000
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388299 19412 388365 19413
rect 388299 19348 388300 19412
rect 388364 19348 388365 19412
rect 388299 19347 388365 19348
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 70954 393914 94000
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 75454 398414 94000
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 79954 402914 94000
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 84454 407414 94000
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 88954 411914 94000
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 93454 416414 94000
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 61954 420914 94000
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 66454 425414 94000
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 70954 429914 94000
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 75454 434414 94000
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 79954 438914 94000
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 84454 443414 94000
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 88954 447914 94000
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 93454 452414 94000
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 61954 456914 94000
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 66454 461414 94000
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 70954 465914 94000
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 75454 470414 94000
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 79954 474914 94000
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 84454 479414 94000
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 88954 483914 94000
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 93454 488414 94000
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 61954 492914 94000
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 66454 497414 94000
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 70954 501914 94000
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 75454 506414 94000
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 79954 510914 94000
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 84454 515414 94000
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 88954 519914 94000
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 93454 524414 94000
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 61954 528914 94000
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 66454 533414 94000
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 70954 537914 94000
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 75454 542414 94000
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 79954 546914 94000
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 84454 551414 94000
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 88954 555914 94000
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 93454 560414 94000
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 61954 564914 94000
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 66454 569414 94000
rect 571382 84149 571442 244291
rect 571566 200837 571626 284819
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 571563 200836 571629 200837
rect 571563 200772 571564 200836
rect 571628 200772 571629 200836
rect 571563 200771 571629 200772
rect 571563 193900 571629 193901
rect 571563 193836 571564 193900
rect 571628 193836 571629 193900
rect 571563 193835 571629 193836
rect 571566 96389 571626 193835
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 571563 96388 571629 96389
rect 571563 96324 571564 96388
rect 571628 96324 571629 96388
rect 571563 96323 571629 96324
rect 571379 84148 571445 84149
rect 571379 84084 571380 84148
rect 571444 84084 571445 84148
rect 571379 84083 571445 84084
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 70954 573914 106398
rect 574694 93669 574754 294475
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 574691 93668 574757 93669
rect 574691 93604 574692 93668
rect 574756 93604 574757 93668
rect 574691 93603 574757 93604
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 75454 578414 110898
rect 579662 97205 579722 510579
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 579659 97204 579725 97205
rect 579659 97140 579660 97204
rect 579724 97140 579725 97204
rect 579659 97139 579725 97140
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< obsm4 >>
rect 68800 174494 96960 174600
rect 97020 174494 98320 174600
rect 98380 174494 99408 174600
rect 99468 174494 100768 174600
rect 100828 174494 101992 174600
rect 102052 174494 103352 174600
rect 103412 174494 104576 174600
rect 104636 174494 105664 174600
rect 105724 174494 107024 174600
rect 107084 174494 108112 174600
rect 108172 174494 109472 174600
rect 109532 174494 110696 174600
rect 110756 174494 112056 174600
rect 112116 174494 113144 174600
rect 113204 174494 114368 174600
rect 114428 174494 115728 174600
rect 115788 174494 116952 174600
rect 117012 174494 118312 174600
rect 118372 174494 119400 174600
rect 119460 174494 120760 174600
rect 120820 174494 121848 174600
rect 121908 174494 123072 174600
rect 123132 174494 124432 174600
rect 124492 174494 125656 174600
rect 125716 174494 127016 174600
rect 127076 174494 128104 174600
rect 128164 174494 129464 174600
rect 129524 174494 130688 174600
rect 130748 174494 132048 174600
rect 132108 174494 133136 174600
rect 133196 174494 134360 174600
rect 134420 174494 135720 174600
rect 135780 174494 148232 174600
rect 148292 174494 158840 174600
rect 158900 174494 164756 174600
rect 68800 151986 164756 174494
rect 68800 151366 69072 151986
rect 69420 151366 164136 151986
rect 164484 151366 164756 151986
rect 68800 147486 164756 151366
rect 68800 146866 69752 147486
rect 70100 146866 163456 147486
rect 163804 146866 164756 147486
rect 68800 115986 164756 146866
rect 68800 115366 69072 115986
rect 69420 115366 164136 115986
rect 164484 115366 164756 115986
rect 68800 111486 164756 115366
rect 68800 110866 69752 111486
rect 70100 110866 163456 111486
rect 163804 110866 164756 111486
rect 68800 95200 164756 110866
rect 68800 95100 74656 95200
rect 74716 95100 84312 95200
rect 84372 95100 85536 95200
rect 85596 95100 86624 95200
rect 86684 95100 87984 95200
rect 88044 95100 88936 95200
rect 88996 95100 90160 95200
rect 90220 95100 91384 95200
rect 91444 95100 92472 95200
rect 92532 95100 93832 95200
rect 93892 95100 94920 95200
rect 94980 95100 96008 95200
rect 96068 95100 96688 95200
rect 96748 95100 97096 95200
rect 97156 95100 98048 95200
rect 98108 95100 98456 95200
rect 98516 95100 99136 95200
rect 99196 95100 99544 95200
rect 99604 95100 100632 95200
rect 100692 95100 100768 95200
rect 100828 95100 101856 95200
rect 101916 95100 101992 95200
rect 102052 95100 102944 95200
rect 103004 95100 103216 95200
rect 103276 95100 104304 95200
rect 104364 95100 104440 95200
rect 104500 95100 105392 95200
rect 105452 95100 105664 95200
rect 105724 95100 106480 95200
rect 106540 95100 106616 95200
rect 106676 95100 107704 95200
rect 107764 95100 108112 95200
rect 108172 95100 109064 95200
rect 109124 95100 109472 95200
rect 109532 95100 110152 95200
rect 110212 95100 110696 95200
rect 110756 95100 111240 95200
rect 111300 95100 111920 95200
rect 111980 95100 112328 95200
rect 112388 95100 113144 95200
rect 113204 95100 113688 95200
rect 113748 95100 114368 95200
rect 114428 95100 114776 95200
rect 114836 95100 115456 95200
rect 115516 95100 115864 95200
rect 115924 95100 116680 95200
rect 116740 95100 117088 95200
rect 117148 95100 117904 95200
rect 117964 95100 118176 95200
rect 118236 95100 119400 95200
rect 119460 95100 119536 95200
rect 119596 95100 120216 95200
rect 120276 95100 120624 95200
rect 120684 95100 121712 95200
rect 121772 95100 121984 95200
rect 122044 95100 122800 95200
rect 122860 95100 123208 95200
rect 123268 95100 124024 95200
rect 124084 95100 124432 95200
rect 124492 95100 125384 95200
rect 125444 95100 125656 95200
rect 125716 95100 126472 95200
rect 126532 95100 126608 95200
rect 126668 95100 128104 95200
rect 128164 95100 129328 95200
rect 129388 95100 130688 95200
rect 130748 95100 131912 95200
rect 131972 95100 133136 95200
rect 133196 95100 134360 95200
rect 134420 95100 135584 95200
rect 135644 95100 151496 95200
rect 151556 95100 151632 95200
rect 151692 95100 151768 95200
rect 151828 95100 151904 95200
rect 151964 95100 164756 95200
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 89610 259718 89846 259954
rect 89610 259398 89846 259634
rect 74250 255218 74486 255454
rect 74250 254898 74486 255134
rect 104970 255218 105206 255454
rect 104970 254898 105206 255134
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 118826 228218 119062 228454
rect 119146 228218 119382 228454
rect 118826 227898 119062 228134
rect 119146 227898 119382 228134
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 123326 232718 123562 232954
rect 123646 232718 123882 232954
rect 123326 232398 123562 232634
rect 123646 232398 123882 232634
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 132326 241718 132562 241954
rect 132646 241718 132882 241954
rect 132326 241398 132562 241634
rect 132646 241398 132882 241634
rect 132326 205718 132562 205954
rect 132646 205718 132882 205954
rect 132326 205398 132562 205634
rect 132646 205398 132882 205634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 136826 246218 137062 246454
rect 137146 246218 137382 246454
rect 136826 245898 137062 246134
rect 137146 245898 137382 246134
rect 136826 210218 137062 210454
rect 137146 210218 137382 210454
rect 136826 209898 137062 210134
rect 137146 209898 137382 210134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 141326 214718 141562 214954
rect 141646 214718 141882 214954
rect 141326 214398 141562 214634
rect 141646 214398 141882 214634
rect 141326 178718 141562 178954
rect 141646 178718 141882 178954
rect 141326 178398 141562 178634
rect 141646 178398 141882 178634
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 150326 223718 150562 223954
rect 150646 223718 150882 223954
rect 150326 223398 150562 223634
rect 150646 223398 150882 223634
rect 150326 187718 150562 187954
rect 150646 187718 150882 187954
rect 150326 187398 150562 187634
rect 150646 187398 150882 187634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 154826 228218 155062 228454
rect 155146 228218 155382 228454
rect 154826 227898 155062 228134
rect 155146 227898 155382 228134
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 159326 232718 159562 232954
rect 159646 232718 159882 232954
rect 159326 232398 159562 232634
rect 159646 232398 159882 232634
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 168326 241718 168562 241954
rect 168646 241718 168882 241954
rect 168326 241398 168562 241634
rect 168646 241398 168882 241634
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 168326 205718 168562 205954
rect 168646 205718 168882 205954
rect 168326 205398 168562 205634
rect 168646 205398 168882 205634
rect 69128 151718 69364 151954
rect 69128 151398 69364 151634
rect 164192 151718 164428 151954
rect 164192 151398 164428 151634
rect 69808 147218 70044 147454
rect 69808 146898 70044 147134
rect 163512 147218 163748 147454
rect 163512 146898 163748 147134
rect 69128 115718 69364 115954
rect 69128 115398 69364 115634
rect 164192 115718 164428 115954
rect 164192 115398 164428 115634
rect 69808 111218 70044 111454
rect 69808 110898 70044 111134
rect 163512 111218 163748 111454
rect 163512 110898 163748 111134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 84218 119062 84454
rect 119146 84218 119382 84454
rect 118826 83898 119062 84134
rect 119146 83898 119382 84134
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 88718 123562 88954
rect 123646 88718 123882 88954
rect 123326 88398 123562 88634
rect 123646 88398 123882 88634
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 79718 150562 79954
rect 150646 79718 150882 79954
rect 150326 79398 150562 79634
rect 150646 79398 150882 79634
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 154826 84218 155062 84454
rect 155146 84218 155382 84454
rect 154826 83898 155062 84134
rect 155146 83898 155382 84134
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 159326 88718 159562 88954
rect 159646 88718 159882 88954
rect 159326 88398 159562 88634
rect 159646 88398 159882 88634
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 168326 169718 168562 169954
rect 168646 169718 168882 169954
rect 168326 169398 168562 169634
rect 168646 169398 168882 169634
rect 168326 133718 168562 133954
rect 168646 133718 168882 133954
rect 168326 133398 168562 133634
rect 168646 133398 168882 133634
rect 168326 97718 168562 97954
rect 168646 97718 168882 97954
rect 168326 97398 168562 97634
rect 168646 97398 168882 97634
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 172826 246218 173062 246454
rect 173146 246218 173382 246454
rect 172826 245898 173062 246134
rect 173146 245898 173382 246134
rect 172826 210218 173062 210454
rect 173146 210218 173382 210454
rect 172826 209898 173062 210134
rect 173146 209898 173382 210134
rect 172826 174218 173062 174454
rect 173146 174218 173382 174454
rect 172826 173898 173062 174134
rect 173146 173898 173382 174134
rect 172826 138218 173062 138454
rect 173146 138218 173382 138454
rect 172826 137898 173062 138134
rect 173146 137898 173382 138134
rect 172826 102218 173062 102454
rect 173146 102218 173382 102454
rect 172826 101898 173062 102134
rect 173146 101898 173382 102134
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 222326 547718 222562 547954
rect 222646 547718 222882 547954
rect 222326 547398 222562 547634
rect 222646 547398 222882 547634
rect 222326 511718 222562 511954
rect 222646 511718 222882 511954
rect 222326 511398 222562 511634
rect 222646 511398 222882 511634
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 226826 552218 227062 552454
rect 227146 552218 227382 552454
rect 226826 551898 227062 552134
rect 227146 551898 227382 552134
rect 226826 516218 227062 516454
rect 227146 516218 227382 516454
rect 226826 515898 227062 516134
rect 227146 515898 227382 516134
rect 226826 480218 227062 480454
rect 227146 480218 227382 480454
rect 226826 479898 227062 480134
rect 227146 479898 227382 480134
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 231326 556718 231562 556954
rect 231646 556718 231882 556954
rect 231326 556398 231562 556634
rect 231646 556398 231882 556634
rect 231326 520718 231562 520954
rect 231646 520718 231882 520954
rect 231326 520398 231562 520634
rect 231646 520398 231882 520634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 231326 412718 231562 412954
rect 231646 412718 231882 412954
rect 231326 412398 231562 412634
rect 231646 412398 231882 412634
rect 231326 376718 231562 376954
rect 231646 376718 231882 376954
rect 231326 376398 231562 376634
rect 231646 376398 231882 376634
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 240326 529718 240562 529954
rect 240646 529718 240882 529954
rect 240326 529398 240562 529634
rect 240646 529398 240882 529634
rect 240326 493718 240562 493954
rect 240646 493718 240882 493954
rect 240326 493398 240562 493634
rect 240646 493398 240882 493634
rect 240326 457718 240562 457954
rect 240646 457718 240882 457954
rect 240326 457398 240562 457634
rect 240646 457398 240882 457634
rect 240326 421718 240562 421954
rect 240646 421718 240882 421954
rect 240326 421398 240562 421634
rect 240646 421398 240882 421634
rect 240326 385718 240562 385954
rect 240646 385718 240882 385954
rect 240326 385398 240562 385634
rect 240646 385398 240882 385634
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 244826 534218 245062 534454
rect 245146 534218 245382 534454
rect 244826 533898 245062 534134
rect 245146 533898 245382 534134
rect 244826 498218 245062 498454
rect 245146 498218 245382 498454
rect 244826 497898 245062 498134
rect 245146 497898 245382 498134
rect 244826 462218 245062 462454
rect 245146 462218 245382 462454
rect 244826 461898 245062 462134
rect 245146 461898 245382 462134
rect 244826 426218 245062 426454
rect 245146 426218 245382 426454
rect 244826 425898 245062 426134
rect 245146 425898 245382 426134
rect 244826 390218 245062 390454
rect 245146 390218 245382 390454
rect 244826 389898 245062 390134
rect 245146 389898 245382 390134
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 249326 538718 249562 538954
rect 249646 538718 249882 538954
rect 249326 538398 249562 538634
rect 249646 538398 249882 538634
rect 249326 502718 249562 502954
rect 249646 502718 249882 502954
rect 249326 502398 249562 502634
rect 249646 502398 249882 502634
rect 249326 466718 249562 466954
rect 249646 466718 249882 466954
rect 249326 466398 249562 466634
rect 249646 466398 249882 466634
rect 249326 430718 249562 430954
rect 249646 430718 249882 430954
rect 249326 430398 249562 430634
rect 249646 430398 249882 430634
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 249326 358718 249562 358954
rect 249646 358718 249882 358954
rect 249326 358398 249562 358634
rect 249646 358398 249882 358634
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 276326 529718 276562 529954
rect 276646 529718 276882 529954
rect 276326 529398 276562 529634
rect 276646 529398 276882 529634
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 280826 534218 281062 534454
rect 281146 534218 281382 534454
rect 280826 533898 281062 534134
rect 281146 533898 281382 534134
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 177326 214718 177562 214954
rect 177646 214718 177882 214954
rect 177326 214398 177562 214634
rect 177646 214398 177882 214634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 177326 106718 177562 106954
rect 177646 106718 177882 106954
rect 177326 106398 177562 106634
rect 177646 106398 177882 106634
rect 199610 331718 199846 331954
rect 199610 331398 199846 331634
rect 230330 331718 230566 331954
rect 230330 331398 230566 331634
rect 261050 331718 261286 331954
rect 261050 331398 261286 331634
rect 184250 327218 184486 327454
rect 184250 326898 184486 327134
rect 214970 327218 215206 327454
rect 214970 326898 215206 327134
rect 245690 327218 245926 327454
rect 245690 326898 245926 327134
rect 276410 327218 276646 327454
rect 276410 326898 276646 327134
rect 199610 295718 199846 295954
rect 199610 295398 199846 295634
rect 230330 295718 230566 295954
rect 230330 295398 230566 295634
rect 261050 295718 261286 295954
rect 261050 295398 261286 295634
rect 184250 291218 184486 291454
rect 184250 290898 184486 291134
rect 214970 291218 215206 291454
rect 214970 290898 215206 291134
rect 245690 291218 245926 291454
rect 245690 290898 245926 291134
rect 276410 291218 276646 291454
rect 276410 290898 276646 291134
rect 199610 259718 199846 259954
rect 199610 259398 199846 259634
rect 230330 259718 230566 259954
rect 230330 259398 230566 259634
rect 261050 259718 261286 259954
rect 261050 259398 261286 259634
rect 184250 255218 184486 255454
rect 184250 254898 184486 255134
rect 214970 255218 215206 255454
rect 214970 254898 215206 255134
rect 245690 255218 245926 255454
rect 245690 254898 245926 255134
rect 276410 255218 276646 255454
rect 276410 254898 276646 255134
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 186326 115718 186562 115954
rect 186646 115718 186882 115954
rect 186326 115398 186562 115634
rect 186646 115398 186882 115634
rect 186326 79718 186562 79954
rect 186646 79718 186882 79954
rect 186326 79398 186562 79634
rect 186646 79398 186882 79634
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 228218 191062 228454
rect 191146 228218 191382 228454
rect 190826 227898 191062 228134
rect 191146 227898 191382 228134
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 190826 120218 191062 120454
rect 191146 120218 191382 120454
rect 190826 119898 191062 120134
rect 191146 119898 191382 120134
rect 190826 84218 191062 84454
rect 191146 84218 191382 84454
rect 190826 83898 191062 84134
rect 191146 83898 191382 84134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 232718 195562 232954
rect 195646 232718 195882 232954
rect 195326 232398 195562 232634
rect 195646 232398 195882 232634
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 226826 228218 227062 228454
rect 227146 228218 227382 228454
rect 226826 227898 227062 228134
rect 227146 227898 227382 228134
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 231326 232718 231562 232954
rect 231646 232718 231882 232954
rect 231326 232398 231562 232634
rect 231646 232398 231882 232634
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 227916 151718 228152 151954
rect 227916 151398 228152 151634
rect 237847 151718 238083 151954
rect 237847 151398 238083 151634
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 222952 147218 223188 147454
rect 222952 146898 223188 147134
rect 232882 147218 233118 147454
rect 232882 146898 233118 147134
rect 242813 147218 243049 147454
rect 242813 146898 243049 147134
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 227916 115718 228152 115954
rect 227916 115398 228152 115634
rect 237847 115718 238083 115954
rect 237847 115398 238083 115634
rect 222952 111218 223188 111454
rect 222952 110898 223188 111134
rect 232882 111218 233118 111454
rect 232882 110898 233118 111134
rect 242813 111218 243049 111454
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 242813 110898 243049 111134
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 262826 228218 263062 228454
rect 263146 228218 263382 228454
rect 262826 227898 263062 228134
rect 263146 227898 263382 228134
rect 267326 232718 267562 232954
rect 267646 232718 267882 232954
rect 267326 232398 267562 232634
rect 267646 232398 267882 232634
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 298826 516218 299062 516454
rect 299146 516218 299382 516454
rect 298826 515898 299062 516134
rect 299146 515898 299382 516134
rect 298826 480218 299062 480454
rect 299146 480218 299382 480454
rect 298826 479898 299062 480134
rect 299146 479898 299382 480134
rect 298826 444218 299062 444454
rect 299146 444218 299382 444454
rect 298826 443898 299062 444134
rect 299146 443898 299382 444134
rect 298826 408218 299062 408454
rect 299146 408218 299382 408454
rect 298826 407898 299062 408134
rect 299146 407898 299382 408134
rect 298826 372218 299062 372454
rect 299146 372218 299382 372454
rect 298826 371898 299062 372134
rect 299146 371898 299382 372134
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 298826 228218 299062 228454
rect 299146 228218 299382 228454
rect 298826 227898 299062 228134
rect 299146 227898 299382 228134
rect 298826 192218 299062 192454
rect 299146 192218 299382 192454
rect 298826 191898 299062 192134
rect 299146 191898 299382 192134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 303326 556718 303562 556954
rect 303646 556718 303882 556954
rect 303326 556398 303562 556634
rect 303646 556398 303882 556634
rect 303326 520718 303562 520954
rect 303646 520718 303882 520954
rect 303326 520398 303562 520634
rect 303646 520398 303882 520634
rect 303326 484718 303562 484954
rect 303646 484718 303882 484954
rect 303326 484398 303562 484634
rect 303646 484398 303882 484634
rect 303326 448718 303562 448954
rect 303646 448718 303882 448954
rect 303326 448398 303562 448634
rect 303646 448398 303882 448634
rect 303326 412718 303562 412954
rect 303646 412718 303882 412954
rect 303326 412398 303562 412634
rect 303646 412398 303882 412634
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 303326 232718 303562 232954
rect 303646 232718 303882 232954
rect 303326 232398 303562 232634
rect 303646 232398 303882 232634
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 312326 529718 312562 529954
rect 312646 529718 312882 529954
rect 312326 529398 312562 529634
rect 312646 529398 312882 529634
rect 312326 493718 312562 493954
rect 312646 493718 312882 493954
rect 312326 493398 312562 493634
rect 312646 493398 312882 493634
rect 312326 457718 312562 457954
rect 312646 457718 312882 457954
rect 312326 457398 312562 457634
rect 312646 457398 312882 457634
rect 312326 421718 312562 421954
rect 312646 421718 312882 421954
rect 312326 421398 312562 421634
rect 312646 421398 312882 421634
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 312326 313718 312562 313954
rect 312646 313718 312882 313954
rect 312326 313398 312562 313634
rect 312646 313398 312882 313634
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 312326 241718 312562 241954
rect 312646 241718 312882 241954
rect 312326 241398 312562 241634
rect 312646 241398 312882 241634
rect 312326 205718 312562 205954
rect 312646 205718 312882 205954
rect 312326 205398 312562 205634
rect 312646 205398 312882 205634
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 316826 534218 317062 534454
rect 317146 534218 317382 534454
rect 316826 533898 317062 534134
rect 317146 533898 317382 534134
rect 316826 498218 317062 498454
rect 317146 498218 317382 498454
rect 316826 497898 317062 498134
rect 317146 497898 317382 498134
rect 316826 462218 317062 462454
rect 317146 462218 317382 462454
rect 316826 461898 317062 462134
rect 317146 461898 317382 462134
rect 316826 426218 317062 426454
rect 317146 426218 317382 426454
rect 316826 425898 317062 426134
rect 317146 425898 317382 426134
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 316826 318218 317062 318454
rect 317146 318218 317382 318454
rect 316826 317898 317062 318134
rect 317146 317898 317382 318134
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 316826 246218 317062 246454
rect 317146 246218 317382 246454
rect 316826 245898 317062 246134
rect 317146 245898 317382 246134
rect 316826 210218 317062 210454
rect 317146 210218 317382 210454
rect 316826 209898 317062 210134
rect 317146 209898 317382 210134
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 321326 538718 321562 538954
rect 321646 538718 321882 538954
rect 321326 538398 321562 538634
rect 321646 538398 321882 538634
rect 321326 502718 321562 502954
rect 321646 502718 321882 502954
rect 321326 502398 321562 502634
rect 321646 502398 321882 502634
rect 321326 466718 321562 466954
rect 321646 466718 321882 466954
rect 321326 466398 321562 466634
rect 321646 466398 321882 466634
rect 321326 430718 321562 430954
rect 321646 430718 321882 430954
rect 321326 430398 321562 430634
rect 321646 430398 321882 430634
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 321326 322718 321562 322954
rect 321646 322718 321882 322954
rect 321326 322398 321562 322634
rect 321646 322398 321882 322634
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 321326 214718 321562 214954
rect 321646 214718 321882 214954
rect 321326 214398 321562 214634
rect 321646 214398 321882 214634
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 321326 178718 321562 178954
rect 321646 178718 321882 178954
rect 321326 178398 321562 178634
rect 321646 178398 321882 178634
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 314250 151718 314486 151954
rect 314250 151398 314486 151634
rect 317514 151718 317750 151954
rect 317514 151398 317750 151634
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 330326 511718 330562 511954
rect 330646 511718 330882 511954
rect 330326 511398 330562 511634
rect 330646 511398 330882 511634
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 330326 439718 330562 439954
rect 330646 439718 330882 439954
rect 330326 439398 330562 439634
rect 330646 439398 330882 439634
rect 330326 403718 330562 403954
rect 330646 403718 330882 403954
rect 330326 403398 330562 403634
rect 330646 403398 330882 403634
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 330326 223718 330562 223954
rect 330646 223718 330882 223954
rect 330326 223398 330562 223634
rect 330646 223398 330882 223634
rect 330326 187718 330562 187954
rect 330646 187718 330882 187954
rect 330326 187398 330562 187634
rect 330646 187398 330882 187634
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 312618 147218 312854 147454
rect 312618 146898 312854 147134
rect 315882 147218 316118 147454
rect 315882 146898 316118 147134
rect 319146 147218 319382 147454
rect 319146 146898 319382 147134
rect 314250 115718 314486 115954
rect 314250 115398 314486 115634
rect 317514 115718 317750 115954
rect 317514 115398 317750 115634
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 312618 111218 312854 111454
rect 312618 110898 312854 111134
rect 315882 111218 316118 111454
rect 315882 110898 316118 111134
rect 319146 111218 319382 111454
rect 319146 110898 319382 111134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 334826 516218 335062 516454
rect 335146 516218 335382 516454
rect 334826 515898 335062 516134
rect 335146 515898 335382 516134
rect 334826 480218 335062 480454
rect 335146 480218 335382 480454
rect 334826 479898 335062 480134
rect 335146 479898 335382 480134
rect 334826 444218 335062 444454
rect 335146 444218 335382 444454
rect 334826 443898 335062 444134
rect 335146 443898 335382 444134
rect 334826 408218 335062 408454
rect 335146 408218 335382 408454
rect 334826 407898 335062 408134
rect 335146 407898 335382 408134
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 339326 556718 339562 556954
rect 339646 556718 339882 556954
rect 339326 556398 339562 556634
rect 339646 556398 339882 556634
rect 339326 520718 339562 520954
rect 339646 520718 339882 520954
rect 339326 520398 339562 520634
rect 339646 520398 339882 520634
rect 339326 484718 339562 484954
rect 339646 484718 339882 484954
rect 339326 484398 339562 484634
rect 339646 484398 339882 484634
rect 339326 448718 339562 448954
rect 339646 448718 339882 448954
rect 339326 448398 339562 448634
rect 339646 448398 339882 448634
rect 339326 412718 339562 412954
rect 339646 412718 339882 412954
rect 339326 412398 339562 412634
rect 339646 412398 339882 412634
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 334826 228218 335062 228454
rect 335146 228218 335382 228454
rect 334826 227898 335062 228134
rect 335146 227898 335382 228134
rect 334826 192218 335062 192454
rect 335146 192218 335382 192454
rect 334826 191898 335062 192134
rect 335146 191898 335382 192134
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 339326 232718 339562 232954
rect 339646 232718 339882 232954
rect 339326 232398 339562 232634
rect 339646 232398 339882 232634
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 348326 529718 348562 529954
rect 348646 529718 348882 529954
rect 348326 529398 348562 529634
rect 348646 529398 348882 529634
rect 348326 493718 348562 493954
rect 348646 493718 348882 493954
rect 348326 493398 348562 493634
rect 348646 493398 348882 493634
rect 348326 457718 348562 457954
rect 348646 457718 348882 457954
rect 348326 457398 348562 457634
rect 348646 457398 348882 457634
rect 348326 421718 348562 421954
rect 348646 421718 348882 421954
rect 348326 421398 348562 421634
rect 348646 421398 348882 421634
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 348326 313718 348562 313954
rect 348646 313718 348882 313954
rect 348326 313398 348562 313634
rect 348646 313398 348882 313634
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 348326 241718 348562 241954
rect 348646 241718 348882 241954
rect 348326 241398 348562 241634
rect 348646 241398 348882 241634
rect 348326 205718 348562 205954
rect 348646 205718 348882 205954
rect 348326 205398 348562 205634
rect 348646 205398 348882 205634
rect 348326 169718 348562 169954
rect 348646 169718 348882 169954
rect 348326 169398 348562 169634
rect 348646 169398 348882 169634
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 352826 426218 353062 426454
rect 353146 426218 353382 426454
rect 352826 425898 353062 426134
rect 353146 425898 353382 426134
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 357326 538718 357562 538954
rect 357646 538718 357882 538954
rect 357326 538398 357562 538634
rect 357646 538398 357882 538634
rect 357326 502718 357562 502954
rect 357646 502718 357882 502954
rect 357326 502398 357562 502634
rect 357646 502398 357882 502634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 384326 241718 384562 241954
rect 384646 241718 384882 241954
rect 384326 241398 384562 241634
rect 384646 241398 384882 241634
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 409610 259718 409846 259954
rect 409610 259398 409846 259634
rect 440330 259718 440566 259954
rect 440330 259398 440566 259634
rect 471050 259718 471286 259954
rect 471050 259398 471286 259634
rect 501770 259718 502006 259954
rect 501770 259398 502006 259634
rect 532490 259718 532726 259954
rect 532490 259398 532726 259634
rect 563210 259718 563446 259954
rect 563210 259398 563446 259634
rect 394250 255218 394486 255454
rect 394250 254898 394486 255134
rect 424970 255218 425206 255454
rect 424970 254898 425206 255134
rect 455690 255218 455926 255454
rect 455690 254898 455926 255134
rect 486410 255218 486646 255454
rect 486410 254898 486646 255134
rect 517130 255218 517366 255454
rect 517130 254898 517366 255134
rect 547850 255218 548086 255454
rect 547850 254898 548086 255134
rect 409610 223718 409846 223954
rect 409610 223398 409846 223634
rect 440330 223718 440566 223954
rect 440330 223398 440566 223634
rect 471050 223718 471286 223954
rect 471050 223398 471286 223634
rect 501770 223718 502006 223954
rect 501770 223398 502006 223634
rect 532490 223718 532726 223954
rect 532490 223398 532726 223634
rect 563210 223718 563446 223954
rect 563210 223398 563446 223634
rect 394250 219218 394486 219454
rect 394250 218898 394486 219134
rect 424970 219218 425206 219454
rect 424970 218898 425206 219134
rect 455690 219218 455926 219454
rect 455690 218898 455926 219134
rect 486410 219218 486646 219454
rect 486410 218898 486646 219134
rect 517130 219218 517366 219454
rect 517130 218898 517366 219134
rect 547850 219218 548086 219454
rect 547850 218898 548086 219134
rect 409610 187718 409846 187954
rect 409610 187398 409846 187634
rect 440330 187718 440566 187954
rect 440330 187398 440566 187634
rect 471050 187718 471286 187954
rect 471050 187398 471286 187634
rect 501770 187718 502006 187954
rect 501770 187398 502006 187634
rect 532490 187718 532726 187954
rect 532490 187398 532726 187634
rect 563210 187718 563446 187954
rect 563210 187398 563446 187634
rect 394250 183218 394486 183454
rect 394250 182898 394486 183134
rect 424970 183218 425206 183454
rect 424970 182898 425206 183134
rect 455690 183218 455926 183454
rect 455690 182898 455926 183134
rect 486410 183218 486646 183454
rect 486410 182898 486646 183134
rect 517130 183218 517366 183454
rect 517130 182898 517366 183134
rect 547850 183218 548086 183454
rect 547850 182898 548086 183134
rect 409610 151718 409846 151954
rect 409610 151398 409846 151634
rect 440330 151718 440566 151954
rect 440330 151398 440566 151634
rect 471050 151718 471286 151954
rect 471050 151398 471286 151634
rect 501770 151718 502006 151954
rect 501770 151398 502006 151634
rect 532490 151718 532726 151954
rect 532490 151398 532726 151634
rect 563210 151718 563446 151954
rect 563210 151398 563446 151634
rect 394250 147218 394486 147454
rect 394250 146898 394486 147134
rect 424970 147218 425206 147454
rect 424970 146898 425206 147134
rect 455690 147218 455926 147454
rect 455690 146898 455926 147134
rect 486410 147218 486646 147454
rect 486410 146898 486646 147134
rect 517130 147218 517366 147454
rect 517130 146898 517366 147134
rect 547850 147218 548086 147454
rect 547850 146898 548086 147134
rect 409610 115718 409846 115954
rect 409610 115398 409846 115634
rect 440330 115718 440566 115954
rect 440330 115398 440566 115634
rect 471050 115718 471286 115954
rect 471050 115398 471286 115634
rect 501770 115718 502006 115954
rect 501770 115398 502006 115634
rect 532490 115718 532726 115954
rect 532490 115398 532726 115634
rect 563210 115718 563446 115954
rect 563210 115398 563446 115634
rect 394250 111218 394486 111454
rect 394250 110898 394486 111134
rect 424970 111218 425206 111454
rect 424970 110898 425206 111134
rect 455690 111218 455926 111454
rect 455690 110898 455926 111134
rect 486410 111218 486646 111454
rect 486410 110898 486646 111134
rect 517130 111218 517366 111454
rect 517130 110898 517366 111134
rect 547850 111218 548086 111454
rect 547850 110898 548086 111134
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 199610 331954
rect 199846 331718 230330 331954
rect 230566 331718 261050 331954
rect 261286 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 199610 331634
rect 199846 331398 230330 331634
rect 230566 331398 261050 331634
rect 261286 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 184250 327454
rect 184486 327218 214970 327454
rect 215206 327218 245690 327454
rect 245926 327218 276410 327454
rect 276646 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 184250 327134
rect 184486 326898 214970 327134
rect 215206 326898 245690 327134
rect 245926 326898 276410 327134
rect 276646 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 199610 295954
rect 199846 295718 230330 295954
rect 230566 295718 261050 295954
rect 261286 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 199610 295634
rect 199846 295398 230330 295634
rect 230566 295398 261050 295634
rect 261286 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 184250 291454
rect 184486 291218 214970 291454
rect 215206 291218 245690 291454
rect 245926 291218 276410 291454
rect 276646 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 184250 291134
rect 184486 290898 214970 291134
rect 215206 290898 245690 291134
rect 245926 290898 276410 291134
rect 276646 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 89610 259954
rect 89846 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 199610 259954
rect 199846 259718 230330 259954
rect 230566 259718 261050 259954
rect 261286 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 409610 259954
rect 409846 259718 440330 259954
rect 440566 259718 471050 259954
rect 471286 259718 501770 259954
rect 502006 259718 532490 259954
rect 532726 259718 563210 259954
rect 563446 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 89610 259634
rect 89846 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 199610 259634
rect 199846 259398 230330 259634
rect 230566 259398 261050 259634
rect 261286 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 409610 259634
rect 409846 259398 440330 259634
rect 440566 259398 471050 259634
rect 471286 259398 501770 259634
rect 502006 259398 532490 259634
rect 532726 259398 563210 259634
rect 563446 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 74250 255454
rect 74486 255218 104970 255454
rect 105206 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 184250 255454
rect 184486 255218 214970 255454
rect 215206 255218 245690 255454
rect 245926 255218 276410 255454
rect 276646 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 394250 255454
rect 394486 255218 424970 255454
rect 425206 255218 455690 255454
rect 455926 255218 486410 255454
rect 486646 255218 517130 255454
rect 517366 255218 547850 255454
rect 548086 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 74250 255134
rect 74486 254898 104970 255134
rect 105206 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 184250 255134
rect 184486 254898 214970 255134
rect 215206 254898 245690 255134
rect 245926 254898 276410 255134
rect 276646 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 394250 255134
rect 394486 254898 424970 255134
rect 425206 254898 455690 255134
rect 455926 254898 486410 255134
rect 486646 254898 517130 255134
rect 517366 254898 547850 255134
rect 548086 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 409610 223954
rect 409846 223718 440330 223954
rect 440566 223718 471050 223954
rect 471286 223718 501770 223954
rect 502006 223718 532490 223954
rect 532726 223718 563210 223954
rect 563446 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 409610 223634
rect 409846 223398 440330 223634
rect 440566 223398 471050 223634
rect 471286 223398 501770 223634
rect 502006 223398 532490 223634
rect 532726 223398 563210 223634
rect 563446 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 394250 219454
rect 394486 219218 424970 219454
rect 425206 219218 455690 219454
rect 455926 219218 486410 219454
rect 486646 219218 517130 219454
rect 517366 219218 547850 219454
rect 548086 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 394250 219134
rect 394486 218898 424970 219134
rect 425206 218898 455690 219134
rect 455926 218898 486410 219134
rect 486646 218898 517130 219134
rect 517366 218898 547850 219134
rect 548086 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 409610 187954
rect 409846 187718 440330 187954
rect 440566 187718 471050 187954
rect 471286 187718 501770 187954
rect 502006 187718 532490 187954
rect 532726 187718 563210 187954
rect 563446 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 409610 187634
rect 409846 187398 440330 187634
rect 440566 187398 471050 187634
rect 471286 187398 501770 187634
rect 502006 187398 532490 187634
rect 532726 187398 563210 187634
rect 563446 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 394250 183454
rect 394486 183218 424970 183454
rect 425206 183218 455690 183454
rect 455926 183218 486410 183454
rect 486646 183218 517130 183454
rect 517366 183218 547850 183454
rect 548086 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 394250 183134
rect 394486 182898 424970 183134
rect 425206 182898 455690 183134
rect 455926 182898 486410 183134
rect 486646 182898 517130 183134
rect 517366 182898 547850 183134
rect 548086 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 69128 151954
rect 69364 151718 164192 151954
rect 164428 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 227916 151954
rect 228152 151718 237847 151954
rect 238083 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 314250 151954
rect 314486 151718 317514 151954
rect 317750 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 409610 151954
rect 409846 151718 440330 151954
rect 440566 151718 471050 151954
rect 471286 151718 501770 151954
rect 502006 151718 532490 151954
rect 532726 151718 563210 151954
rect 563446 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 69128 151634
rect 69364 151398 164192 151634
rect 164428 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 227916 151634
rect 228152 151398 237847 151634
rect 238083 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 314250 151634
rect 314486 151398 317514 151634
rect 317750 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 409610 151634
rect 409846 151398 440330 151634
rect 440566 151398 471050 151634
rect 471286 151398 501770 151634
rect 502006 151398 532490 151634
rect 532726 151398 563210 151634
rect 563446 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 69808 147454
rect 70044 147218 163512 147454
rect 163748 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 222952 147454
rect 223188 147218 232882 147454
rect 233118 147218 242813 147454
rect 243049 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 312618 147454
rect 312854 147218 315882 147454
rect 316118 147218 319146 147454
rect 319382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 394250 147454
rect 394486 147218 424970 147454
rect 425206 147218 455690 147454
rect 455926 147218 486410 147454
rect 486646 147218 517130 147454
rect 517366 147218 547850 147454
rect 548086 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 69808 147134
rect 70044 146898 163512 147134
rect 163748 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 222952 147134
rect 223188 146898 232882 147134
rect 233118 146898 242813 147134
rect 243049 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 312618 147134
rect 312854 146898 315882 147134
rect 316118 146898 319146 147134
rect 319382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 394250 147134
rect 394486 146898 424970 147134
rect 425206 146898 455690 147134
rect 455926 146898 486410 147134
rect 486646 146898 517130 147134
rect 517366 146898 547850 147134
rect 548086 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 69128 115954
rect 69364 115718 164192 115954
rect 164428 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 227916 115954
rect 228152 115718 237847 115954
rect 238083 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 314250 115954
rect 314486 115718 317514 115954
rect 317750 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 409610 115954
rect 409846 115718 440330 115954
rect 440566 115718 471050 115954
rect 471286 115718 501770 115954
rect 502006 115718 532490 115954
rect 532726 115718 563210 115954
rect 563446 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 69128 115634
rect 69364 115398 164192 115634
rect 164428 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 227916 115634
rect 228152 115398 237847 115634
rect 238083 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 314250 115634
rect 314486 115398 317514 115634
rect 317750 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 409610 115634
rect 409846 115398 440330 115634
rect 440566 115398 471050 115634
rect 471286 115398 501770 115634
rect 502006 115398 532490 115634
rect 532726 115398 563210 115634
rect 563446 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 69808 111454
rect 70044 111218 163512 111454
rect 163748 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 222952 111454
rect 223188 111218 232882 111454
rect 233118 111218 242813 111454
rect 243049 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 312618 111454
rect 312854 111218 315882 111454
rect 316118 111218 319146 111454
rect 319382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 394250 111454
rect 394486 111218 424970 111454
rect 425206 111218 455690 111454
rect 455926 111218 486410 111454
rect 486646 111218 517130 111454
rect 517366 111218 547850 111454
rect 548086 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 69808 111134
rect 70044 110898 163512 111134
rect 163748 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 222952 111134
rect 223188 110898 232882 111134
rect 233118 110898 242813 111134
rect 243049 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 312618 111134
rect 312854 110898 315882 111134
rect 316118 110898 319146 111134
rect 319382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 394250 111134
rect 394486 110898 424970 111134
rect 425206 110898 455690 111134
rect 455926 110898 486410 111134
rect 486646 110898 517130 111134
rect 517366 110898 547850 111134
rect 548086 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use sky130_sram_1kbyte_1rw1r_32x256_8  openram_1kB
timestamp 0
transform 1 0 68800 0 1 95100
box 0 0 95956 79500
use wb_bridge_2way  wb_bridge_2way
timestamp 0
transform 1 0 310000 0 1 96000
box 0 144 12000 80000
use wb_openram_wrapper  wb_openram_wrapper
timestamp 0
transform 1 0 217000 0 1 96000
box 0 144 32000 79688
use wrapped_etpu  wrapped_etpu_3
timestamp 0
transform 1 0 390000 0 1 96000
box -10 0 180000 180000
use wrapped_function_generator  wrapped_function_generator_0
timestamp 0
transform 1 0 70000 0 1 240000
box 0 0 50000 52000
use wrapped_ibnalhaytham  wrapped_ibnalhaytham_1
timestamp 0
transform 1 0 180000 0 1 240000
box 0 0 113010 115154
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 93100 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 176600 74414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 294000 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 93100 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 176600 110414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 294000 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 93100 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 176600 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 357154 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 94000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 178000 218414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 357154 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 357154 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 357154 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 94000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 278000 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 94000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 278000 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 94000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 278000 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 94000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 278000 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 94000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 278000 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 93100 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 176600 83414 238000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 294000 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 93100 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 176600 119414 238000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 294000 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 93100 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 176600 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 238000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 357154 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 94000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 178000 227414 238000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 357154 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 238000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 357154 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 94000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 278000 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 94000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 278000 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 94000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 278000 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 94000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 278000 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 94000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 278000 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 93100 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 176600 92414 238000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 294000 92414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 93100 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 176600 128414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 93100 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 176600 164414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 238000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 357154 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 94000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 178000 236414 238000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 357154 236414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 238000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 357154 272414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 94000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 178000 308414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 94000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 278000 416414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 94000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 278000 452414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 94000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 278000 488414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 94000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 278000 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 94000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 278000 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 -7654 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 -7654 101414 93100 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 294000 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 93100 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 176600 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 -7654 209414 238000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 357154 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 -7654 245414 94000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 357154 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 -7654 281414 238000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 357154 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 -7654 317414 94000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 178000 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 -7654 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 -7654 389414 94000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 278000 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 94000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 278000 425414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 94000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 278000 461414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 94000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 278000 497414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 94000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 278000 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 94000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 278000 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 93100 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 294000 96914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 93100 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 176600 132914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 238000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 357154 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 94000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 357154 240914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 238000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 357154 276914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 94000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 178000 312914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 94000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 278000 420914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 94000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 278000 456914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 94000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 278000 492914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 94000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 278000 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 94000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 278000 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 93100 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 176600 69914 238000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 294000 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 93100 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 176600 105914 238000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 294000 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 93100 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 176600 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 238000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 357154 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 94000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 178000 249914 238000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 357154 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 238000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 357154 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 94000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 178000 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 94000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 278000 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 94000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 278000 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 94000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 278000 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 94000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 278000 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 94000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 278000 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 93100 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 176600 78914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 294000 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 93100 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 176600 114914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 294000 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 93100 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 176600 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 357154 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 94000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 178000 222914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 357154 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 357154 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 357154 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 94000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 278000 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 94000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 278000 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 94000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 278000 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 94000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 278000 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 94000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 278000 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 93100 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 176600 87914 238000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 294000 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 93100 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 176600 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 93100 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 176600 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 238000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 357154 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 94000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 178000 231914 238000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 357154 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 238000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 357154 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 94000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 278000 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 94000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 278000 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 94000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 278000 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 94000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 278000 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 94000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 278000 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
