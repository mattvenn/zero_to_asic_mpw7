magic
tech sky130B
magscale 1 2
timestamp 1661625863
<< obsli1 >>
rect 0 0 584000 704000
<< metal1 >>
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 301498 702652 301504 702704
rect 301556 702692 301562 702704
rect 494790 702692 494796 702704
rect 301556 702664 494796 702692
rect 301556 702652 301562 702664
rect 494790 702652 494796 702664
rect 494848 702652 494854 702704
rect 209774 702584 209780 702636
rect 209832 702624 209838 702636
rect 462314 702624 462320 702636
rect 209832 702596 462320 702624
rect 209832 702584 209838 702596
rect 462314 702584 462320 702596
rect 462372 702584 462378 702636
rect 177942 702516 177948 702568
rect 178000 702556 178006 702568
rect 478506 702556 478512 702568
rect 178000 702528 478512 702556
rect 178000 702516 178006 702528
rect 478506 702516 478512 702528
rect 478564 702516 478570 702568
rect 206278 702448 206284 702500
rect 206336 702488 206342 702500
rect 559650 702488 559656 702500
rect 206336 702460 559656 702488
rect 206336 702448 206342 702460
rect 559650 702448 559656 702460
rect 559708 702448 559714 702500
rect 72970 700340 72976 700392
rect 73028 700380 73034 700392
rect 82078 700380 82084 700392
rect 73028 700352 82084 700380
rect 73028 700340 73034 700352
rect 82078 700340 82084 700352
rect 82136 700340 82142 700392
rect 105446 700340 105452 700392
rect 105504 700380 105510 700392
rect 193214 700380 193220 700392
rect 105504 700352 193220 700380
rect 105504 700340 105510 700352
rect 193214 700340 193220 700352
rect 193272 700340 193278 700392
rect 235166 700340 235172 700392
rect 235224 700380 235230 700392
rect 304994 700380 305000 700392
rect 235224 700352 305000 700380
rect 235224 700340 235230 700352
rect 304994 700340 305000 700352
rect 305052 700340 305058 700392
rect 24302 700272 24308 700324
rect 24360 700312 24366 700324
rect 43438 700312 43444 700324
rect 24360 700284 43444 700312
rect 24360 700272 24366 700284
rect 43438 700272 43444 700284
rect 43496 700272 43502 700324
rect 62758 700272 62764 700324
rect 62816 700312 62822 700324
rect 170306 700312 170312 700324
rect 62816 700284 170312 700312
rect 62816 700272 62822 700284
rect 170306 700272 170312 700284
rect 170364 700272 170370 700324
rect 218974 700272 218980 700324
rect 219032 700312 219038 700324
rect 310514 700312 310520 700324
rect 219032 700284 310520 700312
rect 219032 700272 219038 700284
rect 310514 700272 310520 700284
rect 310572 700272 310578 700324
rect 319438 700272 319444 700324
rect 319496 700312 319502 700324
rect 429838 700312 429844 700324
rect 319496 700284 429844 700312
rect 319496 700272 319502 700284
rect 429838 700272 429844 700284
rect 429896 700272 429902 700324
rect 300118 699660 300124 699712
rect 300176 699700 300182 699712
rect 306466 699700 306472 699712
rect 300176 699672 306472 699700
rect 300176 699660 300182 699672
rect 306466 699660 306472 699672
rect 306524 699660 306530 699712
rect 525058 699660 525064 699712
rect 525116 699700 525122 699712
rect 527174 699700 527180 699712
rect 525116 699672 527180 699700
rect 525116 699660 525122 699672
rect 527174 699660 527180 699672
rect 527232 699660 527238 699712
rect 324958 698912 324964 698964
rect 325016 698952 325022 698964
rect 397454 698952 397460 698964
rect 325016 698924 397460 698952
rect 325016 698912 325022 698924
rect 397454 698912 397460 698924
rect 397512 698912 397518 698964
rect 266354 697620 266360 697672
rect 266412 697660 266418 697672
rect 267642 697660 267648 697672
rect 266412 697632 267648 697660
rect 266412 697620 266418 697632
rect 267642 697620 267648 697632
rect 267700 697620 267706 697672
rect 211798 697552 211804 697604
rect 211856 697592 211862 697604
rect 348786 697592 348792 697604
rect 211856 697564 348792 697592
rect 211856 697552 211862 697564
rect 348786 697552 348792 697564
rect 348844 697552 348850 697604
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 189718 683176 189724 683188
rect 3476 683148 189724 683176
rect 3476 683136 3482 683148
rect 189718 683136 189724 683148
rect 189776 683136 189782 683188
rect 297358 683136 297364 683188
rect 297416 683176 297422 683188
rect 580166 683176 580172 683188
rect 297416 683148 580172 683176
rect 297416 683136 297422 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 22738 670732 22744 670744
rect 3568 670704 22744 670732
rect 3568 670692 3574 670704
rect 22738 670692 22744 670704
rect 22796 670692 22802 670744
rect 2774 656956 2780 657008
rect 2832 656996 2838 657008
rect 4798 656996 4804 657008
rect 2832 656968 4804 656996
rect 2832 656956 2838 656968
rect 4798 656956 4804 656968
rect 4856 656956 4862 657008
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 44818 632108 44824 632120
rect 3476 632080 44824 632108
rect 3476 632068 3482 632080
rect 44818 632068 44824 632080
rect 44876 632068 44882 632120
rect 179322 630640 179328 630692
rect 179380 630680 179386 630692
rect 579982 630680 579988 630692
rect 179380 630652 579988 630680
rect 179380 630640 179386 630652
rect 579982 630640 579988 630652
rect 580040 630640 580046 630692
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 18598 618304 18604 618316
rect 3200 618276 18604 618304
rect 3200 618264 3206 618276
rect 18598 618264 18604 618276
rect 18656 618264 18662 618316
rect 337378 616836 337384 616888
rect 337436 616876 337442 616888
rect 580166 616876 580172 616888
rect 337436 616848 580172 616876
rect 337436 616836 337442 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3418 606024 3424 606076
rect 3476 606064 3482 606076
rect 8938 606064 8944 606076
rect 3476 606036 8944 606064
rect 3476 606024 3482 606036
rect 8938 606024 8944 606036
rect 8996 606024 9002 606076
rect 309778 590656 309784 590708
rect 309836 590696 309842 590708
rect 580166 590696 580172 590708
rect 309836 590668 580172 590696
rect 309836 590656 309842 590668
rect 580166 590656 580172 590668
rect 580224 590656 580230 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 116578 579680 116584 579692
rect 3384 579652 116584 579680
rect 3384 579640 3390 579652
rect 116578 579640 116584 579652
rect 116636 579640 116642 579692
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 21358 565876 21364 565888
rect 3476 565848 21364 565876
rect 3476 565836 3482 565848
rect 21358 565836 21364 565848
rect 21416 565836 21422 565888
rect 158622 563048 158628 563100
rect 158680 563088 158686 563100
rect 579890 563088 579896 563100
rect 158680 563060 579896 563088
rect 158680 563048 158686 563060
rect 579890 563048 579896 563060
rect 579948 563048 579954 563100
rect 3418 553392 3424 553444
rect 3476 553432 3482 553444
rect 17218 553432 17224 553444
rect 3476 553404 17224 553432
rect 3476 553392 3482 553404
rect 17218 553392 17224 553404
rect 17276 553392 17282 553444
rect 3418 527144 3424 527196
rect 3476 527184 3482 527196
rect 13078 527184 13084 527196
rect 3476 527156 13084 527184
rect 3476 527144 3482 527156
rect 13078 527144 13084 527156
rect 13136 527144 13142 527196
rect 347038 524424 347044 524476
rect 347096 524464 347102 524476
rect 580166 524464 580172 524476
rect 347096 524436 580172 524464
rect 347096 524424 347102 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 400858 510620 400864 510672
rect 400916 510660 400922 510672
rect 580166 510660 580172 510672
rect 400916 510632 580172 510660
rect 400916 510620 400922 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3050 474716 3056 474768
rect 3108 474756 3114 474768
rect 202874 474756 202880 474768
rect 3108 474728 202880 474756
rect 3108 474716 3114 474728
rect 202874 474716 202880 474728
rect 202932 474716 202938 474768
rect 278038 470568 278044 470620
rect 278096 470608 278102 470620
rect 580166 470608 580172 470620
rect 278096 470580 580172 470608
rect 278096 470568 278102 470580
rect 580166 470568 580172 470580
rect 580224 470568 580230 470620
rect 3510 462340 3516 462392
rect 3568 462380 3574 462392
rect 111058 462380 111064 462392
rect 3568 462352 111064 462380
rect 3568 462340 3574 462352
rect 111058 462340 111064 462352
rect 111116 462340 111122 462392
rect 166902 456764 166908 456816
rect 166960 456804 166966 456816
rect 580166 456804 580172 456816
rect 166960 456776 580172 456804
rect 166960 456764 166966 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 39298 448576 39304 448588
rect 3200 448548 39304 448576
rect 3200 448536 3206 448548
rect 39298 448536 39304 448548
rect 39356 448536 39362 448588
rect 3510 422288 3516 422340
rect 3568 422328 3574 422340
rect 32398 422328 32404 422340
rect 3568 422300 32404 422328
rect 3568 422288 3574 422300
rect 32398 422288 32404 422300
rect 32456 422288 32462 422340
rect 2866 409844 2872 409896
rect 2924 409884 2930 409896
rect 53098 409884 53104 409896
rect 2924 409856 53104 409884
rect 2924 409844 2930 409856
rect 53098 409844 53104 409856
rect 53156 409844 53162 409896
rect 160830 404336 160836 404388
rect 160888 404376 160894 404388
rect 579982 404376 579988 404388
rect 160888 404348 579988 404376
rect 160888 404336 160894 404348
rect 579982 404336 579988 404348
rect 580040 404336 580046 404388
rect 3510 397468 3516 397520
rect 3568 397508 3574 397520
rect 58618 397508 58624 397520
rect 3568 397480 58624 397508
rect 3568 397468 3574 397480
rect 58618 397468 58624 397480
rect 58676 397468 58682 397520
rect 220078 378156 220084 378208
rect 220136 378196 220142 378208
rect 580166 378196 580172 378208
rect 220136 378168 580172 378196
rect 220136 378156 220142 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 179414 377408 179420 377460
rect 179472 377448 179478 377460
rect 266354 377448 266360 377460
rect 179472 377420 266360 377448
rect 179472 377408 179478 377420
rect 266354 377408 266360 377420
rect 266412 377408 266418 377460
rect 195882 375980 195888 376032
rect 195940 376020 195946 376032
rect 331214 376020 331220 376032
rect 195940 375992 331220 376020
rect 195940 375980 195946 375992
rect 331214 375980 331220 375992
rect 331272 375980 331278 376032
rect 179046 374620 179052 374672
rect 179104 374660 179110 374672
rect 580258 374660 580264 374672
rect 179104 374632 580264 374660
rect 179104 374620 179110 374632
rect 580258 374620 580264 374632
rect 580316 374620 580322 374672
rect 122742 373260 122748 373312
rect 122800 373300 122806 373312
rect 201494 373300 201500 373312
rect 122800 373272 201500 373300
rect 122800 373260 122806 373272
rect 201494 373260 201500 373272
rect 201552 373260 201558 373312
rect 189718 371832 189724 371884
rect 189776 371872 189782 371884
rect 198734 371872 198740 371884
rect 189776 371844 198740 371872
rect 189776 371832 189782 371844
rect 198734 371832 198740 371844
rect 198792 371832 198798 371884
rect 3510 371220 3516 371272
rect 3568 371260 3574 371272
rect 128354 371260 128360 371272
rect 3568 371232 128360 371260
rect 3568 371220 3574 371232
rect 128354 371220 128360 371232
rect 128412 371220 128418 371272
rect 206370 371220 206376 371272
rect 206428 371260 206434 371272
rect 327718 371260 327724 371272
rect 206428 371232 327724 371260
rect 206428 371220 206434 371232
rect 327718 371220 327724 371232
rect 327776 371220 327782 371272
rect 179138 370472 179144 370524
rect 179196 370512 179202 370524
rect 580350 370512 580356 370524
rect 179196 370484 580356 370512
rect 179196 370472 179202 370484
rect 580350 370472 580356 370484
rect 580408 370472 580414 370524
rect 209038 369112 209044 369164
rect 209096 369152 209102 369164
rect 220078 369152 220084 369164
rect 209096 369124 220084 369152
rect 209096 369112 209102 369124
rect 220078 369112 220084 369124
rect 220136 369112 220142 369164
rect 39298 368908 39304 368960
rect 39356 368948 39362 368960
rect 39942 368948 39948 368960
rect 39356 368920 39948 368948
rect 39356 368908 39362 368920
rect 39942 368908 39948 368920
rect 40000 368908 40006 368960
rect 194594 368908 194600 368960
rect 194652 368948 194658 368960
rect 195882 368948 195888 368960
rect 194652 368920 195888 368948
rect 194652 368908 194658 368920
rect 195882 368908 195888 368920
rect 195940 368908 195946 368960
rect 64690 368568 64696 368620
rect 64748 368608 64754 368620
rect 194594 368608 194600 368620
rect 64748 368580 194600 368608
rect 64748 368568 64754 368580
rect 194594 368568 194600 368580
rect 194652 368568 194658 368620
rect 39942 368500 39948 368552
rect 40000 368540 40006 368552
rect 295610 368540 295616 368552
rect 40000 368512 295616 368540
rect 40000 368500 40006 368512
rect 295610 368500 295616 368512
rect 295668 368500 295674 368552
rect 109034 367072 109040 367124
rect 109092 367112 109098 367124
rect 254578 367112 254584 367124
rect 109092 367084 254584 367112
rect 109092 367072 109098 367084
rect 254578 367072 254584 367084
rect 254636 367072 254642 367124
rect 142798 365780 142804 365832
rect 142856 365820 142862 365832
rect 276014 365820 276020 365832
rect 142856 365792 276020 365820
rect 142856 365780 142862 365792
rect 276014 365780 276020 365792
rect 276072 365780 276078 365832
rect 124858 365712 124864 365764
rect 124916 365752 124922 365764
rect 287054 365752 287060 365764
rect 124916 365724 287060 365752
rect 124916 365712 124922 365724
rect 287054 365712 287060 365724
rect 287112 365712 287118 365764
rect 190454 364488 190460 364540
rect 190512 364528 190518 364540
rect 315298 364528 315304 364540
rect 190512 364500 315304 364528
rect 190512 364488 190518 364500
rect 315298 364488 315304 364500
rect 315356 364488 315362 364540
rect 69198 364420 69204 364472
rect 69256 364460 69262 364472
rect 242894 364460 242900 364472
rect 69256 364432 242900 364460
rect 69256 364420 69262 364432
rect 242894 364420 242900 364432
rect 242952 364420 242958 364472
rect 179874 364352 179880 364404
rect 179932 364392 179938 364404
rect 580166 364392 580172 364404
rect 179932 364364 580172 364392
rect 179932 364352 179938 364364
rect 580166 364352 580172 364364
rect 580224 364352 580230 364404
rect 117958 363060 117964 363112
rect 118016 363100 118022 363112
rect 214466 363100 214472 363112
rect 118016 363072 214472 363100
rect 118016 363060 118022 363072
rect 214466 363060 214472 363072
rect 214524 363060 214530 363112
rect 130378 362992 130384 363044
rect 130436 363032 130442 363044
rect 295334 363032 295340 363044
rect 130436 363004 295340 363032
rect 130436 362992 130442 363004
rect 295334 362992 295340 363004
rect 295392 362992 295398 363044
rect 179230 362924 179236 362976
rect 179288 362964 179294 362976
rect 580258 362964 580264 362976
rect 179288 362936 580264 362964
rect 179288 362924 179294 362936
rect 580258 362924 580264 362936
rect 580316 362924 580322 362976
rect 282914 362176 282920 362228
rect 282972 362216 282978 362228
rect 295426 362216 295432 362228
rect 282972 362188 295432 362216
rect 282972 362176 282978 362188
rect 295426 362176 295432 362188
rect 295484 362176 295490 362228
rect 174722 361700 174728 361752
rect 174780 361740 174786 361752
rect 237466 361740 237472 361752
rect 174780 361712 237472 361740
rect 174780 361700 174786 361712
rect 237466 361700 237472 361712
rect 237524 361700 237530 361752
rect 273530 361700 273536 361752
rect 273588 361740 273594 361752
rect 278038 361740 278044 361752
rect 273588 361712 278044 361740
rect 273588 361700 273594 361712
rect 278038 361700 278044 361712
rect 278096 361700 278102 361752
rect 134518 361632 134524 361684
rect 134576 361672 134582 361684
rect 256786 361672 256792 361684
rect 134576 361644 256792 361672
rect 134576 361632 134582 361644
rect 256786 361632 256792 361644
rect 256844 361632 256850 361684
rect 79318 361564 79324 361616
rect 79376 361604 79382 361616
rect 245838 361604 245844 361616
rect 79376 361576 245844 361604
rect 79376 361564 79382 361576
rect 245838 361564 245844 361576
rect 245896 361564 245902 361616
rect 162762 360476 162768 360528
rect 162820 360516 162826 360528
rect 197722 360516 197728 360528
rect 162820 360488 197728 360516
rect 162820 360476 162826 360488
rect 197722 360476 197728 360488
rect 197780 360476 197786 360528
rect 126238 360408 126244 360460
rect 126296 360448 126302 360460
rect 201586 360448 201592 360460
rect 126296 360420 201592 360448
rect 126296 360408 126302 360420
rect 201586 360408 201592 360420
rect 201644 360408 201650 360460
rect 225414 360408 225420 360460
rect 225472 360448 225478 360460
rect 303614 360448 303620 360460
rect 225472 360420 303620 360448
rect 225472 360408 225478 360420
rect 303614 360408 303620 360420
rect 303672 360408 303678 360460
rect 167638 360340 167644 360392
rect 167696 360380 167702 360392
rect 279326 360380 279332 360392
rect 167696 360352 279332 360380
rect 167696 360340 167702 360352
rect 279326 360340 279332 360352
rect 279384 360340 279390 360392
rect 170398 360272 170404 360324
rect 170456 360312 170462 360324
rect 291838 360312 291844 360324
rect 170456 360284 291844 360312
rect 170456 360272 170462 360284
rect 291838 360272 291844 360284
rect 291896 360272 291902 360324
rect 69106 360204 69112 360256
rect 69164 360244 69170 360256
rect 220262 360244 220268 360256
rect 69164 360216 220268 360244
rect 69164 360204 69170 360216
rect 220262 360204 220268 360216
rect 220320 360204 220326 360256
rect 254394 360204 254400 360256
rect 254452 360244 254458 360256
rect 254578 360244 254584 360256
rect 254452 360216 254584 360244
rect 254452 360204 254458 360216
rect 254578 360204 254584 360216
rect 254636 360244 254642 360256
rect 373258 360244 373264 360256
rect 254636 360216 373264 360244
rect 254636 360204 254642 360216
rect 373258 360204 373264 360216
rect 373316 360204 373322 360256
rect 144178 359048 144184 359100
rect 144236 359088 144242 359100
rect 283374 359088 283380 359100
rect 144236 359060 283380 359088
rect 144236 359048 144242 359060
rect 283374 359048 283380 359060
rect 283432 359048 283438 359100
rect 157242 358980 157248 359032
rect 157300 359020 157306 359032
rect 184934 359020 184940 359032
rect 157300 358992 184940 359020
rect 157300 358980 157306 358992
rect 184934 358980 184940 358992
rect 184992 358980 184998 359032
rect 282086 358912 282092 358964
rect 282144 358952 282150 358964
rect 311894 358952 311900 358964
rect 282144 358924 311900 358952
rect 282144 358912 282150 358924
rect 311894 358912 311900 358924
rect 311952 358912 311958 358964
rect 181622 358844 181628 358896
rect 181680 358884 181686 358896
rect 349154 358884 349160 358896
rect 181680 358856 349160 358884
rect 181680 358844 181686 358856
rect 349154 358844 349160 358856
rect 349212 358844 349218 358896
rect 101398 358776 101404 358828
rect 101456 358816 101462 358828
rect 294138 358816 294144 358828
rect 101456 358788 294144 358816
rect 101456 358776 101462 358788
rect 294138 358776 294144 358788
rect 294196 358776 294202 358828
rect 187418 358028 187424 358080
rect 187476 358068 187482 358080
rect 206370 358068 206376 358080
rect 187476 358040 206376 358068
rect 187476 358028 187482 358040
rect 206370 358028 206376 358040
rect 206428 358028 206434 358080
rect 269022 357824 269028 357876
rect 269080 357864 269086 357876
rect 349246 357864 349252 357876
rect 269080 357836 349252 357864
rect 269080 357824 269086 357836
rect 349246 357824 349252 357836
rect 349304 357824 349310 357876
rect 242802 357756 242808 357808
rect 242860 357796 242866 357808
rect 270494 357796 270500 357808
rect 242860 357768 270500 357796
rect 242860 357756 242866 357768
rect 270494 357756 270500 357768
rect 270552 357756 270558 357808
rect 174630 357688 174636 357740
rect 174688 357728 174694 357740
rect 241514 357728 241520 357740
rect 174688 357700 241520 357728
rect 174688 357688 174694 357700
rect 241514 357688 241520 357700
rect 241572 357688 241578 357740
rect 260742 357688 260748 357740
rect 260800 357728 260806 357740
rect 296806 357728 296812 357740
rect 260800 357700 296812 357728
rect 260800 357688 260806 357700
rect 296806 357688 296812 357700
rect 296864 357688 296870 357740
rect 179782 357620 179788 357672
rect 179840 357660 179846 357672
rect 211798 357660 211804 357672
rect 179840 357632 211804 357660
rect 179840 357620 179846 357632
rect 211798 357620 211804 357632
rect 211856 357620 211862 357672
rect 223482 357620 223488 357672
rect 223540 357660 223546 357672
rect 291746 357660 291752 357672
rect 223540 357632 291752 357660
rect 223540 357620 223546 357632
rect 291746 357620 291752 357632
rect 291804 357620 291810 357672
rect 148318 357552 148324 357604
rect 148376 357592 148382 357604
rect 193214 357592 193220 357604
rect 148376 357564 193220 357592
rect 148376 357552 148382 357564
rect 193214 357552 193220 357564
rect 193272 357552 193278 357604
rect 217042 357552 217048 357604
rect 217100 357592 217106 357604
rect 317414 357592 317420 357604
rect 217100 357564 317420 357592
rect 217100 357552 217106 357564
rect 317414 357552 317420 357564
rect 317472 357552 317478 357604
rect 3050 357484 3056 357536
rect 3108 357524 3114 357536
rect 90358 357524 90364 357536
rect 3108 357496 90364 357524
rect 3108 357484 3114 357496
rect 90358 357484 90364 357496
rect 90416 357484 90422 357536
rect 107654 357484 107660 357536
rect 107712 357524 107718 357536
rect 289446 357524 289452 357536
rect 107712 357496 289452 357524
rect 107712 357484 107718 357496
rect 289446 357484 289452 357496
rect 289504 357484 289510 357536
rect 290458 357484 290464 357536
rect 290516 357524 290522 357536
rect 308398 357524 308404 357536
rect 290516 357496 308404 357524
rect 290516 357484 290522 357496
rect 308398 357484 308404 357496
rect 308456 357484 308462 357536
rect 55030 357416 55036 357468
rect 55088 357456 55094 357468
rect 265158 357456 265164 357468
rect 55088 357428 265164 357456
rect 55088 357416 55094 357428
rect 265158 357416 265164 357428
rect 265216 357416 265222 357468
rect 287146 357416 287152 357468
rect 287204 357456 287210 357468
rect 293310 357456 293316 357468
rect 287204 357428 293316 357456
rect 287204 357416 287210 357428
rect 293310 357416 293316 357428
rect 293368 357416 293374 357468
rect 154022 357348 154028 357400
rect 154080 357388 154086 357400
rect 242802 357388 242808 357400
rect 154080 357360 242808 357388
rect 154080 357348 154086 357360
rect 242802 357348 242808 357360
rect 242860 357348 242866 357400
rect 68646 356668 68652 356720
rect 68704 356708 68710 356720
rect 153194 356708 153200 356720
rect 68704 356680 153200 356708
rect 68704 356668 68710 356680
rect 153194 356668 153200 356680
rect 153252 356708 153258 356720
rect 154022 356708 154028 356720
rect 153252 356680 154028 356708
rect 153252 356668 153258 356680
rect 154022 356668 154028 356680
rect 154080 356668 154086 356720
rect 174538 356328 174544 356380
rect 174596 356368 174602 356380
rect 208762 356368 208768 356380
rect 174596 356340 208768 356368
rect 174596 356328 174602 356340
rect 208762 356328 208768 356340
rect 208820 356328 208826 356380
rect 258902 356328 258908 356380
rect 258960 356368 258966 356380
rect 299566 356368 299572 356380
rect 258960 356340 299572 356368
rect 258960 356328 258966 356340
rect 299566 356328 299572 356340
rect 299624 356328 299630 356380
rect 171870 356260 171876 356312
rect 171928 356300 171934 356312
rect 273530 356300 273536 356312
rect 171928 356272 273536 356300
rect 171928 356260 171934 356272
rect 273530 356260 273536 356272
rect 273588 356260 273594 356312
rect 285950 356260 285956 356312
rect 286008 356300 286014 356312
rect 313274 356300 313280 356312
rect 286008 356272 313280 356300
rect 286008 356260 286014 356272
rect 313274 356260 313280 356272
rect 313332 356260 313338 356312
rect 140130 356192 140136 356244
rect 140188 356232 140194 356244
rect 247954 356232 247960 356244
rect 140188 356204 247960 356232
rect 140188 356192 140194 356204
rect 247954 356192 247960 356204
rect 248012 356192 248018 356244
rect 252462 356192 252468 356244
rect 252520 356232 252526 356244
rect 301590 356232 301596 356244
rect 252520 356204 301596 356232
rect 252520 356192 252526 356204
rect 301590 356192 301596 356204
rect 301648 356192 301654 356244
rect 111150 356124 111156 356176
rect 111208 356164 111214 356176
rect 295518 356164 295524 356176
rect 111208 356136 295524 356164
rect 111208 356124 111214 356136
rect 295518 356124 295524 356136
rect 295576 356124 295582 356176
rect 80054 356056 80060 356108
rect 80112 356096 80118 356108
rect 298186 356096 298192 356108
rect 80112 356068 298192 356096
rect 80112 356056 80118 356068
rect 298186 356056 298192 356068
rect 298244 356056 298250 356108
rect 289446 355988 289452 356040
rect 289504 356028 289510 356040
rect 294230 356028 294236 356040
rect 289504 356000 294236 356028
rect 289504 355988 289510 356000
rect 294230 355988 294236 356000
rect 294288 355988 294294 356040
rect 111058 355308 111064 355360
rect 111116 355348 111122 355360
rect 135254 355348 135260 355360
rect 111116 355320 135260 355348
rect 111116 355308 111122 355320
rect 135254 355308 135260 355320
rect 135312 355308 135318 355360
rect 202874 355240 202880 355292
rect 202932 355280 202938 355292
rect 203840 355280 203846 355292
rect 202932 355252 203846 355280
rect 202932 355240 202938 355252
rect 203840 355240 203846 355252
rect 203898 355240 203904 355292
rect 171778 355036 171784 355088
rect 171836 355076 171842 355088
rect 198734 355076 198740 355088
rect 171836 355048 198740 355076
rect 171836 355036 171842 355048
rect 198734 355036 198740 355048
rect 198792 355076 198798 355088
rect 199654 355076 199660 355088
rect 198792 355048 199660 355076
rect 198792 355036 198798 355048
rect 199654 355036 199660 355048
rect 199712 355036 199718 355088
rect 169018 354968 169024 355020
rect 169076 355008 169082 355020
rect 202874 355008 202880 355020
rect 169076 354980 202880 355008
rect 169076 354968 169082 354980
rect 202874 354968 202880 354980
rect 202932 354968 202938 355020
rect 275646 354968 275652 355020
rect 275704 355008 275710 355020
rect 299750 355008 299756 355020
rect 275704 354980 299756 355008
rect 275704 354968 275710 354980
rect 299750 354968 299756 354980
rect 299808 354968 299814 355020
rect 175918 354900 175924 354952
rect 175976 354940 175982 354952
rect 235074 354940 235080 354952
rect 175976 354912 235080 354940
rect 175976 354900 175982 354912
rect 235074 354900 235080 354912
rect 235132 354900 235138 354952
rect 256786 354900 256792 354952
rect 256844 354940 256850 354952
rect 297450 354940 297456 354952
rect 256844 354912 297456 354940
rect 256844 354900 256850 354912
rect 297450 354900 297456 354912
rect 297508 354900 297514 354952
rect 97258 354832 97264 354884
rect 97316 354872 97322 354884
rect 293034 354872 293040 354884
rect 97316 354844 293040 354872
rect 97316 354832 97322 354844
rect 293034 354832 293040 354844
rect 293092 354832 293098 354884
rect 75914 354764 75920 354816
rect 75972 354804 75978 354816
rect 294046 354804 294052 354816
rect 75972 354776 294052 354804
rect 75972 354764 75978 354776
rect 294046 354764 294052 354776
rect 294104 354764 294110 354816
rect 135254 354696 135260 354748
rect 135312 354736 135318 354748
rect 266630 354736 266636 354748
rect 135312 354708 266636 354736
rect 135312 354696 135318 354708
rect 266630 354696 266636 354708
rect 266688 354696 266694 354748
rect 279510 354696 279516 354748
rect 279568 354736 279574 354748
rect 449158 354736 449164 354748
rect 279568 354708 449164 354736
rect 279568 354696 279574 354708
rect 449158 354696 449164 354708
rect 449216 354696 449222 354748
rect 84286 354016 84292 354068
rect 84344 354056 84350 354068
rect 179782 354056 179788 354068
rect 84344 354028 179788 354056
rect 84344 354016 84350 354028
rect 179782 354016 179788 354028
rect 179840 354016 179846 354068
rect 44818 353948 44824 354000
rect 44876 353988 44882 354000
rect 45462 353988 45468 354000
rect 44876 353960 45468 353988
rect 44876 353948 44882 353960
rect 45462 353948 45468 353960
rect 45520 353988 45526 354000
rect 176654 353988 176660 354000
rect 45520 353960 176660 353988
rect 45520 353948 45526 353960
rect 176654 353948 176660 353960
rect 176712 353948 176718 354000
rect 293310 353948 293316 354000
rect 293368 353988 293374 354000
rect 580350 353988 580356 354000
rect 293368 353960 580356 353988
rect 293368 353948 293374 353960
rect 580350 353948 580356 353960
rect 580408 353948 580414 354000
rect 177850 353268 177856 353320
rect 177908 353308 177914 353320
rect 179874 353308 179880 353320
rect 177908 353280 179880 353308
rect 177908 353268 177914 353280
rect 179874 353268 179880 353280
rect 179932 353268 179938 353320
rect 113174 352520 113180 352572
rect 113232 352560 113238 352572
rect 179598 352560 179604 352572
rect 113232 352532 179604 352560
rect 113232 352520 113238 352532
rect 179598 352520 179604 352532
rect 179656 352520 179662 352572
rect 50890 351160 50896 351212
rect 50948 351200 50954 351212
rect 174722 351200 174728 351212
rect 50948 351172 174728 351200
rect 50948 351160 50954 351172
rect 174722 351160 174728 351172
rect 174780 351160 174786 351212
rect 293126 351160 293132 351212
rect 293184 351200 293190 351212
rect 580258 351200 580264 351212
rect 293184 351172 580264 351200
rect 293184 351160 293190 351172
rect 580258 351160 580264 351172
rect 580316 351160 580322 351212
rect 127710 347760 127716 347812
rect 127768 347800 127774 347812
rect 176654 347800 176660 347812
rect 127768 347772 176660 347800
rect 127768 347760 127774 347772
rect 176654 347760 176660 347772
rect 176712 347760 176718 347812
rect 6914 347012 6920 347064
rect 6972 347052 6978 347064
rect 62850 347052 62856 347064
rect 6972 347024 62856 347052
rect 6972 347012 6978 347024
rect 62850 347012 62856 347024
rect 62908 347012 62914 347064
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 25498 345080 25504 345092
rect 3384 345052 25504 345080
rect 3384 345040 3390 345052
rect 25498 345040 25504 345052
rect 25556 345040 25562 345092
rect 296162 345040 296168 345092
rect 296220 345080 296226 345092
rect 472618 345080 472624 345092
rect 296220 345052 472624 345080
rect 296220 345040 296226 345052
rect 472618 345040 472624 345052
rect 472676 345040 472682 345092
rect 72418 344292 72424 344344
rect 72476 344332 72482 344344
rect 174630 344332 174636 344344
rect 72476 344304 174636 344332
rect 72476 344292 72482 344304
rect 174630 344292 174636 344304
rect 174688 344292 174694 344344
rect 295334 343544 295340 343596
rect 295392 343584 295398 343596
rect 295610 343584 295616 343596
rect 295392 343556 295616 343584
rect 295392 343544 295398 343556
rect 295610 343544 295616 343556
rect 295668 343544 295674 343596
rect 295334 342864 295340 342916
rect 295392 342904 295398 342916
rect 295392 342876 296714 342904
rect 295392 342864 295398 342876
rect 296686 342768 296714 342876
rect 300854 342768 300860 342780
rect 296686 342740 300860 342768
rect 300854 342728 300860 342740
rect 300912 342768 300918 342780
rect 301498 342768 301504 342780
rect 300912 342740 301504 342768
rect 300912 342728 300918 342740
rect 301498 342728 301504 342740
rect 301556 342728 301562 342780
rect 175182 342252 175188 342304
rect 175240 342292 175246 342304
rect 176654 342292 176660 342304
rect 175240 342264 176660 342292
rect 175240 342252 175246 342264
rect 176654 342252 176660 342264
rect 176712 342252 176718 342304
rect 124122 340892 124128 340944
rect 124180 340932 124186 340944
rect 176654 340932 176660 340944
rect 124180 340904 176660 340932
rect 124180 340892 124186 340904
rect 176654 340892 176660 340904
rect 176712 340892 176718 340944
rect 295334 339464 295340 339516
rect 295392 339504 295398 339516
rect 308490 339504 308496 339516
rect 295392 339476 308496 339504
rect 295392 339464 295398 339476
rect 308490 339464 308496 339476
rect 308548 339464 308554 339516
rect 90358 335996 90364 336048
rect 90416 336036 90422 336048
rect 98638 336036 98644 336048
rect 90416 336008 98644 336036
rect 90416 335996 90422 336008
rect 98638 335996 98644 336008
rect 98696 335996 98702 336048
rect 161566 334568 161572 334620
rect 161624 334608 161630 334620
rect 177942 334608 177948 334620
rect 161624 334580 177948 334608
rect 161624 334568 161630 334580
rect 177942 334568 177948 334580
rect 178000 334568 178006 334620
rect 104158 332596 104164 332648
rect 104216 332636 104222 332648
rect 176654 332636 176660 332648
rect 104216 332608 176660 332636
rect 104216 332596 104222 332608
rect 176654 332596 176660 332608
rect 176712 332596 176718 332648
rect 106274 330488 106280 330540
rect 106332 330528 106338 330540
rect 161566 330528 161572 330540
rect 106332 330500 161572 330528
rect 106332 330488 106338 330500
rect 161566 330488 161572 330500
rect 161624 330488 161630 330540
rect 374638 330488 374644 330540
rect 374696 330528 374702 330540
rect 412634 330528 412640 330540
rect 374696 330500 412640 330528
rect 374696 330488 374702 330500
rect 412634 330488 412640 330500
rect 412692 330488 412698 330540
rect 294414 327088 294420 327140
rect 294472 327128 294478 327140
rect 311158 327128 311164 327140
rect 294472 327100 311164 327128
rect 294472 327088 294478 327100
rect 311158 327088 311164 327100
rect 311216 327088 311222 327140
rect 130562 325660 130568 325712
rect 130620 325700 130626 325712
rect 179506 325700 179512 325712
rect 130620 325672 179512 325700
rect 130620 325660 130626 325672
rect 179506 325660 179512 325672
rect 179564 325660 179570 325712
rect 355318 324300 355324 324352
rect 355376 324340 355382 324352
rect 580166 324340 580172 324352
rect 355376 324312 580172 324340
rect 355376 324300 355382 324312
rect 580166 324300 580172 324312
rect 580224 324300 580230 324352
rect 173802 321580 173808 321632
rect 173860 321620 173866 321632
rect 176654 321620 176660 321632
rect 173860 321592 176660 321620
rect 173860 321580 173866 321592
rect 176654 321580 176660 321592
rect 176712 321580 176718 321632
rect 3418 320832 3424 320884
rect 3476 320872 3482 320884
rect 120074 320872 120080 320884
rect 3476 320844 120080 320872
rect 3476 320832 3482 320844
rect 120074 320832 120080 320844
rect 120132 320832 120138 320884
rect 295518 320152 295524 320204
rect 295576 320192 295582 320204
rect 305638 320192 305644 320204
rect 295576 320164 305644 320192
rect 295576 320152 295582 320164
rect 305638 320152 305644 320164
rect 305696 320152 305702 320204
rect 3418 318792 3424 318844
rect 3476 318832 3482 318844
rect 100018 318832 100024 318844
rect 3476 318804 100024 318832
rect 3476 318792 3482 318804
rect 100018 318792 100024 318804
rect 100076 318792 100082 318844
rect 295518 318792 295524 318844
rect 295576 318832 295582 318844
rect 350534 318832 350540 318844
rect 295576 318804 350540 318832
rect 295576 318792 295582 318804
rect 350534 318792 350540 318804
rect 350592 318792 350598 318844
rect 295610 316684 295616 316736
rect 295668 316724 295674 316736
rect 468478 316724 468484 316736
rect 295668 316696 468484 316724
rect 295668 316684 295674 316696
rect 468478 316684 468484 316696
rect 468536 316684 468542 316736
rect 166258 314644 166264 314696
rect 166316 314684 166322 314696
rect 176654 314684 176660 314696
rect 166316 314656 176660 314684
rect 166316 314644 166322 314656
rect 176654 314644 176660 314656
rect 176712 314644 176718 314696
rect 295518 314576 295524 314628
rect 295576 314616 295582 314628
rect 299474 314616 299480 314628
rect 295576 314588 299480 314616
rect 295576 314576 295582 314588
rect 299474 314576 299480 314588
rect 299532 314576 299538 314628
rect 25498 313896 25504 313948
rect 25556 313936 25562 313948
rect 119614 313936 119620 313948
rect 25556 313908 119620 313936
rect 25556 313896 25562 313908
rect 119614 313896 119620 313908
rect 119672 313896 119678 313948
rect 299474 313896 299480 313948
rect 299532 313936 299538 313948
rect 418798 313936 418804 313948
rect 299532 313908 418804 313936
rect 299532 313896 299538 313908
rect 418798 313896 418804 313908
rect 418856 313896 418862 313948
rect 116578 312740 116584 312792
rect 116636 312780 116642 312792
rect 121454 312780 121460 312792
rect 116636 312752 121460 312780
rect 116636 312740 116642 312752
rect 121454 312740 121460 312752
rect 121512 312740 121518 312792
rect 8938 312536 8944 312588
rect 8996 312576 9002 312588
rect 94498 312576 94504 312588
rect 8996 312548 94504 312576
rect 8996 312536 9002 312548
rect 94498 312536 94504 312548
rect 94556 312536 94562 312588
rect 302234 312536 302240 312588
rect 302292 312576 302298 312588
rect 309778 312576 309784 312588
rect 302292 312548 309784 312576
rect 302292 312536 302298 312548
rect 309778 312536 309784 312548
rect 309836 312536 309842 312588
rect 129182 311924 129188 311976
rect 129240 311964 129246 311976
rect 166258 311964 166264 311976
rect 129240 311936 166264 311964
rect 129240 311924 129246 311936
rect 166258 311924 166264 311936
rect 166316 311924 166322 311976
rect 138106 311856 138112 311908
rect 138164 311896 138170 311908
rect 178954 311896 178960 311908
rect 138164 311868 178960 311896
rect 138164 311856 138170 311868
rect 178954 311856 178960 311868
rect 179012 311856 179018 311908
rect 295518 311856 295524 311908
rect 295576 311896 295582 311908
rect 302234 311896 302240 311908
rect 295576 311868 302240 311896
rect 295576 311856 295582 311868
rect 302234 311856 302240 311868
rect 302292 311856 302298 311908
rect 4798 311108 4804 311160
rect 4856 311148 4862 311160
rect 121546 311148 121552 311160
rect 4856 311120 121552 311148
rect 4856 311108 4862 311120
rect 121546 311108 121552 311120
rect 121604 311108 121610 311160
rect 295518 309748 295524 309800
rect 295576 309788 295582 309800
rect 298186 309788 298192 309800
rect 295576 309760 298192 309788
rect 295576 309748 295582 309760
rect 298186 309748 298192 309760
rect 298244 309788 298250 309800
rect 471238 309788 471244 309800
rect 298244 309760 471244 309788
rect 298244 309748 298250 309760
rect 471238 309748 471244 309760
rect 471296 309748 471302 309800
rect 173158 309136 173164 309188
rect 173216 309176 173222 309188
rect 176654 309176 176660 309188
rect 173216 309148 176660 309176
rect 173216 309136 173222 309148
rect 176654 309136 176660 309148
rect 176712 309136 176718 309188
rect 158530 307844 158536 307896
rect 158588 307884 158594 307896
rect 176654 307884 176660 307896
rect 158588 307856 176660 307884
rect 158588 307844 158594 307856
rect 176654 307844 176660 307856
rect 176712 307844 176718 307896
rect 82170 307776 82176 307828
rect 82228 307816 82234 307828
rect 164970 307816 164976 307828
rect 82228 307788 164976 307816
rect 82228 307776 82234 307788
rect 164970 307776 164976 307788
rect 165028 307776 165034 307828
rect 295518 307776 295524 307828
rect 295576 307816 295582 307828
rect 303706 307816 303712 307828
rect 295576 307788 303712 307816
rect 295576 307776 295582 307788
rect 303706 307776 303712 307788
rect 303764 307776 303770 307828
rect 91094 307028 91100 307080
rect 91152 307068 91158 307080
rect 138106 307068 138112 307080
rect 91152 307040 138112 307068
rect 91152 307028 91158 307040
rect 138106 307028 138112 307040
rect 138164 307028 138170 307080
rect 85574 306348 85580 306400
rect 85632 306388 85638 306400
rect 140222 306388 140228 306400
rect 85632 306360 140228 306388
rect 85632 306348 85638 306360
rect 140222 306348 140228 306360
rect 140280 306348 140286 306400
rect 314654 305600 314660 305652
rect 314712 305640 314718 305652
rect 347038 305640 347044 305652
rect 314712 305612 347044 305640
rect 314712 305600 314718 305612
rect 347038 305600 347044 305612
rect 347096 305600 347102 305652
rect 75362 305056 75368 305108
rect 75420 305096 75426 305108
rect 147030 305096 147036 305108
rect 75420 305068 147036 305096
rect 75420 305056 75426 305068
rect 147030 305056 147036 305068
rect 147088 305056 147094 305108
rect 3234 304988 3240 305040
rect 3292 305028 3298 305040
rect 120166 305028 120172 305040
rect 3292 305000 120172 305028
rect 3292 304988 3298 305000
rect 120166 304988 120172 305000
rect 120224 305028 120230 305040
rect 176654 305028 176660 305040
rect 120224 305000 176660 305028
rect 120224 304988 120230 305000
rect 176654 304988 176660 305000
rect 176712 304988 176718 305040
rect 295426 304988 295432 305040
rect 295484 305028 295490 305040
rect 314654 305028 314660 305040
rect 295484 305000 314660 305028
rect 295484 304988 295490 305000
rect 314654 304988 314660 305000
rect 314712 304988 314718 305040
rect 32398 304920 32404 304972
rect 32456 304960 32462 304972
rect 72234 304960 72240 304972
rect 32456 304932 72240 304960
rect 32456 304920 32462 304932
rect 72234 304920 72240 304932
rect 72292 304920 72298 304972
rect 82078 304240 82084 304292
rect 82136 304280 82142 304292
rect 115842 304280 115848 304292
rect 82136 304252 115848 304280
rect 82136 304240 82142 304252
rect 115842 304240 115848 304252
rect 115900 304240 115906 304292
rect 98730 303696 98736 303748
rect 98788 303736 98794 303748
rect 149698 303736 149704 303748
rect 98788 303708 149704 303736
rect 98788 303696 98794 303708
rect 149698 303696 149704 303708
rect 149756 303696 149762 303748
rect 94590 303628 94596 303680
rect 94648 303668 94654 303680
rect 146938 303668 146944 303680
rect 94648 303640 146944 303668
rect 94648 303628 94654 303640
rect 146938 303628 146944 303640
rect 146996 303628 147002 303680
rect 88334 303560 88340 303612
rect 88392 303600 88398 303612
rect 104158 303600 104164 303612
rect 88392 303572 104164 303600
rect 88392 303560 88398 303572
rect 104158 303560 104164 303572
rect 104216 303600 104222 303612
rect 104434 303600 104440 303612
rect 104216 303572 104440 303600
rect 104216 303560 104222 303572
rect 104434 303560 104440 303572
rect 104492 303560 104498 303612
rect 294230 303560 294236 303612
rect 294288 303600 294294 303612
rect 374638 303600 374644 303612
rect 294288 303572 374644 303600
rect 294288 303560 294294 303572
rect 374638 303560 374644 303572
rect 374696 303560 374702 303612
rect 43438 302880 43444 302932
rect 43496 302920 43502 302932
rect 84378 302920 84384 302932
rect 43496 302892 84384 302920
rect 43496 302880 43502 302892
rect 84378 302880 84384 302892
rect 84436 302880 84442 302932
rect 89714 302268 89720 302320
rect 89772 302308 89778 302320
rect 163590 302308 163596 302320
rect 89772 302280 163596 302308
rect 89772 302268 89778 302280
rect 163590 302268 163596 302280
rect 163648 302268 163654 302320
rect 74534 302200 74540 302252
rect 74592 302240 74598 302252
rect 162210 302240 162216 302252
rect 74592 302212 162216 302240
rect 74592 302200 74598 302212
rect 162210 302200 162216 302212
rect 162268 302200 162274 302252
rect 114738 302132 114744 302184
rect 114796 302172 114802 302184
rect 115842 302172 115848 302184
rect 114796 302144 115848 302172
rect 114796 302132 114802 302144
rect 115842 302132 115848 302144
rect 115900 302172 115906 302184
rect 173158 302172 173164 302184
rect 115900 302144 173164 302172
rect 115900 302132 115906 302144
rect 173158 302132 173164 302144
rect 173216 302132 173222 302184
rect 100018 301452 100024 301504
rect 100076 301492 100082 301504
rect 116578 301492 116584 301504
rect 100076 301464 116584 301492
rect 100076 301452 100082 301464
rect 116578 301452 116584 301464
rect 116636 301452 116642 301504
rect 106918 301044 106924 301096
rect 106976 301084 106982 301096
rect 133138 301084 133144 301096
rect 106976 301056 133144 301084
rect 106976 301044 106982 301056
rect 133138 301044 133144 301056
rect 133196 301044 133202 301096
rect 103698 300976 103704 301028
rect 103756 301016 103762 301028
rect 143074 301016 143080 301028
rect 103756 300988 143080 301016
rect 103756 300976 103762 300988
rect 143074 300976 143080 300988
rect 143132 300976 143138 301028
rect 90266 300908 90272 300960
rect 90324 300948 90330 300960
rect 142890 300948 142896 300960
rect 90324 300920 142896 300948
rect 90324 300908 90330 300920
rect 142890 300908 142896 300920
rect 142948 300908 142954 300960
rect 7558 300840 7564 300892
rect 7616 300880 7622 300892
rect 117958 300880 117964 300892
rect 7616 300852 117964 300880
rect 7616 300840 7622 300852
rect 117958 300840 117964 300852
rect 118016 300840 118022 300892
rect 160002 300772 160008 300824
rect 160060 300812 160066 300824
rect 160830 300812 160836 300824
rect 160060 300784 160836 300812
rect 160060 300772 160066 300784
rect 160830 300772 160836 300784
rect 160888 300772 160894 300824
rect 39942 300092 39948 300144
rect 40000 300132 40006 300144
rect 70946 300132 70952 300144
rect 40000 300104 70952 300132
rect 40000 300092 40006 300104
rect 70946 300092 70952 300104
rect 71004 300092 71010 300144
rect 99374 299820 99380 299872
rect 99432 299860 99438 299872
rect 124950 299860 124956 299872
rect 99432 299832 124956 299860
rect 99432 299820 99438 299832
rect 124950 299820 124956 299832
rect 125008 299820 125014 299872
rect 92842 299752 92848 299804
rect 92900 299792 92906 299804
rect 130470 299792 130476 299804
rect 92900 299764 130476 299792
rect 92900 299752 92906 299764
rect 130470 299752 130476 299764
rect 130528 299752 130534 299804
rect 109126 299684 109132 299736
rect 109184 299724 109190 299736
rect 153930 299724 153936 299736
rect 109184 299696 153936 299724
rect 109184 299684 109190 299696
rect 153930 299684 153936 299696
rect 153988 299684 153994 299736
rect 85666 299616 85672 299668
rect 85724 299656 85730 299668
rect 137278 299656 137284 299668
rect 85724 299628 137284 299656
rect 85724 299616 85730 299628
rect 137278 299616 137284 299628
rect 137336 299616 137342 299668
rect 81434 299548 81440 299600
rect 81492 299588 81498 299600
rect 157978 299588 157984 299600
rect 81492 299560 157984 299588
rect 81492 299548 81498 299560
rect 157978 299548 157984 299560
rect 158036 299548 158042 299600
rect 66162 299480 66168 299532
rect 66220 299520 66226 299532
rect 160002 299520 160008 299532
rect 66220 299492 160008 299520
rect 66220 299480 66226 299492
rect 160002 299480 160008 299492
rect 160060 299480 160066 299532
rect 166442 299412 166448 299464
rect 166500 299452 166506 299464
rect 166902 299452 166908 299464
rect 166500 299424 166908 299452
rect 166500 299412 166506 299424
rect 166902 299412 166908 299424
rect 166960 299452 166966 299464
rect 176654 299452 176660 299464
rect 166960 299424 176660 299452
rect 166960 299412 166966 299424
rect 176654 299412 176660 299424
rect 176712 299412 176718 299464
rect 297450 299412 297456 299464
rect 297508 299452 297514 299464
rect 579614 299452 579620 299464
rect 297508 299424 579620 299452
rect 297508 299412 297514 299424
rect 579614 299412 579620 299424
rect 579672 299412 579678 299464
rect 102226 298392 102232 298444
rect 102284 298432 102290 298444
rect 145650 298432 145656 298444
rect 102284 298404 145656 298432
rect 102284 298392 102290 298404
rect 145650 298392 145656 298404
rect 145708 298392 145714 298444
rect 106734 298324 106740 298376
rect 106792 298364 106798 298376
rect 151078 298364 151084 298376
rect 106792 298336 151084 298364
rect 106792 298324 106798 298336
rect 151078 298324 151084 298336
rect 151136 298324 151142 298376
rect 88058 298256 88064 298308
rect 88116 298296 88122 298308
rect 133230 298296 133236 298308
rect 88116 298268 133236 298296
rect 88116 298256 88122 298268
rect 133230 298256 133236 298268
rect 133288 298256 133294 298308
rect 88702 298188 88708 298240
rect 88760 298228 88766 298240
rect 135898 298228 135904 298240
rect 88760 298200 135904 298228
rect 88760 298188 88766 298200
rect 135898 298188 135904 298200
rect 135956 298188 135962 298240
rect 67542 298120 67548 298172
rect 67600 298160 67606 298172
rect 151262 298160 151268 298172
rect 67600 298132 151268 298160
rect 67600 298120 67606 298132
rect 151262 298120 151268 298132
rect 151320 298120 151326 298172
rect 157334 298052 157340 298104
rect 157392 298092 157398 298104
rect 158622 298092 158628 298104
rect 157392 298064 158628 298092
rect 157392 298052 157398 298064
rect 158622 298052 158628 298064
rect 158680 298092 158686 298104
rect 176654 298092 176660 298104
rect 158680 298064 176660 298092
rect 158680 298052 158686 298064
rect 176654 298052 176660 298064
rect 176712 298052 176718 298104
rect 84194 297032 84200 297084
rect 84252 297072 84258 297084
rect 153838 297072 153844 297084
rect 84252 297044 153844 297072
rect 84252 297032 84258 297044
rect 153838 297032 153844 297044
rect 153896 297032 153902 297084
rect 99006 296964 99012 297016
rect 99064 297004 99070 297016
rect 123478 297004 123484 297016
rect 99064 296976 123484 297004
rect 99064 296964 99070 296976
rect 123478 296964 123484 296976
rect 123536 296964 123542 297016
rect 94498 296896 94504 296948
rect 94556 296936 94562 296948
rect 144362 296936 144368 296948
rect 94556 296908 144368 296936
rect 94556 296896 94562 296908
rect 144362 296896 144368 296908
rect 144420 296896 144426 296948
rect 75178 296828 75184 296880
rect 75236 296868 75242 296880
rect 134610 296868 134616 296880
rect 75236 296840 134616 296868
rect 75236 296828 75242 296840
rect 134610 296828 134616 296840
rect 134668 296828 134674 296880
rect 31018 296760 31024 296812
rect 31076 296800 31082 296812
rect 97074 296800 97080 296812
rect 31076 296772 97080 296800
rect 31076 296760 31082 296772
rect 97074 296760 97080 296772
rect 97132 296760 97138 296812
rect 111242 296760 111248 296812
rect 111300 296800 111306 296812
rect 159358 296800 159364 296812
rect 111300 296772 159364 296800
rect 111300 296760 111306 296772
rect 159358 296760 159364 296772
rect 159416 296760 159422 296812
rect 113818 296692 113824 296744
rect 113876 296732 113882 296744
rect 120718 296732 120724 296744
rect 113876 296704 120724 296732
rect 113876 296692 113882 296704
rect 120718 296692 120724 296704
rect 120776 296692 120782 296744
rect 97718 295672 97724 295724
rect 97776 295712 97782 295724
rect 128998 295712 129004 295724
rect 97776 295684 129004 295712
rect 97776 295672 97782 295684
rect 128998 295672 129004 295684
rect 129056 295672 129062 295724
rect 83550 295604 83556 295656
rect 83608 295644 83614 295656
rect 126330 295644 126336 295656
rect 83608 295616 126336 295644
rect 83608 295604 83614 295616
rect 126330 295604 126336 295616
rect 126388 295604 126394 295656
rect 82262 295536 82268 295588
rect 82320 295576 82326 295588
rect 138750 295576 138756 295588
rect 82320 295548 138756 295576
rect 82320 295536 82326 295548
rect 138750 295536 138756 295548
rect 138808 295536 138814 295588
rect 68554 295468 68560 295520
rect 68612 295508 68618 295520
rect 129274 295508 129280 295520
rect 68612 295480 129280 295508
rect 68612 295468 68618 295480
rect 129274 295468 129280 295480
rect 129332 295468 129338 295520
rect 14458 295400 14464 295452
rect 14516 295440 14522 295452
rect 92566 295440 92572 295452
rect 14516 295412 92572 295440
rect 14516 295400 14522 295412
rect 92566 295400 92572 295412
rect 92624 295440 92630 295452
rect 167730 295440 167736 295452
rect 92624 295412 167736 295440
rect 92624 295400 92630 295412
rect 167730 295400 167736 295412
rect 167788 295400 167794 295452
rect 67266 295332 67272 295384
rect 67324 295372 67330 295384
rect 147122 295372 147128 295384
rect 67324 295344 147128 295372
rect 67324 295332 67330 295344
rect 147122 295332 147128 295344
rect 147180 295332 147186 295384
rect 295426 295332 295432 295384
rect 295484 295372 295490 295384
rect 309870 295372 309876 295384
rect 295484 295344 309876 295372
rect 295484 295332 295490 295344
rect 309870 295332 309876 295344
rect 309928 295332 309934 295384
rect 73246 294720 73252 294772
rect 73304 294760 73310 294772
rect 82170 294760 82176 294772
rect 73304 294732 82176 294760
rect 73304 294720 73310 294732
rect 82170 294720 82176 294732
rect 82228 294720 82234 294772
rect 79686 294652 79692 294704
rect 79744 294692 79750 294704
rect 94590 294692 94596 294704
rect 79744 294664 94596 294692
rect 79744 294652 79750 294664
rect 94590 294652 94596 294664
rect 94648 294652 94654 294704
rect 71958 294584 71964 294636
rect 72016 294624 72022 294636
rect 106918 294624 106924 294636
rect 72016 294596 106924 294624
rect 72016 294584 72022 294596
rect 106918 294584 106924 294596
rect 106976 294584 106982 294636
rect 111886 294312 111892 294364
rect 111944 294352 111950 294364
rect 126422 294352 126428 294364
rect 111944 294324 126428 294352
rect 111944 294312 111950 294324
rect 126422 294312 126428 294324
rect 126480 294312 126486 294364
rect 91922 294244 91928 294296
rect 91980 294284 91986 294296
rect 131758 294284 131764 294296
rect 91980 294256 131764 294284
rect 91980 294244 91986 294256
rect 131758 294244 131764 294256
rect 131816 294244 131822 294296
rect 80974 294176 80980 294228
rect 81032 294216 81038 294228
rect 125042 294216 125048 294228
rect 81032 294188 125048 294216
rect 81032 294176 81038 294188
rect 125042 294176 125048 294188
rect 125100 294176 125106 294228
rect 78582 294108 78588 294160
rect 78640 294148 78646 294160
rect 101398 294148 101404 294160
rect 78640 294120 101404 294148
rect 78640 294108 78646 294120
rect 101398 294108 101404 294120
rect 101456 294108 101462 294160
rect 105446 294108 105452 294160
rect 105504 294148 105510 294160
rect 152458 294148 152464 294160
rect 105504 294120 152464 294148
rect 105504 294108 105510 294120
rect 152458 294108 152464 294120
rect 152516 294108 152522 294160
rect 65610 294040 65616 294092
rect 65668 294080 65674 294092
rect 79318 294080 79324 294092
rect 65668 294052 79324 294080
rect 65668 294040 65674 294052
rect 79318 294040 79324 294052
rect 79376 294040 79382 294092
rect 93854 294040 93860 294092
rect 93912 294080 93918 294092
rect 115842 294080 115848 294092
rect 93912 294052 115848 294080
rect 93912 294040 93918 294052
rect 115842 294040 115848 294052
rect 115900 294040 115906 294092
rect 116578 294040 116584 294092
rect 116636 294080 116642 294092
rect 172054 294080 172060 294092
rect 116636 294052 172060 294080
rect 116636 294040 116642 294052
rect 172054 294040 172060 294052
rect 172112 294040 172118 294092
rect 75914 293972 75920 294024
rect 75972 294012 75978 294024
rect 76742 294012 76748 294024
rect 75972 293984 76748 294012
rect 75972 293972 75978 293984
rect 76742 293972 76748 293984
rect 76800 293972 76806 294024
rect 82906 293972 82912 294024
rect 82964 294012 82970 294024
rect 148410 294012 148416 294024
rect 82964 293984 148416 294012
rect 82964 293972 82970 293984
rect 148410 293972 148416 293984
rect 148468 293972 148474 294024
rect 158622 293972 158628 294024
rect 158680 294012 158686 294024
rect 176654 294012 176660 294024
rect 158680 293984 176660 294012
rect 158680 293972 158686 293984
rect 176654 293972 176660 293984
rect 176712 293972 176718 294024
rect 295334 293972 295340 294024
rect 295392 294012 295398 294024
rect 306374 294012 306380 294024
rect 295392 293984 306380 294012
rect 295392 293972 295398 293984
rect 306374 293972 306380 293984
rect 306432 293972 306438 294024
rect 84286 293904 84292 293956
rect 84344 293944 84350 293956
rect 85206 293944 85212 293956
rect 84344 293916 85212 293944
rect 84344 293904 84350 293916
rect 85206 293904 85212 293916
rect 85264 293904 85270 293956
rect 85574 293904 85580 293956
rect 85632 293944 85638 293956
rect 86494 293944 86500 293956
rect 85632 293916 86500 293944
rect 85632 293904 85638 293916
rect 86494 293904 86500 293916
rect 86552 293904 86558 293956
rect 109034 293904 109040 293956
rect 109092 293944 109098 293956
rect 109678 293944 109684 293956
rect 109092 293916 109684 293944
rect 109092 293904 109098 293916
rect 109678 293904 109684 293916
rect 109736 293904 109742 293956
rect 114554 293904 114560 293956
rect 114612 293944 114618 293956
rect 115382 293944 115388 293956
rect 114612 293916 115388 293944
rect 114612 293904 114618 293916
rect 115382 293904 115388 293916
rect 115440 293904 115446 293956
rect 3418 293224 3424 293276
rect 3476 293264 3482 293276
rect 78582 293264 78588 293276
rect 3476 293236 78588 293264
rect 3476 293224 3482 293236
rect 78582 293224 78588 293236
rect 78640 293224 78646 293276
rect 87414 293224 87420 293276
rect 87472 293264 87478 293276
rect 98730 293264 98736 293276
rect 87472 293236 98736 293264
rect 87472 293224 87478 293236
rect 98730 293224 98736 293236
rect 98788 293224 98794 293276
rect 115842 293224 115848 293276
rect 115900 293264 115906 293276
rect 140038 293264 140044 293276
rect 115900 293236 140044 293264
rect 115900 293224 115906 293236
rect 140038 293224 140044 293236
rect 140096 293224 140102 293276
rect 3326 292816 3332 292868
rect 3384 292856 3390 292868
rect 8938 292856 8944 292868
rect 3384 292828 8944 292856
rect 3384 292816 3390 292828
rect 8938 292816 8944 292828
rect 8996 292816 9002 292868
rect 112530 292816 112536 292868
rect 112588 292856 112594 292868
rect 141418 292856 141424 292868
rect 112588 292828 141424 292856
rect 112588 292816 112594 292828
rect 141418 292816 141424 292828
rect 141476 292816 141482 292868
rect 102870 292748 102876 292800
rect 102928 292788 102934 292800
rect 134702 292788 134708 292800
rect 102928 292760 134708 292788
rect 102928 292748 102934 292760
rect 134702 292748 134708 292760
rect 134760 292748 134766 292800
rect 117038 292680 117044 292732
rect 117096 292720 117102 292732
rect 166258 292720 166264 292732
rect 117096 292692 166264 292720
rect 117096 292680 117102 292692
rect 166258 292680 166264 292692
rect 166316 292680 166322 292732
rect 68830 292612 68836 292664
rect 68888 292652 68894 292664
rect 123662 292652 123668 292664
rect 68888 292624 123668 292652
rect 68888 292612 68894 292624
rect 123662 292612 123668 292624
rect 123720 292612 123726 292664
rect 67358 292544 67364 292596
rect 67416 292584 67422 292596
rect 70670 292584 70676 292596
rect 67416 292556 70676 292584
rect 67416 292544 67422 292556
rect 70670 292544 70676 292556
rect 70728 292544 70734 292596
rect 98638 292544 98644 292596
rect 98696 292584 98702 292596
rect 170490 292584 170496 292596
rect 98696 292556 170496 292584
rect 98696 292544 98702 292556
rect 170490 292544 170496 292556
rect 170548 292544 170554 292596
rect 71682 292476 71688 292528
rect 71740 292516 71746 292528
rect 111150 292516 111156 292528
rect 71740 292488 111156 292516
rect 71740 292476 71746 292488
rect 111150 292476 111156 292488
rect 111208 292476 111214 292528
rect 121546 292476 121552 292528
rect 121604 292516 121610 292528
rect 175918 292516 175924 292528
rect 121604 292488 175924 292516
rect 121604 292476 121610 292488
rect 175918 292476 175924 292488
rect 175976 292476 175982 292528
rect 103486 291944 103744 291972
rect 101306 291864 101312 291916
rect 101364 291904 101370 291916
rect 103486 291904 103514 291944
rect 101364 291876 103514 291904
rect 101364 291864 101370 291876
rect 103606 291864 103612 291916
rect 103664 291864 103670 291916
rect 67450 291184 67456 291236
rect 67508 291224 67514 291236
rect 69750 291224 69756 291236
rect 67508 291196 69756 291224
rect 67508 291184 67514 291196
rect 69750 291184 69756 291196
rect 69808 291184 69814 291236
rect 103624 291224 103652 291864
rect 103716 291360 103744 291944
rect 110874 291864 110880 291916
rect 110932 291904 110938 291916
rect 110932 291876 113174 291904
rect 110932 291864 110938 291876
rect 113146 291428 113174 291876
rect 119338 291864 119344 291916
rect 119396 291904 119402 291916
rect 119706 291904 119712 291916
rect 119396 291876 119712 291904
rect 119396 291864 119402 291876
rect 119706 291864 119712 291876
rect 119764 291864 119770 291916
rect 135990 291428 135996 291440
rect 113146 291400 135996 291428
rect 135990 291388 135996 291400
rect 136048 291388 136054 291440
rect 127618 291360 127624 291372
rect 103716 291332 127624 291360
rect 127618 291320 127624 291332
rect 127676 291320 127682 291372
rect 119798 291252 119804 291304
rect 119856 291292 119862 291304
rect 152642 291292 152648 291304
rect 119856 291264 152648 291292
rect 119856 291252 119862 291264
rect 152642 291252 152648 291264
rect 152700 291252 152706 291304
rect 156598 291224 156604 291236
rect 103624 291196 156604 291224
rect 156598 291184 156604 291196
rect 156656 291184 156662 291236
rect 168282 291184 168288 291236
rect 168340 291224 168346 291236
rect 176654 291224 176660 291236
rect 168340 291196 176660 291224
rect 168340 291184 168346 291196
rect 176654 291184 176660 291196
rect 176712 291184 176718 291236
rect 26878 290436 26884 290488
rect 26936 290476 26942 290488
rect 67726 290476 67732 290488
rect 26936 290448 67732 290476
rect 26936 290436 26942 290448
rect 67726 290436 67732 290448
rect 67784 290436 67790 290488
rect 302326 290436 302332 290488
rect 302384 290476 302390 290488
rect 400858 290476 400864 290488
rect 302384 290448 400864 290476
rect 302384 290436 302390 290448
rect 400858 290436 400864 290448
rect 400916 290436 400922 290488
rect 121638 289960 121644 290012
rect 121696 290000 121702 290012
rect 138658 290000 138664 290012
rect 121696 289972 138664 290000
rect 121696 289960 121702 289972
rect 138658 289960 138664 289972
rect 138716 289960 138722 290012
rect 121546 289892 121552 289944
rect 121604 289932 121610 289944
rect 144270 289932 144276 289944
rect 121604 289904 144276 289932
rect 121604 289892 121610 289904
rect 144270 289892 144276 289904
rect 144328 289892 144334 289944
rect 53650 289824 53656 289876
rect 53708 289864 53714 289876
rect 67634 289864 67640 289876
rect 53708 289836 67640 289864
rect 53708 289824 53714 289836
rect 67634 289824 67640 289836
rect 67692 289824 67698 289876
rect 120810 289824 120816 289876
rect 120868 289864 120874 289876
rect 176654 289864 176660 289876
rect 120868 289836 176660 289864
rect 120868 289824 120874 289836
rect 176654 289824 176660 289836
rect 176712 289824 176718 289876
rect 295518 289824 295524 289876
rect 295576 289864 295582 289876
rect 302326 289864 302332 289876
rect 295576 289836 302332 289864
rect 295576 289824 295582 289836
rect 302326 289824 302332 289836
rect 302384 289824 302390 289876
rect 121546 289756 121552 289808
rect 121604 289796 121610 289808
rect 174538 289796 174544 289808
rect 121604 289768 174544 289796
rect 121604 289756 121610 289768
rect 174538 289756 174544 289768
rect 174596 289756 174602 289808
rect 67266 289280 67272 289332
rect 67324 289320 67330 289332
rect 67542 289320 67548 289332
rect 67324 289292 67548 289320
rect 67324 289280 67330 289292
rect 67542 289280 67548 289292
rect 67600 289280 67606 289332
rect 64782 288396 64788 288448
rect 64840 288436 64846 288448
rect 67634 288436 67640 288448
rect 64840 288408 67640 288436
rect 64840 288396 64846 288408
rect 67634 288396 67640 288408
rect 67692 288396 67698 288448
rect 121546 288396 121552 288448
rect 121604 288436 121610 288448
rect 148502 288436 148508 288448
rect 121604 288408 148508 288436
rect 121604 288396 121610 288408
rect 148502 288396 148508 288408
rect 148560 288396 148566 288448
rect 121638 288328 121644 288380
rect 121696 288368 121702 288380
rect 167638 288368 167644 288380
rect 121696 288340 167644 288368
rect 121696 288328 121702 288340
rect 167638 288328 167644 288340
rect 167696 288328 167702 288380
rect 3510 287648 3516 287700
rect 3568 287688 3574 287700
rect 65610 287688 65616 287700
rect 3568 287660 65616 287688
rect 3568 287648 3574 287660
rect 65610 287648 65616 287660
rect 65668 287648 65674 287700
rect 52362 287036 52368 287088
rect 52420 287076 52426 287088
rect 67634 287076 67640 287088
rect 52420 287048 67640 287076
rect 52420 287036 52426 287048
rect 67634 287036 67640 287048
rect 67692 287036 67698 287088
rect 121730 287036 121736 287088
rect 121788 287076 121794 287088
rect 145558 287076 145564 287088
rect 121788 287048 145564 287076
rect 121788 287036 121794 287048
rect 145558 287036 145564 287048
rect 145616 287036 145622 287088
rect 22738 286968 22744 287020
rect 22796 287008 22802 287020
rect 67542 287008 67548 287020
rect 22796 286980 67548 287008
rect 22796 286968 22802 286980
rect 67542 286968 67548 286980
rect 67600 286968 67606 287020
rect 121454 286424 121460 286476
rect 121512 286464 121518 286476
rect 124122 286464 124128 286476
rect 121512 286436 124128 286464
rect 121512 286424 121518 286436
rect 124122 286424 124128 286436
rect 124180 286464 124186 286476
rect 136082 286464 136088 286476
rect 124180 286436 136088 286464
rect 124180 286424 124186 286436
rect 136082 286424 136088 286436
rect 136140 286424 136146 286476
rect 122742 286356 122748 286408
rect 122800 286396 122806 286408
rect 171962 286396 171968 286408
rect 122800 286368 171968 286396
rect 122800 286356 122806 286368
rect 171962 286356 171968 286368
rect 172020 286356 172026 286408
rect 123570 286288 123576 286340
rect 123628 286328 123634 286340
rect 177850 286328 177856 286340
rect 123628 286300 177856 286328
rect 123628 286288 123634 286300
rect 177850 286288 177856 286300
rect 177908 286288 177914 286340
rect 60642 285744 60648 285796
rect 60700 285784 60706 285796
rect 67726 285784 67732 285796
rect 60700 285756 67732 285784
rect 60700 285744 60706 285756
rect 67726 285744 67732 285756
rect 67784 285744 67790 285796
rect 39942 285676 39948 285728
rect 40000 285716 40006 285728
rect 67634 285716 67640 285728
rect 40000 285688 67640 285716
rect 40000 285676 40006 285688
rect 67634 285676 67640 285688
rect 67692 285676 67698 285728
rect 295518 285676 295524 285728
rect 295576 285716 295582 285728
rect 309686 285716 309692 285728
rect 295576 285688 309692 285716
rect 295576 285676 295582 285688
rect 309686 285676 309692 285688
rect 309744 285676 309750 285728
rect 121546 285608 121552 285660
rect 121604 285648 121610 285660
rect 171870 285648 171876 285660
rect 121604 285620 171876 285648
rect 121604 285608 121610 285620
rect 171870 285608 171876 285620
rect 171928 285608 171934 285660
rect 121454 284316 121460 284368
rect 121512 284356 121518 284368
rect 167822 284356 167828 284368
rect 121512 284328 167828 284356
rect 121512 284316 121518 284328
rect 167822 284316 167828 284328
rect 167880 284316 167886 284368
rect 66162 284248 66168 284300
rect 66220 284288 66226 284300
rect 67634 284288 67640 284300
rect 66220 284260 67640 284288
rect 66220 284248 66226 284260
rect 67634 284248 67640 284260
rect 67692 284248 67698 284300
rect 310974 283568 310980 283620
rect 311032 283608 311038 283620
rect 355318 283608 355324 283620
rect 311032 283580 355324 283608
rect 311032 283568 311038 283580
rect 355318 283568 355324 283580
rect 355376 283568 355382 283620
rect 121454 282888 121460 282940
rect 121512 282928 121518 282940
rect 174538 282928 174544 282940
rect 121512 282900 174544 282928
rect 121512 282888 121518 282900
rect 174538 282888 174544 282900
rect 174596 282888 174602 282940
rect 295518 282888 295524 282940
rect 295576 282928 295582 282940
rect 310606 282928 310612 282940
rect 295576 282900 310612 282928
rect 295576 282888 295582 282900
rect 310606 282888 310612 282900
rect 310664 282928 310670 282940
rect 310974 282928 310980 282940
rect 310664 282900 310980 282928
rect 310664 282888 310670 282900
rect 310974 282888 310980 282900
rect 311032 282888 311038 282940
rect 64690 282820 64696 282872
rect 64748 282860 64754 282872
rect 67634 282860 67640 282872
rect 64748 282832 67640 282860
rect 64748 282820 64754 282832
rect 67634 282820 67640 282832
rect 67692 282820 67698 282872
rect 167730 282820 167736 282872
rect 167788 282860 167794 282872
rect 176654 282860 176660 282872
rect 167788 282832 176660 282860
rect 167788 282820 167794 282832
rect 176654 282820 176660 282832
rect 176712 282820 176718 282872
rect 121546 281596 121552 281648
rect 121604 281636 121610 281648
rect 164878 281636 164884 281648
rect 121604 281608 164884 281636
rect 121604 281596 121610 281608
rect 164878 281596 164884 281608
rect 164936 281596 164942 281648
rect 121454 281528 121460 281580
rect 121512 281568 121518 281580
rect 167638 281568 167644 281580
rect 121512 281540 167644 281568
rect 121512 281528 121518 281540
rect 167638 281528 167644 281540
rect 167696 281528 167702 281580
rect 295518 281528 295524 281580
rect 295576 281568 295582 281580
rect 353938 281568 353944 281580
rect 295576 281540 353944 281568
rect 295576 281528 295582 281540
rect 353938 281528 353944 281540
rect 353996 281528 354002 281580
rect 54938 280236 54944 280288
rect 54996 280276 55002 280288
rect 67634 280276 67640 280288
rect 54996 280248 67640 280276
rect 54996 280236 55002 280248
rect 67634 280236 67640 280248
rect 67692 280236 67698 280288
rect 121546 280236 121552 280288
rect 121604 280276 121610 280288
rect 137370 280276 137376 280288
rect 121604 280248 137376 280276
rect 121604 280236 121610 280248
rect 137370 280236 137376 280248
rect 137428 280236 137434 280288
rect 55122 280168 55128 280220
rect 55180 280208 55186 280220
rect 67726 280208 67732 280220
rect 55180 280180 67732 280208
rect 55180 280168 55186 280180
rect 67726 280168 67732 280180
rect 67784 280168 67790 280220
rect 121454 280168 121460 280220
rect 121512 280208 121518 280220
rect 156690 280208 156696 280220
rect 121512 280180 156696 280208
rect 121512 280168 121518 280180
rect 156690 280168 156696 280180
rect 156748 280168 156754 280220
rect 129274 280100 129280 280152
rect 129332 280140 129338 280152
rect 176746 280140 176752 280152
rect 129332 280112 176752 280140
rect 129332 280100 129338 280112
rect 176746 280100 176752 280112
rect 176804 280100 176810 280152
rect 48958 279420 48964 279472
rect 49016 279460 49022 279472
rect 67910 279460 67916 279472
rect 49016 279432 67916 279460
rect 49016 279420 49022 279432
rect 67910 279420 67916 279432
rect 67968 279420 67974 279472
rect 121454 278740 121460 278792
rect 121512 278780 121518 278792
rect 129090 278780 129096 278792
rect 121512 278752 129096 278780
rect 121512 278740 121518 278752
rect 129090 278740 129096 278752
rect 129148 278740 129154 278792
rect 295518 278740 295524 278792
rect 295576 278780 295582 278792
rect 299474 278780 299480 278792
rect 295576 278752 299480 278780
rect 295576 278740 295582 278752
rect 299474 278740 299480 278752
rect 299532 278740 299538 278792
rect 152458 278060 152464 278112
rect 152516 278100 152522 278112
rect 162670 278100 162676 278112
rect 152516 278072 162676 278100
rect 152516 278060 152522 278072
rect 162670 278060 162676 278072
rect 162728 278060 162734 278112
rect 121730 277992 121736 278044
rect 121788 278032 121794 278044
rect 167730 278032 167736 278044
rect 121788 278004 167736 278032
rect 121788 277992 121794 278004
rect 167730 277992 167736 278004
rect 167788 277992 167794 278044
rect 56502 277448 56508 277500
rect 56560 277488 56566 277500
rect 67634 277488 67640 277500
rect 56560 277460 67640 277488
rect 56560 277448 56566 277460
rect 67634 277448 67640 277460
rect 67692 277448 67698 277500
rect 46842 277380 46848 277432
rect 46900 277420 46906 277432
rect 67726 277420 67732 277432
rect 46900 277392 67732 277420
rect 46900 277380 46906 277392
rect 67726 277380 67732 277392
rect 67784 277380 67790 277432
rect 121454 277380 121460 277432
rect 121512 277420 121518 277432
rect 149882 277420 149888 277432
rect 121512 277392 149888 277420
rect 121512 277380 121518 277392
rect 149882 277380 149888 277392
rect 149940 277380 149946 277432
rect 162670 277380 162676 277432
rect 162728 277420 162734 277432
rect 176654 277420 176660 277432
rect 162728 277392 176660 277420
rect 162728 277380 162734 277392
rect 176654 277380 176660 277392
rect 176712 277380 176718 277432
rect 305086 276632 305092 276684
rect 305144 276672 305150 276684
rect 337378 276672 337384 276684
rect 305144 276644 337384 276672
rect 305144 276632 305150 276644
rect 337378 276632 337384 276644
rect 337436 276632 337442 276684
rect 64690 276088 64696 276140
rect 64748 276128 64754 276140
rect 67634 276128 67640 276140
rect 64748 276100 67640 276128
rect 64748 276088 64754 276100
rect 67634 276088 67640 276100
rect 67692 276088 67698 276140
rect 121546 276088 121552 276140
rect 121604 276128 121610 276140
rect 147214 276128 147220 276140
rect 121604 276100 147220 276128
rect 121604 276088 121610 276100
rect 147214 276088 147220 276100
rect 147272 276088 147278 276140
rect 53742 276020 53748 276072
rect 53800 276060 53806 276072
rect 67726 276060 67732 276072
rect 53800 276032 67732 276060
rect 53800 276020 53806 276032
rect 67726 276020 67732 276032
rect 67784 276020 67790 276072
rect 121454 276020 121460 276072
rect 121512 276060 121518 276072
rect 166534 276060 166540 276072
rect 121512 276032 166540 276060
rect 121512 276020 121518 276032
rect 166534 276020 166540 276032
rect 166592 276020 166598 276072
rect 295610 276020 295616 276072
rect 295668 276060 295674 276072
rect 305086 276060 305092 276072
rect 295668 276032 305092 276060
rect 295668 276020 295674 276032
rect 305086 276020 305092 276032
rect 305144 276020 305150 276072
rect 172054 275952 172060 276004
rect 172112 275992 172118 276004
rect 176654 275992 176660 276004
rect 172112 275964 176660 275992
rect 172112 275952 172118 275964
rect 176654 275952 176660 275964
rect 176712 275952 176718 276004
rect 121454 274728 121460 274780
rect 121512 274768 121518 274780
rect 151170 274768 151176 274780
rect 121512 274740 151176 274768
rect 121512 274728 121518 274740
rect 151170 274728 151176 274740
rect 151228 274728 151234 274780
rect 63402 274660 63408 274712
rect 63460 274700 63466 274712
rect 67634 274700 67640 274712
rect 63460 274672 67640 274700
rect 63460 274660 63466 274672
rect 67634 274660 67640 274672
rect 67692 274660 67698 274712
rect 121546 274660 121552 274712
rect 121604 274700 121610 274712
rect 155494 274700 155500 274712
rect 121604 274672 155500 274700
rect 121604 274660 121610 274672
rect 155494 274660 155500 274672
rect 155552 274660 155558 274712
rect 121454 274388 121460 274440
rect 121512 274428 121518 274440
rect 124858 274428 124864 274440
rect 121512 274400 124864 274428
rect 121512 274388 121518 274400
rect 124858 274388 124864 274400
rect 124916 274388 124922 274440
rect 18598 273912 18604 273964
rect 18656 273952 18662 273964
rect 57238 273952 57244 273964
rect 18656 273924 57244 273952
rect 18656 273912 18662 273924
rect 57238 273912 57244 273924
rect 57296 273912 57302 273964
rect 64598 273300 64604 273352
rect 64656 273340 64662 273352
rect 67634 273340 67640 273352
rect 64656 273312 67640 273340
rect 64656 273300 64662 273312
rect 67634 273300 67640 273312
rect 67692 273300 67698 273352
rect 57238 273232 57244 273284
rect 57296 273272 57302 273284
rect 57606 273272 57612 273284
rect 57296 273244 57612 273272
rect 57296 273232 57302 273244
rect 57606 273232 57612 273244
rect 57664 273272 57670 273284
rect 67726 273272 67732 273284
rect 57664 273244 67732 273272
rect 57664 273232 57670 273244
rect 67726 273232 67732 273244
rect 67784 273232 67790 273284
rect 121454 273232 121460 273284
rect 121512 273272 121518 273284
rect 143166 273272 143172 273284
rect 121512 273244 143172 273272
rect 121512 273232 121518 273244
rect 143166 273232 143172 273244
rect 143224 273232 143230 273284
rect 128354 273164 128360 273216
rect 128412 273204 128418 273216
rect 176654 273204 176660 273216
rect 128412 273176 176660 273204
rect 128412 273164 128418 273176
rect 176654 273164 176660 273176
rect 176712 273164 176718 273216
rect 120902 272484 120908 272536
rect 120960 272524 120966 272536
rect 128354 272524 128360 272536
rect 120960 272496 128360 272524
rect 120960 272484 120966 272496
rect 128354 272484 128360 272496
rect 128412 272484 128418 272536
rect 62022 271940 62028 271992
rect 62080 271980 62086 271992
rect 67726 271980 67732 271992
rect 62080 271952 67732 271980
rect 62080 271940 62086 271952
rect 67726 271940 67732 271952
rect 67784 271940 67790 271992
rect 45370 271872 45376 271924
rect 45428 271912 45434 271924
rect 67634 271912 67640 271924
rect 45428 271884 67640 271912
rect 45428 271872 45434 271884
rect 67634 271872 67640 271884
rect 67692 271872 67698 271924
rect 121454 271872 121460 271924
rect 121512 271912 121518 271924
rect 155218 271912 155224 271924
rect 121512 271884 155224 271912
rect 121512 271872 121518 271884
rect 155218 271872 155224 271884
rect 155276 271872 155282 271924
rect 295610 271872 295616 271924
rect 295668 271912 295674 271924
rect 300946 271912 300952 271924
rect 295668 271884 300952 271912
rect 295668 271872 295674 271884
rect 300946 271872 300952 271884
rect 301004 271872 301010 271924
rect 62298 271804 62304 271856
rect 62356 271844 62362 271856
rect 62758 271844 62764 271856
rect 62356 271816 62764 271844
rect 62356 271804 62362 271816
rect 62758 271804 62764 271816
rect 62816 271844 62822 271856
rect 67726 271844 67732 271856
rect 62816 271816 67732 271844
rect 62816 271804 62822 271816
rect 67726 271804 67732 271816
rect 67784 271804 67790 271856
rect 50982 270512 50988 270564
rect 51040 270552 51046 270564
rect 67634 270552 67640 270564
rect 51040 270524 67640 270552
rect 51040 270512 51046 270524
rect 67634 270512 67640 270524
rect 67692 270512 67698 270564
rect 121454 270512 121460 270564
rect 121512 270552 121518 270564
rect 138842 270552 138848 270564
rect 121512 270524 138848 270552
rect 121512 270512 121518 270524
rect 138842 270512 138848 270524
rect 138900 270512 138906 270564
rect 66070 269152 66076 269204
rect 66128 269192 66134 269204
rect 68186 269192 68192 269204
rect 66128 269164 68192 269192
rect 66128 269152 66134 269164
rect 68186 269152 68192 269164
rect 68244 269152 68250 269204
rect 121454 269152 121460 269204
rect 121512 269192 121518 269204
rect 145742 269192 145748 269204
rect 121512 269164 145748 269192
rect 121512 269152 121518 269164
rect 145742 269152 145748 269164
rect 145800 269152 145806 269204
rect 44082 269084 44088 269136
rect 44140 269124 44146 269136
rect 67634 269124 67640 269136
rect 44140 269096 67640 269124
rect 44140 269084 44146 269096
rect 67634 269084 67640 269096
rect 67692 269084 67698 269136
rect 121546 269084 121552 269136
rect 121604 269124 121610 269136
rect 165062 269124 165068 269136
rect 121604 269096 165068 269124
rect 121604 269084 121610 269096
rect 165062 269084 165068 269096
rect 165120 269084 165126 269136
rect 295610 269084 295616 269136
rect 295668 269124 295674 269136
rect 345658 269124 345664 269136
rect 295668 269096 345664 269124
rect 295668 269084 295674 269096
rect 345658 269084 345664 269096
rect 345716 269084 345722 269136
rect 66162 268200 66168 268252
rect 66220 268240 66226 268252
rect 68186 268240 68192 268252
rect 66220 268212 68192 268240
rect 66220 268200 66226 268212
rect 68186 268200 68192 268212
rect 68244 268200 68250 268252
rect 121454 267792 121460 267844
rect 121512 267832 121518 267844
rect 134794 267832 134800 267844
rect 121512 267804 134800 267832
rect 121512 267792 121518 267804
rect 134794 267792 134800 267804
rect 134852 267792 134858 267844
rect 161382 267792 161388 267844
rect 161440 267832 161446 267844
rect 176654 267832 176660 267844
rect 161440 267804 176660 267832
rect 161440 267792 161446 267804
rect 176654 267792 176660 267804
rect 176712 267792 176718 267844
rect 46750 267724 46756 267776
rect 46808 267764 46814 267776
rect 67634 267764 67640 267776
rect 46808 267736 67640 267764
rect 46808 267724 46814 267736
rect 67634 267724 67640 267736
rect 67692 267724 67698 267776
rect 120074 267724 120080 267776
rect 120132 267764 120138 267776
rect 163682 267764 163688 267776
rect 120132 267736 163688 267764
rect 120132 267724 120138 267736
rect 163682 267724 163688 267736
rect 163740 267724 163746 267776
rect 63218 266976 63224 267028
rect 63276 267016 63282 267028
rect 67634 267016 67640 267028
rect 63276 266988 67640 267016
rect 63276 266976 63282 266988
rect 67634 266976 67640 266988
rect 67692 266976 67698 267028
rect 121546 266432 121552 266484
rect 121604 266472 121610 266484
rect 152458 266472 152464 266484
rect 121604 266444 152464 266472
rect 121604 266432 121610 266444
rect 152458 266432 152464 266444
rect 152516 266432 152522 266484
rect 121454 266364 121460 266416
rect 121512 266404 121518 266416
rect 163498 266404 163504 266416
rect 121512 266376 163504 266404
rect 121512 266364 121518 266376
rect 163498 266364 163504 266376
rect 163556 266364 163562 266416
rect 45462 266296 45468 266348
rect 45520 266336 45526 266348
rect 67726 266336 67732 266348
rect 45520 266308 67732 266336
rect 45520 266296 45526 266308
rect 67726 266296 67732 266308
rect 67784 266296 67790 266348
rect 123662 266296 123668 266348
rect 123720 266336 123726 266348
rect 176654 266336 176660 266348
rect 123720 266308 176660 266336
rect 123720 266296 123726 266308
rect 176654 266296 176660 266308
rect 176712 266296 176718 266348
rect 121546 265004 121552 265056
rect 121604 265044 121610 265056
rect 127802 265044 127808 265056
rect 121604 265016 127808 265044
rect 121604 265004 121610 265016
rect 127802 265004 127808 265016
rect 127860 265004 127866 265056
rect 53558 264936 53564 264988
rect 53616 264976 53622 264988
rect 67634 264976 67640 264988
rect 53616 264948 67640 264976
rect 53616 264936 53622 264948
rect 67634 264936 67640 264948
rect 67692 264936 67698 264988
rect 121454 264936 121460 264988
rect 121512 264976 121518 264988
rect 178678 264976 178684 264988
rect 121512 264948 178684 264976
rect 121512 264936 121518 264948
rect 178678 264936 178684 264948
rect 178736 264936 178742 264988
rect 295610 264936 295616 264988
rect 295668 264976 295674 264988
rect 331858 264976 331864 264988
rect 295668 264948 331864 264976
rect 295668 264936 295674 264948
rect 331858 264936 331864 264948
rect 331916 264936 331922 264988
rect 48222 263644 48228 263696
rect 48280 263684 48286 263696
rect 67634 263684 67640 263696
rect 48280 263656 67640 263684
rect 48280 263644 48286 263656
rect 67634 263644 67640 263656
rect 67692 263644 67698 263696
rect 21358 263576 21364 263628
rect 21416 263616 21422 263628
rect 60458 263616 60464 263628
rect 21416 263588 60464 263616
rect 21416 263576 21422 263588
rect 60458 263576 60464 263588
rect 60516 263616 60522 263628
rect 67726 263616 67732 263628
rect 60516 263588 67732 263616
rect 60516 263576 60522 263588
rect 67726 263576 67732 263588
rect 67784 263576 67790 263628
rect 121546 263576 121552 263628
rect 121604 263616 121610 263628
rect 148594 263616 148600 263628
rect 121604 263588 148600 263616
rect 121604 263576 121610 263588
rect 148594 263576 148600 263588
rect 148652 263576 148658 263628
rect 295610 263576 295616 263628
rect 295668 263616 295674 263628
rect 305086 263616 305092 263628
rect 295668 263588 305092 263616
rect 295668 263576 295674 263588
rect 305086 263576 305092 263588
rect 305144 263576 305150 263628
rect 121454 263508 121460 263560
rect 121512 263548 121518 263560
rect 169018 263548 169024 263560
rect 121512 263520 169024 263548
rect 121512 263508 121518 263520
rect 169018 263508 169024 263520
rect 169076 263508 169082 263560
rect 17218 262828 17224 262880
rect 17276 262868 17282 262880
rect 53834 262868 53840 262880
rect 17276 262840 53840 262868
rect 17276 262828 17282 262840
rect 53834 262828 53840 262840
rect 53892 262828 53898 262880
rect 56410 262284 56416 262336
rect 56468 262324 56474 262336
rect 67634 262324 67640 262336
rect 56468 262296 67640 262324
rect 56468 262284 56474 262296
rect 67634 262284 67640 262296
rect 67692 262284 67698 262336
rect 53834 262216 53840 262268
rect 53892 262256 53898 262268
rect 54846 262256 54852 262268
rect 53892 262228 54852 262256
rect 53892 262216 53898 262228
rect 54846 262216 54852 262228
rect 54904 262256 54910 262268
rect 67726 262256 67732 262268
rect 54904 262228 67732 262256
rect 54904 262216 54910 262228
rect 67726 262216 67732 262228
rect 67784 262216 67790 262268
rect 121454 262216 121460 262268
rect 121512 262256 121518 262268
rect 129274 262256 129280 262268
rect 121512 262228 129280 262256
rect 121512 262216 121518 262228
rect 129274 262216 129280 262228
rect 129332 262216 129338 262268
rect 121546 262148 121552 262200
rect 121604 262188 121610 262200
rect 171778 262188 171784 262200
rect 121604 262160 171784 262188
rect 121604 262148 121610 262160
rect 171778 262148 171784 262160
rect 171836 262148 171842 262200
rect 160002 262080 160008 262132
rect 160060 262120 160066 262132
rect 176654 262120 176660 262132
rect 160060 262092 176660 262120
rect 160060 262080 160066 262092
rect 176654 262080 176660 262092
rect 176712 262080 176718 262132
rect 3050 261468 3056 261520
rect 3108 261508 3114 261520
rect 62758 261508 62764 261520
rect 3108 261480 62764 261508
rect 3108 261468 3114 261480
rect 62758 261468 62764 261480
rect 62816 261468 62822 261520
rect 121638 260856 121644 260908
rect 121696 260896 121702 260908
rect 170582 260896 170588 260908
rect 121696 260868 170588 260896
rect 121696 260856 121702 260868
rect 170582 260856 170588 260868
rect 170640 260856 170646 260908
rect 295610 260856 295616 260908
rect 295668 260896 295674 260908
rect 309778 260896 309784 260908
rect 295668 260868 309784 260896
rect 295668 260856 295674 260868
rect 309778 260856 309784 260868
rect 309836 260856 309842 260908
rect 13078 260788 13084 260840
rect 13136 260828 13142 260840
rect 55030 260828 55036 260840
rect 13136 260800 55036 260828
rect 13136 260788 13142 260800
rect 55030 260788 55036 260800
rect 55088 260828 55094 260840
rect 67634 260828 67640 260840
rect 55088 260800 67640 260828
rect 55088 260788 55094 260800
rect 67634 260788 67640 260800
rect 67692 260788 67698 260840
rect 121454 260788 121460 260840
rect 121512 260828 121518 260840
rect 170398 260828 170404 260840
rect 121512 260800 170404 260828
rect 121512 260788 121518 260800
rect 170398 260788 170404 260800
rect 170456 260788 170462 260840
rect 160002 259496 160008 259548
rect 160060 259536 160066 259548
rect 176654 259536 176660 259548
rect 160060 259508 176660 259536
rect 160060 259496 160066 259508
rect 176654 259496 176660 259508
rect 176712 259496 176718 259548
rect 121454 259428 121460 259480
rect 121512 259468 121518 259480
rect 169018 259468 169024 259480
rect 121512 259440 169024 259468
rect 121512 259428 121518 259440
rect 169018 259428 169024 259440
rect 169076 259428 169082 259480
rect 311158 259360 311164 259412
rect 311216 259400 311222 259412
rect 579614 259400 579620 259412
rect 311216 259372 579620 259400
rect 311216 259360 311222 259372
rect 579614 259360 579620 259372
rect 579672 259360 579678 259412
rect 57698 258136 57704 258188
rect 57756 258176 57762 258188
rect 67726 258176 67732 258188
rect 57756 258148 67732 258176
rect 57756 258136 57762 258148
rect 67726 258136 67732 258148
rect 67784 258136 67790 258188
rect 55030 258068 55036 258120
rect 55088 258108 55094 258120
rect 67634 258108 67640 258120
rect 55088 258080 67640 258108
rect 55088 258068 55094 258080
rect 67634 258068 67640 258080
rect 67692 258068 67698 258120
rect 121454 258068 121460 258120
rect 121512 258108 121518 258120
rect 171870 258108 171876 258120
rect 121512 258080 171876 258108
rect 121512 258068 121518 258080
rect 171870 258068 171876 258080
rect 171928 258068 171934 258120
rect 305638 257320 305644 257372
rect 305696 257360 305702 257372
rect 340874 257360 340880 257372
rect 305696 257332 340880 257360
rect 305696 257320 305702 257332
rect 340874 257320 340880 257332
rect 340932 257320 340938 257372
rect 295702 257048 295708 257100
rect 295760 257088 295766 257100
rect 298186 257088 298192 257100
rect 295760 257060 298192 257088
rect 295760 257048 295766 257060
rect 298186 257048 298192 257060
rect 298244 257048 298250 257100
rect 60366 256776 60372 256828
rect 60424 256816 60430 256828
rect 67634 256816 67640 256828
rect 60424 256788 67640 256816
rect 60424 256776 60430 256788
rect 67634 256776 67640 256788
rect 67692 256776 67698 256828
rect 121546 256776 121552 256828
rect 121604 256816 121610 256828
rect 140314 256816 140320 256828
rect 121604 256788 140320 256816
rect 121604 256776 121610 256788
rect 140314 256776 140320 256788
rect 140372 256776 140378 256828
rect 13078 256708 13084 256760
rect 13136 256748 13142 256760
rect 69014 256748 69020 256760
rect 13136 256720 69020 256748
rect 13136 256708 13142 256720
rect 69014 256708 69020 256720
rect 69072 256708 69078 256760
rect 121454 256708 121460 256760
rect 121512 256748 121518 256760
rect 159450 256748 159456 256760
rect 121512 256720 159456 256748
rect 121512 256708 121518 256720
rect 159450 256708 159456 256720
rect 159508 256708 159514 256760
rect 122098 255960 122104 256012
rect 122156 256000 122162 256012
rect 169202 256000 169208 256012
rect 122156 255972 169208 256000
rect 122156 255960 122162 255972
rect 169202 255960 169208 255972
rect 169260 255960 169266 256012
rect 63310 255280 63316 255332
rect 63368 255320 63374 255332
rect 67634 255320 67640 255332
rect 63368 255292 67640 255320
rect 63368 255280 63374 255292
rect 67634 255280 67640 255292
rect 67692 255280 67698 255332
rect 122466 254532 122472 254584
rect 122524 254572 122530 254584
rect 169110 254572 169116 254584
rect 122524 254544 169116 254572
rect 122524 254532 122530 254544
rect 169110 254532 169116 254544
rect 169168 254532 169174 254584
rect 2774 254056 2780 254108
rect 2832 254096 2838 254108
rect 4798 254096 4804 254108
rect 2832 254068 4804 254096
rect 2832 254056 2838 254068
rect 4798 254056 4804 254068
rect 4856 254056 4862 254108
rect 61930 253988 61936 254040
rect 61988 254028 61994 254040
rect 67634 254028 67640 254040
rect 61988 254000 67640 254028
rect 61988 253988 61994 254000
rect 67634 253988 67640 254000
rect 67692 253988 67698 254040
rect 61838 253920 61844 253972
rect 61896 253960 61902 253972
rect 67726 253960 67732 253972
rect 61896 253932 67732 253960
rect 61896 253920 61902 253932
rect 67726 253920 67732 253932
rect 67784 253920 67790 253972
rect 121454 253920 121460 253972
rect 121512 253960 121518 253972
rect 170398 253960 170404 253972
rect 121512 253932 170404 253960
rect 121512 253920 121518 253932
rect 170398 253920 170404 253932
rect 170456 253920 170462 253972
rect 295702 253920 295708 253972
rect 295760 253960 295766 253972
rect 335354 253960 335360 253972
rect 295760 253932 335360 253960
rect 295760 253920 295766 253932
rect 335354 253920 335360 253932
rect 335412 253920 335418 253972
rect 50522 253852 50528 253904
rect 50580 253892 50586 253904
rect 50890 253892 50896 253904
rect 50580 253864 50896 253892
rect 50580 253852 50586 253864
rect 50890 253852 50896 253864
rect 50948 253892 50954 253904
rect 67634 253892 67640 253904
rect 50948 253864 67640 253892
rect 50948 253852 50954 253864
rect 67634 253852 67640 253864
rect 67692 253852 67698 253904
rect 295518 253444 295524 253496
rect 295576 253484 295582 253496
rect 295702 253484 295708 253496
rect 295576 253456 295708 253484
rect 295576 253444 295582 253456
rect 295702 253444 295708 253456
rect 295760 253444 295766 253496
rect 25498 253172 25504 253224
rect 25556 253212 25562 253224
rect 50522 253212 50528 253224
rect 25556 253184 50528 253212
rect 25556 253172 25562 253184
rect 50522 253172 50528 253184
rect 50580 253172 50586 253224
rect 121546 252628 121552 252680
rect 121604 252668 121610 252680
rect 155310 252668 155316 252680
rect 121604 252640 155316 252668
rect 121604 252628 121610 252640
rect 155310 252628 155316 252640
rect 155368 252628 155374 252680
rect 50890 252560 50896 252612
rect 50948 252600 50954 252612
rect 67634 252600 67640 252612
rect 50948 252572 67640 252600
rect 50948 252560 50954 252572
rect 67634 252560 67640 252572
rect 67692 252560 67698 252612
rect 121454 252560 121460 252612
rect 121512 252600 121518 252612
rect 173250 252600 173256 252612
rect 121512 252572 173256 252600
rect 121512 252560 121518 252572
rect 173250 252560 173256 252572
rect 173308 252560 173314 252612
rect 64506 251880 64512 251932
rect 64564 251920 64570 251932
rect 68094 251920 68100 251932
rect 64564 251892 68100 251920
rect 64564 251880 64570 251892
rect 68094 251880 68100 251892
rect 68152 251880 68158 251932
rect 59262 251812 59268 251864
rect 59320 251852 59326 251864
rect 68370 251852 68376 251864
rect 59320 251824 68376 251852
rect 59320 251812 59326 251824
rect 68370 251812 68376 251824
rect 68428 251812 68434 251864
rect 302418 251812 302424 251864
rect 302476 251852 302482 251864
rect 319438 251852 319444 251864
rect 302476 251824 319444 251852
rect 302476 251812 302482 251824
rect 319438 251812 319444 251824
rect 319496 251812 319502 251864
rect 56318 251268 56324 251320
rect 56376 251308 56382 251320
rect 67634 251308 67640 251320
rect 56376 251280 67640 251308
rect 56376 251268 56382 251280
rect 67634 251268 67640 251280
rect 67692 251268 67698 251320
rect 121454 251200 121460 251252
rect 121512 251240 121518 251252
rect 166442 251240 166448 251252
rect 121512 251212 166448 251240
rect 121512 251200 121518 251212
rect 166442 251200 166448 251212
rect 166500 251200 166506 251252
rect 296438 251200 296444 251252
rect 296496 251240 296502 251252
rect 302418 251240 302424 251252
rect 296496 251212 302424 251240
rect 296496 251200 296502 251212
rect 302418 251200 302424 251212
rect 302476 251200 302482 251252
rect 120626 251132 120632 251184
rect 120684 251172 120690 251184
rect 127710 251172 127716 251184
rect 120684 251144 127716 251172
rect 120684 251132 120690 251144
rect 127710 251132 127716 251144
rect 127768 251132 127774 251184
rect 295334 250860 295340 250912
rect 295392 250900 295398 250912
rect 295518 250900 295524 250912
rect 295392 250872 295524 250900
rect 295392 250860 295398 250872
rect 295518 250860 295524 250872
rect 295576 250860 295582 250912
rect 60550 249772 60556 249824
rect 60608 249812 60614 249824
rect 67634 249812 67640 249824
rect 60608 249784 67640 249812
rect 60608 249772 60614 249784
rect 67634 249772 67640 249784
rect 67692 249772 67698 249824
rect 121454 249772 121460 249824
rect 121512 249812 121518 249824
rect 130654 249812 130660 249824
rect 121512 249784 130660 249812
rect 121512 249772 121518 249784
rect 130654 249772 130660 249784
rect 130712 249772 130718 249824
rect 172422 249772 172428 249824
rect 172480 249812 172486 249824
rect 176654 249812 176660 249824
rect 172480 249784 176660 249812
rect 172480 249772 172486 249784
rect 176654 249772 176660 249784
rect 176712 249772 176718 249824
rect 295794 249772 295800 249824
rect 295852 249812 295858 249824
rect 319438 249812 319444 249824
rect 295852 249784 319444 249812
rect 295852 249772 295858 249784
rect 319438 249772 319444 249784
rect 319496 249772 319502 249824
rect 68922 249704 68928 249756
rect 68980 249744 68986 249756
rect 69658 249744 69664 249756
rect 68980 249716 69664 249744
rect 68980 249704 68986 249716
rect 69658 249704 69664 249716
rect 69716 249704 69722 249756
rect 65978 248616 65984 248668
rect 66036 248656 66042 248668
rect 67818 248656 67824 248668
rect 66036 248628 67824 248656
rect 66036 248616 66042 248628
rect 67818 248616 67824 248628
rect 67876 248616 67882 248668
rect 121546 248480 121552 248532
rect 121604 248520 121610 248532
rect 161014 248520 161020 248532
rect 121604 248492 161020 248520
rect 121604 248480 121610 248492
rect 161014 248480 161020 248492
rect 161072 248480 161078 248532
rect 121454 248412 121460 248464
rect 121512 248452 121518 248464
rect 173342 248452 173348 248464
rect 121512 248424 173348 248452
rect 121512 248412 121518 248424
rect 173342 248412 173348 248424
rect 173400 248412 173406 248464
rect 121546 248344 121552 248396
rect 121604 248384 121610 248396
rect 140130 248384 140136 248396
rect 121604 248356 140136 248384
rect 121604 248344 121610 248356
rect 140130 248344 140136 248356
rect 140188 248344 140194 248396
rect 296622 248344 296628 248396
rect 296680 248384 296686 248396
rect 299658 248384 299664 248396
rect 296680 248356 299664 248384
rect 296680 248344 296686 248356
rect 299658 248344 299664 248356
rect 299716 248384 299722 248396
rect 324958 248384 324964 248396
rect 299716 248356 324964 248384
rect 299716 248344 299722 248356
rect 324958 248344 324964 248356
rect 325016 248344 325022 248396
rect 59170 247120 59176 247172
rect 59228 247160 59234 247172
rect 67634 247160 67640 247172
rect 59228 247132 67640 247160
rect 59228 247120 59234 247132
rect 67634 247120 67640 247132
rect 67692 247120 67698 247172
rect 57790 247052 57796 247104
rect 57848 247092 57854 247104
rect 67726 247092 67732 247104
rect 57848 247064 67732 247092
rect 57848 247052 57854 247064
rect 67726 247052 67732 247064
rect 67784 247052 67790 247104
rect 121454 247052 121460 247104
rect 121512 247092 121518 247104
rect 144546 247092 144552 247104
rect 121512 247064 144552 247092
rect 121512 247052 121518 247064
rect 144546 247052 144552 247064
rect 144604 247052 144610 247104
rect 143074 246304 143080 246356
rect 143132 246344 143138 246356
rect 174630 246344 174636 246356
rect 143132 246316 174636 246344
rect 143132 246304 143138 246316
rect 174630 246304 174636 246316
rect 174688 246304 174694 246356
rect 121454 245692 121460 245744
rect 121512 245732 121518 245744
rect 142982 245732 142988 245744
rect 121512 245704 142988 245732
rect 121512 245692 121518 245704
rect 142982 245692 142988 245704
rect 143040 245692 143046 245744
rect 121546 245624 121552 245676
rect 121604 245664 121610 245676
rect 149790 245664 149796 245676
rect 121604 245636 149796 245664
rect 121604 245624 121610 245636
rect 149790 245624 149796 245636
rect 149848 245624 149854 245676
rect 296898 245624 296904 245676
rect 296956 245664 296962 245676
rect 467098 245664 467104 245676
rect 296956 245636 467104 245664
rect 296956 245624 296962 245636
rect 467098 245624 467104 245636
rect 467156 245624 467162 245676
rect 121454 245556 121460 245608
rect 121512 245596 121518 245608
rect 162118 245596 162124 245608
rect 121512 245568 162124 245596
rect 121512 245556 121518 245568
rect 162118 245556 162124 245568
rect 162176 245556 162182 245608
rect 147030 245012 147036 245064
rect 147088 245052 147094 245064
rect 171778 245052 171784 245064
rect 147088 245024 171784 245052
rect 147088 245012 147094 245024
rect 171778 245012 171784 245024
rect 171836 245012 171842 245064
rect 120718 244944 120724 244996
rect 120776 244984 120782 244996
rect 158070 244984 158076 244996
rect 120776 244956 158076 244984
rect 120776 244944 120782 244956
rect 158070 244944 158076 244956
rect 158128 244944 158134 244996
rect 53098 244876 53104 244928
rect 53156 244916 53162 244928
rect 59078 244916 59084 244928
rect 53156 244888 59084 244916
rect 53156 244876 53162 244888
rect 59078 244876 59084 244888
rect 59136 244876 59142 244928
rect 119798 244876 119804 244928
rect 119856 244916 119862 244928
rect 162302 244916 162308 244928
rect 119856 244888 162308 244916
rect 119856 244876 119862 244888
rect 162302 244876 162308 244888
rect 162360 244876 162366 244928
rect 59078 244264 59084 244316
rect 59136 244304 59142 244316
rect 67634 244304 67640 244316
rect 59136 244276 67640 244304
rect 59136 244264 59142 244276
rect 67634 244264 67640 244276
rect 67692 244264 67698 244316
rect 121546 244264 121552 244316
rect 121604 244304 121610 244316
rect 170674 244304 170680 244316
rect 121604 244276 170680 244304
rect 121604 244264 121610 244276
rect 170674 244264 170680 244276
rect 170732 244264 170738 244316
rect 574738 244264 574744 244316
rect 574796 244304 574802 244316
rect 579890 244304 579896 244316
rect 574796 244276 579896 244304
rect 574796 244264 574802 244276
rect 579890 244264 579896 244276
rect 579948 244264 579954 244316
rect 8938 244196 8944 244248
rect 8996 244236 9002 244248
rect 69198 244236 69204 244248
rect 8996 244208 69204 244236
rect 8996 244196 9002 244208
rect 69198 244196 69204 244208
rect 69256 244196 69262 244248
rect 121546 242972 121552 243024
rect 121604 243012 121610 243024
rect 147030 243012 147036 243024
rect 121604 242984 147036 243012
rect 121604 242972 121610 242984
rect 147030 242972 147036 242984
rect 147088 242972 147094 243024
rect 121454 242904 121460 242956
rect 121512 242944 121518 242956
rect 179690 242944 179696 242956
rect 121512 242916 179696 242944
rect 121512 242904 121518 242916
rect 179690 242904 179696 242916
rect 179748 242904 179754 242956
rect 295334 242904 295340 242956
rect 295392 242944 295398 242956
rect 299658 242944 299664 242956
rect 295392 242916 299664 242944
rect 295392 242904 295398 242916
rect 299658 242904 299664 242916
rect 299716 242944 299722 242956
rect 395338 242944 395344 242956
rect 299716 242916 395344 242944
rect 299716 242904 299722 242916
rect 395338 242904 395344 242916
rect 395396 242904 395402 242956
rect 121546 242836 121552 242888
rect 121604 242876 121610 242888
rect 160738 242876 160744 242888
rect 121604 242848 160744 242876
rect 121604 242836 121610 242848
rect 160738 242836 160744 242848
rect 160796 242836 160802 242888
rect 121454 242768 121460 242820
rect 121512 242808 121518 242820
rect 158622 242808 158628 242820
rect 121512 242780 158628 242808
rect 121512 242768 121518 242780
rect 158622 242768 158628 242780
rect 158680 242808 158686 242820
rect 160922 242808 160928 242820
rect 158680 242780 160928 242808
rect 158680 242768 158686 242780
rect 160922 242768 160928 242780
rect 160980 242768 160986 242820
rect 147122 242700 147128 242752
rect 147180 242740 147186 242752
rect 176838 242740 176844 242752
rect 147180 242712 176844 242740
rect 147180 242700 147186 242712
rect 176838 242700 176844 242712
rect 176896 242700 176902 242752
rect 143166 242224 143172 242276
rect 143224 242264 143230 242276
rect 152734 242264 152740 242276
rect 143224 242236 152740 242264
rect 143224 242224 143230 242236
rect 152734 242224 152740 242236
rect 152792 242224 152798 242276
rect 125042 242156 125048 242208
rect 125100 242196 125106 242208
rect 154114 242196 154120 242208
rect 125100 242168 154120 242196
rect 125100 242156 125106 242168
rect 154114 242156 154120 242168
rect 154172 242156 154178 242208
rect 61746 241476 61752 241528
rect 61804 241516 61810 241528
rect 67726 241516 67732 241528
rect 61804 241488 67732 241516
rect 61804 241476 61810 241488
rect 67726 241476 67732 241488
rect 67784 241476 67790 241528
rect 57882 241408 57888 241460
rect 57940 241448 57946 241460
rect 67634 241448 67640 241460
rect 57940 241420 67640 241448
rect 57940 241408 57946 241420
rect 67634 241408 67640 241420
rect 67692 241408 67698 241460
rect 163682 241408 163688 241460
rect 163740 241448 163746 241460
rect 295518 241448 295524 241460
rect 163740 241420 295524 241448
rect 163740 241408 163746 241420
rect 295518 241408 295524 241420
rect 295576 241408 295582 241460
rect 127802 240796 127808 240848
rect 127860 240836 127866 240848
rect 156782 240836 156788 240848
rect 127860 240808 156788 240836
rect 127860 240796 127866 240808
rect 156782 240796 156788 240808
rect 156840 240796 156846 240848
rect 140222 240728 140228 240780
rect 140280 240768 140286 240780
rect 140280 240740 161474 240768
rect 140280 240728 140286 240740
rect 161446 240632 161474 240740
rect 182818 240632 182824 240644
rect 161446 240604 182824 240632
rect 182818 240592 182824 240604
rect 182876 240592 182882 240644
rect 179690 240320 179696 240372
rect 179748 240360 179754 240372
rect 179748 240332 179920 240360
rect 179748 240320 179754 240332
rect 69842 240184 69848 240236
rect 69900 240184 69906 240236
rect 69860 239952 69888 240184
rect 179892 240168 179920 240332
rect 121454 240116 121460 240168
rect 121512 240156 121518 240168
rect 144454 240156 144460 240168
rect 121512 240128 144460 240156
rect 121512 240116 121518 240128
rect 144454 240116 144460 240128
rect 144512 240116 144518 240168
rect 179874 240116 179880 240168
rect 179932 240116 179938 240168
rect 152642 240048 152648 240100
rect 152700 240088 152706 240100
rect 295702 240088 295708 240100
rect 152700 240060 295708 240088
rect 152700 240048 152706 240060
rect 295702 240048 295708 240060
rect 295760 240048 295766 240100
rect 75270 239952 75276 239964
rect 69860 239924 75276 239952
rect 75270 239912 75276 239924
rect 75328 239912 75334 239964
rect 118970 239912 118976 239964
rect 119028 239952 119034 239964
rect 119798 239952 119804 239964
rect 119028 239924 119804 239952
rect 119028 239912 119034 239924
rect 119798 239912 119804 239924
rect 119856 239912 119862 239964
rect 64506 239436 64512 239488
rect 64564 239476 64570 239488
rect 116578 239476 116584 239488
rect 64564 239448 116584 239476
rect 64564 239436 64570 239448
rect 116578 239436 116584 239448
rect 116636 239436 116642 239488
rect 3326 239368 3332 239420
rect 3384 239408 3390 239420
rect 70302 239408 70308 239420
rect 3384 239380 70308 239408
rect 3384 239368 3390 239380
rect 70302 239368 70308 239380
rect 70360 239368 70366 239420
rect 118602 239368 118608 239420
rect 118660 239408 118666 239420
rect 135254 239408 135260 239420
rect 118660 239380 135260 239408
rect 118660 239368 118666 239380
rect 135254 239368 135260 239380
rect 135312 239368 135318 239420
rect 287698 239368 287704 239420
rect 287756 239408 287762 239420
rect 296806 239408 296812 239420
rect 287756 239380 296812 239408
rect 287756 239368 287762 239380
rect 296806 239368 296812 239380
rect 296864 239368 296870 239420
rect 121546 238960 121552 239012
rect 121604 239000 121610 239012
rect 323578 239000 323584 239012
rect 121604 238972 323584 239000
rect 121604 238960 121610 238972
rect 323578 238960 323584 238972
rect 323636 238960 323642 239012
rect 60458 238892 60464 238944
rect 60516 238932 60522 238944
rect 252554 238932 252560 238944
rect 60516 238904 252560 238932
rect 60516 238892 60522 238904
rect 252554 238892 252560 238904
rect 252612 238892 252618 238944
rect 61930 238824 61936 238876
rect 61988 238864 61994 238876
rect 262214 238864 262220 238876
rect 61988 238836 262220 238864
rect 61988 238824 61994 238836
rect 262214 238824 262220 238836
rect 262272 238864 262278 238876
rect 262766 238864 262772 238876
rect 262272 238836 262772 238864
rect 262272 238824 262278 238836
rect 262766 238824 262772 238836
rect 262824 238824 262830 238876
rect 278866 238824 278872 238876
rect 278924 238864 278930 238876
rect 279970 238864 279976 238876
rect 278924 238836 279976 238864
rect 278924 238824 278930 238836
rect 279970 238824 279976 238836
rect 280028 238864 280034 238876
rect 310514 238864 310520 238876
rect 280028 238836 310520 238864
rect 280028 238824 280034 238836
rect 310514 238824 310520 238836
rect 310572 238824 310578 238876
rect 58618 238756 58624 238808
rect 58676 238796 58682 238808
rect 81526 238796 81532 238808
rect 58676 238768 81532 238796
rect 58676 238756 58682 238768
rect 81526 238756 81532 238768
rect 81584 238796 81590 238808
rect 82262 238796 82268 238808
rect 81584 238768 82268 238796
rect 81584 238756 81590 238768
rect 82262 238756 82268 238768
rect 82320 238756 82326 238808
rect 109034 238756 109040 238808
rect 109092 238796 109098 238808
rect 109954 238796 109960 238808
rect 109092 238768 109960 238796
rect 109092 238756 109098 238768
rect 109954 238756 109960 238768
rect 110012 238796 110018 238808
rect 120810 238796 120816 238808
rect 110012 238768 120816 238796
rect 110012 238756 110018 238768
rect 120810 238756 120816 238768
rect 120868 238756 120874 238808
rect 174538 238756 174544 238808
rect 174596 238796 174602 238808
rect 215294 238796 215300 238808
rect 174596 238768 215300 238796
rect 174596 238756 174602 238768
rect 215294 238756 215300 238768
rect 215352 238796 215358 238808
rect 525058 238796 525064 238808
rect 215352 238768 525064 238796
rect 215352 238756 215358 238768
rect 525058 238756 525064 238768
rect 525116 238756 525122 238808
rect 62758 238688 62764 238740
rect 62816 238728 62822 238740
rect 86770 238728 86776 238740
rect 62816 238700 86776 238728
rect 62816 238688 62822 238700
rect 86770 238688 86776 238700
rect 86828 238688 86834 238740
rect 114462 238688 114468 238740
rect 114520 238728 114526 238740
rect 118602 238728 118608 238740
rect 114520 238700 118608 238728
rect 114520 238688 114526 238700
rect 118602 238688 118608 238700
rect 118660 238688 118666 238740
rect 189994 238688 190000 238740
rect 190052 238728 190058 238740
rect 582558 238728 582564 238740
rect 190052 238700 582564 238728
rect 190052 238688 190058 238700
rect 582558 238688 582564 238700
rect 582616 238688 582622 238740
rect 70302 238620 70308 238672
rect 70360 238660 70366 238672
rect 103514 238660 103520 238672
rect 70360 238632 103520 238660
rect 70360 238620 70366 238632
rect 103514 238620 103520 238632
rect 103572 238660 103578 238672
rect 104710 238660 104716 238672
rect 103572 238632 104716 238660
rect 103572 238620 103578 238632
rect 104710 238620 104716 238632
rect 104768 238620 104774 238672
rect 107378 238620 107384 238672
rect 107436 238660 107442 238672
rect 130562 238660 130568 238672
rect 107436 238632 130568 238660
rect 107436 238620 107442 238632
rect 130562 238620 130568 238632
rect 130620 238620 130626 238672
rect 176010 238620 176016 238672
rect 176068 238660 176074 238672
rect 223850 238660 223856 238672
rect 176068 238632 223856 238660
rect 176068 238620 176074 238632
rect 223850 238620 223856 238632
rect 223908 238620 223914 238672
rect 235994 238620 236000 238672
rect 236052 238660 236058 238672
rect 582466 238660 582472 238672
rect 236052 238632 582472 238660
rect 236052 238620 236058 238632
rect 582466 238620 582472 238632
rect 582524 238620 582530 238672
rect 117682 238552 117688 238604
rect 117740 238592 117746 238604
rect 250806 238592 250812 238604
rect 117740 238564 250812 238592
rect 117740 238552 117746 238564
rect 250806 238552 250812 238564
rect 250864 238552 250870 238604
rect 99006 238484 99012 238536
rect 99064 238524 99070 238536
rect 120902 238524 120908 238536
rect 99064 238496 120908 238524
rect 99064 238484 99070 238496
rect 120902 238484 120908 238496
rect 120960 238484 120966 238536
rect 170490 238484 170496 238536
rect 170548 238524 170554 238536
rect 195974 238524 195980 238536
rect 170548 238496 195980 238524
rect 170548 238484 170554 238496
rect 195974 238484 195980 238496
rect 196032 238484 196038 238536
rect 110598 238416 110604 238468
rect 110656 238456 110662 238468
rect 126238 238456 126244 238468
rect 110656 238428 126244 238456
rect 110656 238416 110662 238428
rect 126238 238416 126244 238428
rect 126296 238416 126302 238468
rect 89346 238348 89352 238400
rect 89404 238388 89410 238400
rect 148318 238388 148324 238400
rect 89404 238360 148324 238388
rect 89404 238348 89410 238360
rect 148318 238348 148324 238360
rect 148376 238348 148382 238400
rect 86126 238212 86132 238264
rect 86184 238252 86190 238264
rect 95694 238252 95700 238264
rect 86184 238224 95700 238252
rect 86184 238212 86190 238224
rect 95694 238212 95700 238224
rect 95752 238212 95758 238264
rect 75822 238144 75828 238196
rect 75880 238184 75886 238196
rect 86218 238184 86224 238196
rect 75880 238156 86224 238184
rect 75880 238144 75886 238156
rect 86218 238144 86224 238156
rect 86276 238144 86282 238196
rect 70670 238076 70676 238128
rect 70728 238116 70734 238128
rect 147122 238116 147128 238128
rect 70728 238088 147128 238116
rect 70728 238076 70734 238088
rect 147122 238076 147128 238088
rect 147180 238076 147186 238128
rect 4798 238008 4804 238060
rect 4856 238048 4862 238060
rect 112530 238048 112536 238060
rect 4856 238020 112536 238048
rect 4856 238008 4862 238020
rect 112530 238008 112536 238020
rect 112588 238008 112594 238060
rect 155402 238008 155408 238060
rect 155460 238048 155466 238060
rect 189718 238048 189724 238060
rect 155460 238020 189724 238048
rect 155460 238008 155466 238020
rect 189718 238008 189724 238020
rect 189776 238008 189782 238060
rect 110598 237804 110604 237856
rect 110656 237844 110662 237856
rect 111058 237844 111064 237856
rect 110656 237816 111064 237844
rect 110656 237804 110662 237816
rect 111058 237804 111064 237816
rect 111116 237804 111122 237856
rect 104158 237396 104164 237448
rect 104216 237436 104222 237448
rect 106918 237436 106924 237448
rect 104216 237408 106924 237436
rect 104216 237396 104222 237408
rect 106918 237396 106924 237408
rect 106976 237396 106982 237448
rect 215938 237396 215944 237448
rect 215996 237436 216002 237448
rect 217042 237436 217048 237448
rect 215996 237408 217048 237436
rect 215996 237396 216002 237408
rect 217042 237396 217048 237408
rect 217100 237396 217106 237448
rect 224126 237396 224132 237448
rect 224184 237436 224190 237448
rect 240042 237436 240048 237448
rect 224184 237408 240048 237436
rect 224184 237396 224190 237408
rect 240042 237396 240048 237408
rect 240100 237396 240106 237448
rect 291838 237396 291844 237448
rect 291896 237436 291902 237448
rect 292574 237436 292580 237448
rect 291896 237408 292580 237436
rect 291896 237396 291902 237408
rect 292574 237396 292580 237408
rect 292632 237396 292638 237448
rect 91922 237328 91928 237380
rect 91980 237368 91986 237380
rect 134518 237368 134524 237380
rect 91980 237340 134524 237368
rect 91980 237328 91986 237340
rect 134518 237328 134524 237340
rect 134576 237328 134582 237380
rect 166350 237328 166356 237380
rect 166408 237368 166414 237380
rect 580350 237368 580356 237380
rect 166408 237340 580356 237368
rect 166408 237328 166414 237340
rect 580350 237328 580356 237340
rect 580408 237328 580414 237380
rect 112530 237260 112536 237312
rect 112588 237300 112594 237312
rect 144178 237300 144184 237312
rect 112588 237272 144184 237300
rect 112588 237260 112594 237272
rect 144178 237260 144184 237272
rect 144236 237260 144242 237312
rect 161014 237260 161020 237312
rect 161072 237300 161078 237312
rect 314654 237300 314660 237312
rect 161072 237272 314660 237300
rect 161072 237260 161078 237272
rect 314654 237260 314660 237272
rect 314712 237260 314718 237312
rect 63218 237192 63224 237244
rect 63276 237232 63282 237244
rect 191926 237232 191932 237244
rect 63276 237204 191932 237232
rect 63276 237192 63282 237204
rect 191926 237192 191932 237204
rect 191984 237192 191990 237244
rect 233878 237192 233884 237244
rect 233936 237232 233942 237244
rect 364334 237232 364340 237244
rect 233936 237204 364340 237232
rect 233936 237192 233942 237204
rect 364334 237192 364340 237204
rect 364392 237192 364398 237244
rect 188338 237124 188344 237176
rect 188396 237164 188402 237176
rect 254394 237164 254400 237176
rect 188396 237136 254400 237164
rect 188396 237124 188402 237136
rect 254394 237124 254400 237136
rect 254452 237124 254458 237176
rect 173342 236716 173348 236768
rect 173400 236756 173406 236768
rect 192478 236756 192484 236768
rect 173400 236728 192484 236756
rect 173400 236716 173406 236728
rect 192478 236716 192484 236728
rect 192536 236716 192542 236768
rect 40034 236648 40040 236700
rect 40092 236688 40098 236700
rect 95050 236688 95056 236700
rect 40092 236660 95056 236688
rect 40092 236648 40098 236660
rect 95050 236648 95056 236660
rect 95108 236688 95114 236700
rect 95786 236688 95792 236700
rect 95108 236660 95792 236688
rect 95108 236648 95114 236660
rect 95786 236648 95792 236660
rect 95844 236648 95850 236700
rect 141510 236648 141516 236700
rect 141568 236688 141574 236700
rect 242250 236688 242256 236700
rect 141568 236660 242256 236688
rect 141568 236648 141574 236660
rect 242250 236648 242256 236660
rect 242308 236648 242314 236700
rect 113818 235900 113824 235952
rect 113876 235940 113882 235952
rect 300854 235940 300860 235952
rect 113876 235912 300860 235940
rect 113876 235900 113882 235912
rect 300854 235900 300860 235912
rect 300912 235900 300918 235952
rect 72602 235832 72608 235884
rect 72660 235872 72666 235884
rect 123570 235872 123576 235884
rect 72660 235844 123576 235872
rect 72660 235832 72666 235844
rect 123570 235832 123576 235844
rect 123628 235832 123634 235884
rect 159450 235832 159456 235884
rect 159508 235872 159514 235884
rect 310606 235872 310612 235884
rect 159508 235844 310612 235872
rect 159508 235832 159514 235844
rect 310606 235832 310612 235844
rect 310664 235832 310670 235884
rect 95050 235764 95056 235816
rect 95108 235804 95114 235816
rect 142798 235804 142804 235816
rect 95108 235776 142804 235804
rect 95108 235764 95114 235776
rect 142798 235764 142804 235776
rect 142856 235764 142862 235816
rect 169202 235764 169208 235816
rect 169260 235804 169266 235816
rect 295610 235804 295616 235816
rect 169260 235776 295616 235804
rect 169260 235764 169266 235776
rect 295610 235764 295616 235776
rect 295668 235764 295674 235816
rect 276290 235696 276296 235748
rect 276348 235736 276354 235748
rect 276658 235736 276664 235748
rect 276348 235708 276664 235736
rect 276348 235696 276354 235708
rect 276658 235696 276664 235708
rect 276716 235736 276722 235748
rect 304994 235736 305000 235748
rect 276716 235708 305000 235736
rect 276716 235696 276722 235708
rect 304994 235696 305000 235708
rect 305052 235696 305058 235748
rect 170582 235356 170588 235408
rect 170640 235396 170646 235408
rect 197998 235396 198004 235408
rect 170640 235368 198004 235396
rect 170640 235356 170646 235368
rect 197998 235356 198004 235368
rect 198056 235356 198062 235408
rect 60366 235288 60372 235340
rect 60424 235328 60430 235340
rect 159542 235328 159548 235340
rect 60424 235300 159548 235328
rect 60424 235288 60430 235300
rect 159542 235288 159548 235300
rect 159600 235288 159606 235340
rect 171870 235288 171876 235340
rect 171928 235328 171934 235340
rect 222838 235328 222844 235340
rect 171928 235300 222844 235328
rect 171928 235288 171934 235300
rect 222838 235288 222844 235300
rect 222896 235288 222902 235340
rect 152550 235220 152556 235272
rect 152608 235260 152614 235272
rect 260098 235260 260104 235272
rect 152608 235232 260104 235260
rect 152608 235220 152614 235232
rect 260098 235220 260104 235232
rect 260156 235220 260162 235272
rect 46750 234540 46756 234592
rect 46808 234580 46814 234592
rect 303706 234580 303712 234592
rect 46808 234552 303712 234580
rect 46808 234540 46814 234552
rect 303706 234540 303712 234552
rect 303764 234540 303770 234592
rect 91278 234472 91284 234524
rect 91336 234512 91342 234524
rect 129182 234512 129188 234524
rect 91336 234484 129188 234512
rect 91336 234472 91342 234484
rect 129182 234472 129188 234484
rect 129240 234472 129246 234524
rect 151262 234472 151268 234524
rect 151320 234512 151326 234524
rect 298186 234512 298192 234524
rect 151320 234484 298192 234512
rect 151320 234472 151326 234484
rect 298186 234472 298192 234484
rect 298244 234472 298250 234524
rect 264974 234404 264980 234456
rect 265032 234444 265038 234456
rect 265618 234444 265624 234456
rect 265032 234416 265624 234444
rect 265032 234404 265038 234416
rect 265618 234404 265624 234416
rect 265676 234444 265682 234456
rect 306466 234444 306472 234456
rect 265676 234416 306472 234444
rect 265676 234404 265682 234416
rect 306466 234404 306472 234416
rect 306524 234404 306530 234456
rect 46198 234132 46204 234184
rect 46256 234172 46262 234184
rect 46750 234172 46756 234184
rect 46256 234144 46756 234172
rect 46256 234132 46262 234144
rect 46750 234132 46756 234144
rect 46808 234132 46814 234184
rect 149882 233996 149888 234048
rect 149940 234036 149946 234048
rect 186958 234036 186964 234048
rect 149940 234008 186964 234036
rect 149940 233996 149946 234008
rect 186958 233996 186964 234008
rect 187016 233996 187022 234048
rect 69014 233928 69020 233980
rect 69072 233968 69078 233980
rect 69750 233968 69756 233980
rect 69072 233940 69756 233968
rect 69072 233928 69078 233940
rect 69750 233928 69756 233940
rect 69808 233928 69814 233980
rect 75914 233928 75920 233980
rect 75972 233968 75978 233980
rect 77110 233968 77116 233980
rect 75972 233940 77116 233968
rect 75972 233928 75978 233940
rect 77110 233928 77116 233940
rect 77168 233928 77174 233980
rect 77294 233928 77300 233980
rect 77352 233968 77358 233980
rect 78398 233968 78404 233980
rect 77352 233940 78404 233968
rect 77352 233928 77358 233940
rect 78398 233928 78404 233940
rect 78456 233928 78462 233980
rect 78674 233928 78680 233980
rect 78732 233968 78738 233980
rect 79686 233968 79692 233980
rect 78732 233940 79692 233968
rect 78732 233928 78738 233940
rect 79686 233928 79692 233940
rect 79744 233928 79750 233980
rect 84286 233928 84292 233980
rect 84344 233968 84350 233980
rect 85482 233968 85488 233980
rect 84344 233940 85488 233968
rect 84344 233928 84350 233940
rect 85482 233928 85488 233940
rect 85540 233928 85546 233980
rect 93854 233928 93860 233980
rect 93912 233968 93918 233980
rect 94498 233968 94504 233980
rect 93912 233940 94504 233968
rect 93912 233928 93918 233940
rect 94498 233928 94504 233940
rect 94556 233928 94562 233980
rect 96614 233928 96620 233980
rect 96672 233968 96678 233980
rect 97718 233968 97724 233980
rect 96672 233940 97724 233968
rect 96672 233928 96678 233940
rect 97718 233928 97724 233940
rect 97776 233928 97782 233980
rect 100754 233928 100760 233980
rect 100812 233968 100818 233980
rect 101582 233968 101588 233980
rect 100812 233940 101588 233968
rect 100812 233928 100818 233940
rect 101582 233928 101588 233940
rect 101640 233928 101646 233980
rect 102134 233928 102140 233980
rect 102192 233968 102198 233980
rect 102870 233968 102876 233980
rect 102192 233940 102876 233968
rect 102192 233928 102198 233940
rect 102870 233928 102876 233940
rect 102928 233928 102934 233980
rect 104894 233928 104900 233980
rect 104952 233968 104958 233980
rect 106090 233968 106096 233980
rect 104952 233940 106096 233968
rect 104952 233928 104958 233940
rect 106090 233928 106096 233940
rect 106148 233928 106154 233980
rect 114554 233928 114560 233980
rect 114612 233968 114618 233980
rect 115750 233968 115756 233980
rect 114612 233940 115756 233968
rect 114612 233928 114618 233940
rect 115750 233928 115756 233940
rect 115808 233928 115814 233980
rect 174630 233928 174636 233980
rect 174688 233968 174694 233980
rect 255958 233968 255964 233980
rect 174688 233940 255964 233968
rect 174688 233928 174694 233940
rect 255958 233928 255964 233940
rect 256016 233928 256022 233980
rect 62022 233860 62028 233912
rect 62080 233900 62086 233912
rect 196710 233900 196716 233912
rect 62080 233872 196716 233900
rect 62080 233860 62086 233872
rect 196710 233860 196716 233872
rect 196768 233860 196774 233912
rect 289814 233656 289820 233708
rect 289872 233696 289878 233708
rect 294138 233696 294144 233708
rect 289872 233668 294144 233696
rect 289872 233656 289878 233668
rect 294138 233656 294144 233668
rect 294196 233656 294202 233708
rect 92474 233384 92480 233436
rect 92532 233424 92538 233436
rect 93210 233424 93216 233436
rect 92532 233396 93216 233424
rect 92532 233384 92538 233396
rect 93210 233384 93216 233396
rect 93268 233384 93274 233436
rect 59078 233180 59084 233232
rect 59136 233220 59142 233232
rect 218974 233220 218980 233232
rect 59136 233192 218980 233220
rect 59136 233180 59142 233192
rect 218974 233180 218980 233192
rect 219032 233180 219038 233232
rect 223850 233180 223856 233232
rect 223908 233220 223914 233232
rect 582650 233220 582656 233232
rect 223908 233192 582656 233220
rect 223908 233180 223914 233192
rect 582650 233180 582656 233192
rect 582708 233180 582714 233232
rect 86770 233112 86776 233164
rect 86828 233152 86834 233164
rect 210602 233152 210608 233164
rect 86828 233124 210608 233152
rect 86828 233112 86834 233124
rect 210602 233112 210608 233124
rect 210660 233112 210666 233164
rect 240042 233112 240048 233164
rect 240100 233152 240106 233164
rect 582374 233152 582380 233164
rect 240100 233124 582380 233152
rect 240100 233112 240106 233124
rect 582374 233112 582380 233124
rect 582432 233112 582438 233164
rect 115106 233044 115112 233096
rect 115164 233084 115170 233096
rect 235994 233084 236000 233096
rect 115164 233056 236000 233084
rect 115164 233044 115170 233056
rect 235994 233044 236000 233056
rect 236052 233044 236058 233096
rect 395338 233044 395344 233096
rect 395396 233084 395402 233096
rect 579614 233084 579620 233096
rect 395396 233056 579620 233084
rect 395396 233044 395402 233056
rect 579614 233044 579620 233056
rect 579672 233044 579678 233096
rect 171962 232976 171968 233028
rect 172020 233016 172026 233028
rect 271138 233016 271144 233028
rect 172020 232988 271144 233016
rect 172020 232976 172026 232988
rect 271138 232976 271144 232988
rect 271196 232976 271202 233028
rect 278774 232636 278780 232688
rect 278832 232676 278838 232688
rect 294230 232676 294236 232688
rect 278832 232648 294236 232676
rect 278832 232636 278838 232648
rect 294230 232636 294236 232648
rect 294288 232636 294294 232688
rect 274634 232568 274640 232620
rect 274692 232608 274698 232620
rect 293218 232608 293224 232620
rect 274692 232580 293224 232608
rect 274692 232568 274698 232580
rect 293218 232568 293224 232580
rect 293276 232568 293282 232620
rect 68646 232500 68652 232552
rect 68704 232540 68710 232552
rect 328546 232540 328552 232552
rect 68704 232512 328552 232540
rect 68704 232500 68710 232512
rect 328546 232500 328552 232512
rect 328604 232500 328610 232552
rect 84102 231820 84108 231872
rect 84160 231860 84166 231872
rect 84838 231860 84844 231872
rect 84160 231832 84844 231860
rect 84160 231820 84166 231832
rect 84838 231820 84844 231832
rect 84896 231820 84902 231872
rect 61838 231752 61844 231804
rect 61896 231792 61902 231804
rect 302418 231792 302424 231804
rect 61896 231764 302424 231792
rect 61896 231752 61902 231764
rect 302418 231752 302424 231764
rect 302476 231752 302482 231804
rect 83550 231684 83556 231736
rect 83608 231724 83614 231736
rect 130378 231724 130384 231736
rect 83608 231696 130384 231724
rect 83608 231684 83614 231696
rect 130378 231684 130384 231696
rect 130436 231684 130442 231736
rect 179874 231684 179880 231736
rect 179932 231724 179938 231736
rect 295426 231724 295432 231736
rect 179932 231696 295432 231724
rect 179932 231684 179938 231696
rect 295426 231684 295432 231696
rect 295484 231684 295490 231736
rect 118326 231616 118332 231668
rect 118384 231656 118390 231668
rect 224126 231656 224132 231668
rect 118384 231628 224132 231656
rect 118384 231616 118390 231628
rect 224126 231616 224132 231628
rect 224184 231616 224190 231668
rect 167822 231072 167828 231124
rect 167880 231112 167886 231124
rect 224218 231112 224224 231124
rect 167880 231084 224224 231112
rect 167880 231072 167886 231084
rect 224218 231072 224224 231084
rect 224276 231072 224282 231124
rect 319438 231072 319444 231124
rect 319496 231112 319502 231124
rect 333974 231112 333980 231124
rect 319496 231084 333980 231112
rect 319496 231072 319502 231084
rect 333974 231072 333980 231084
rect 334032 231072 334038 231124
rect 54846 230392 54852 230444
rect 54904 230432 54910 230444
rect 289906 230432 289912 230444
rect 54904 230404 289912 230432
rect 54904 230392 54910 230404
rect 289906 230392 289912 230404
rect 289964 230392 289970 230444
rect 104710 230324 104716 230376
rect 104768 230364 104774 230376
rect 293126 230364 293132 230376
rect 104768 230336 293132 230364
rect 104768 230324 104774 230336
rect 293126 230324 293132 230336
rect 293184 230324 293190 230376
rect 98362 230256 98368 230308
rect 98420 230296 98426 230308
rect 233878 230296 233884 230308
rect 98420 230268 233884 230296
rect 98420 230256 98426 230268
rect 233878 230256 233884 230268
rect 233936 230256 233942 230308
rect 170674 229712 170680 229764
rect 170732 229752 170738 229764
rect 264330 229752 264336 229764
rect 170732 229724 264336 229752
rect 170732 229712 170738 229724
rect 264330 229712 264336 229724
rect 264388 229712 264394 229764
rect 73154 229304 73160 229356
rect 73212 229344 73218 229356
rect 73890 229344 73896 229356
rect 73212 229316 73896 229344
rect 73212 229304 73218 229316
rect 73890 229304 73896 229316
rect 73948 229304 73954 229356
rect 81526 229032 81532 229084
rect 81584 229072 81590 229084
rect 277394 229072 277400 229084
rect 81584 229044 277400 229072
rect 81584 229032 81590 229044
rect 277394 229032 277400 229044
rect 277452 229032 277458 229084
rect 57606 228964 57612 229016
rect 57664 229004 57670 229016
rect 241514 229004 241520 229016
rect 57664 228976 241520 229004
rect 57664 228964 57670 228976
rect 241514 228964 241520 228976
rect 241572 228964 241578 229016
rect 100294 228488 100300 228540
rect 100352 228528 100358 228540
rect 163682 228528 163688 228540
rect 100352 228500 163688 228528
rect 100352 228488 100358 228500
rect 163682 228488 163688 228500
rect 163740 228488 163746 228540
rect 165062 228488 165068 228540
rect 165120 228528 165126 228540
rect 206278 228528 206284 228540
rect 165120 228500 206284 228528
rect 165120 228488 165126 228500
rect 206278 228488 206284 228500
rect 206336 228488 206342 228540
rect 108666 228420 108672 228472
rect 108724 228460 108730 228472
rect 328454 228460 328460 228472
rect 108724 228432 328460 228460
rect 108724 228420 108730 228432
rect 328454 228420 328460 228432
rect 328512 228420 328518 228472
rect 67358 228352 67364 228404
rect 67416 228392 67422 228404
rect 98638 228392 98644 228404
rect 67416 228364 98644 228392
rect 67416 228352 67422 228364
rect 98638 228352 98644 228364
rect 98696 228352 98702 228404
rect 162670 228352 162676 228404
rect 162728 228392 162734 228404
rect 582374 228392 582380 228404
rect 162728 228364 582380 228392
rect 162728 228352 162734 228364
rect 582374 228352 582380 228364
rect 582432 228352 582438 228404
rect 86218 227672 86224 227724
rect 86276 227712 86282 227724
rect 302234 227712 302240 227724
rect 86276 227684 302240 227712
rect 86276 227672 86282 227684
rect 302234 227672 302240 227684
rect 302292 227672 302298 227724
rect 92566 227128 92572 227180
rect 92624 227168 92630 227180
rect 220078 227168 220084 227180
rect 92624 227140 220084 227168
rect 92624 227128 92630 227140
rect 220078 227128 220084 227140
rect 220136 227128 220142 227180
rect 280154 227128 280160 227180
rect 280212 227168 280218 227180
rect 311894 227168 311900 227180
rect 280212 227140 311900 227168
rect 280212 227128 280218 227140
rect 311894 227128 311900 227140
rect 311952 227128 311958 227180
rect 113174 227060 113180 227112
rect 113232 227100 113238 227112
rect 283558 227100 283564 227112
rect 113232 227072 283564 227100
rect 113232 227060 113238 227072
rect 283558 227060 283564 227072
rect 283616 227060 283622 227112
rect 66070 226992 66076 227044
rect 66128 227032 66134 227044
rect 324590 227032 324596 227044
rect 66128 227004 324596 227032
rect 66128 226992 66134 227004
rect 324590 226992 324596 227004
rect 324648 226992 324654 227044
rect 155494 226244 155500 226296
rect 155552 226284 155558 226296
rect 296898 226284 296904 226296
rect 155552 226256 296904 226284
rect 155552 226244 155558 226256
rect 296898 226244 296904 226256
rect 296956 226244 296962 226296
rect 182818 225700 182824 225752
rect 182876 225740 182882 225752
rect 319438 225740 319444 225752
rect 182876 225712 319444 225740
rect 182876 225700 182882 225712
rect 319438 225700 319444 225712
rect 319496 225700 319502 225752
rect 156782 225632 156788 225684
rect 156840 225672 156846 225684
rect 336734 225672 336740 225684
rect 156840 225644 336740 225672
rect 156840 225632 156846 225644
rect 336734 225632 336740 225644
rect 336792 225632 336798 225684
rect 67266 225564 67272 225616
rect 67324 225604 67330 225616
rect 253198 225604 253204 225616
rect 67324 225576 253204 225604
rect 67324 225564 67330 225576
rect 253198 225564 253204 225576
rect 253256 225564 253262 225616
rect 81434 224884 81440 224936
rect 81492 224924 81498 224936
rect 278866 224924 278872 224936
rect 81492 224896 278872 224924
rect 81492 224884 81498 224896
rect 278866 224884 278872 224896
rect 278924 224884 278930 224936
rect 147214 224816 147220 224868
rect 147272 224856 147278 224868
rect 299658 224856 299664 224868
rect 147272 224828 299664 224856
rect 147272 224816 147278 224828
rect 299658 224816 299664 224828
rect 299716 224816 299722 224868
rect 129274 224340 129280 224392
rect 129332 224380 129338 224392
rect 257338 224380 257344 224392
rect 129332 224352 257344 224380
rect 129332 224340 129338 224352
rect 257338 224340 257344 224352
rect 257396 224340 257402 224392
rect 97074 224272 97080 224324
rect 97132 224312 97138 224324
rect 129182 224312 129188 224324
rect 97132 224284 129188 224312
rect 97132 224272 97138 224284
rect 129182 224272 129188 224284
rect 129240 224272 129246 224324
rect 164970 224272 164976 224324
rect 165028 224312 165034 224324
rect 311158 224312 311164 224324
rect 165028 224284 311164 224312
rect 165028 224272 165034 224284
rect 311158 224272 311164 224284
rect 311216 224272 311222 224324
rect 3602 224204 3608 224256
rect 3660 224244 3666 224256
rect 120166 224244 120172 224256
rect 3660 224216 120172 224244
rect 3660 224204 3666 224216
rect 120166 224204 120172 224216
rect 120224 224204 120230 224256
rect 136082 224204 136088 224256
rect 136140 224244 136146 224256
rect 580350 224244 580356 224256
rect 136140 224216 580356 224244
rect 136140 224204 136146 224216
rect 580350 224204 580356 224216
rect 580408 224204 580414 224256
rect 160922 223524 160928 223576
rect 160980 223564 160986 223576
rect 574738 223564 574744 223576
rect 160980 223536 574744 223564
rect 160980 223524 160986 223536
rect 574738 223524 574744 223536
rect 574796 223524 574802 223576
rect 69106 222980 69112 223032
rect 69164 223020 69170 223032
rect 249794 223020 249800 223032
rect 69164 222992 249800 223020
rect 69164 222980 69170 222992
rect 249794 222980 249800 222992
rect 249852 222980 249858 223032
rect 56410 222912 56416 222964
rect 56468 222952 56474 222964
rect 240778 222952 240784 222964
rect 56468 222924 240784 222952
rect 56468 222912 56474 222924
rect 240778 222912 240784 222924
rect 240836 222912 240842 222964
rect 256694 222912 256700 222964
rect 256752 222952 256758 222964
rect 278038 222952 278044 222964
rect 256752 222924 278044 222952
rect 256752 222912 256758 222924
rect 278038 222912 278044 222924
rect 278096 222912 278102 222964
rect 131850 222844 131856 222896
rect 131908 222884 131914 222896
rect 345014 222884 345020 222896
rect 131908 222856 345020 222884
rect 131908 222844 131914 222856
rect 345014 222844 345020 222856
rect 345072 222844 345078 222896
rect 162210 221620 162216 221672
rect 162268 221660 162274 221672
rect 214558 221660 214564 221672
rect 162268 221632 214564 221660
rect 162268 221620 162274 221632
rect 214558 221620 214564 221632
rect 214616 221620 214622 221672
rect 88058 221552 88064 221604
rect 88116 221592 88122 221604
rect 247678 221592 247684 221604
rect 88116 221564 247684 221592
rect 88116 221552 88122 221564
rect 247678 221552 247684 221564
rect 247736 221552 247742 221604
rect 64690 221484 64696 221536
rect 64748 221524 64754 221536
rect 324406 221524 324412 221536
rect 64748 221496 324412 221524
rect 64748 221484 64754 221496
rect 324406 221484 324412 221496
rect 324464 221484 324470 221536
rect 77754 221416 77760 221468
rect 77812 221456 77818 221468
rect 351914 221456 351920 221468
rect 77812 221428 351920 221456
rect 77812 221416 77818 221428
rect 351914 221416 351920 221428
rect 351972 221416 351978 221468
rect 111886 220328 111892 220380
rect 111944 220368 111950 220380
rect 267734 220368 267740 220380
rect 111944 220340 267740 220368
rect 111944 220328 111950 220340
rect 267734 220328 267740 220340
rect 267792 220328 267798 220380
rect 79042 220260 79048 220312
rect 79100 220300 79106 220312
rect 242158 220300 242164 220312
rect 79100 220272 242164 220300
rect 79100 220260 79106 220272
rect 242158 220260 242164 220272
rect 242216 220260 242222 220312
rect 159358 220192 159364 220244
rect 159416 220232 159422 220244
rect 346486 220232 346492 220244
rect 159416 220204 346492 220232
rect 159416 220192 159422 220204
rect 346486 220192 346492 220204
rect 346544 220192 346550 220244
rect 56318 220124 56324 220176
rect 56376 220164 56382 220176
rect 313918 220164 313924 220176
rect 56376 220136 313924 220164
rect 56376 220124 56382 220136
rect 313918 220124 313924 220136
rect 313976 220124 313982 220176
rect 179046 220056 179052 220108
rect 179104 220096 179110 220108
rect 580442 220096 580448 220108
rect 179104 220068 580448 220096
rect 179104 220056 179110 220068
rect 580442 220056 580448 220068
rect 580500 220056 580506 220108
rect 76006 219376 76012 219428
rect 76064 219416 76070 219428
rect 150342 219416 150348 219428
rect 76064 219388 150348 219416
rect 76064 219376 76070 219388
rect 150342 219376 150348 219388
rect 150400 219376 150406 219428
rect 471238 219376 471244 219428
rect 471296 219416 471302 219428
rect 580166 219416 580172 219428
rect 471296 219388 580172 219416
rect 471296 219376 471302 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 170398 218968 170404 219020
rect 170456 219008 170462 219020
rect 273346 219008 273352 219020
rect 170456 218980 273352 219008
rect 170456 218968 170462 218980
rect 273346 218968 273352 218980
rect 273404 218968 273410 219020
rect 153930 218900 153936 218952
rect 153988 218940 153994 218952
rect 318058 218940 318064 218952
rect 153988 218912 318064 218940
rect 153988 218900 153994 218912
rect 318058 218900 318064 218912
rect 318116 218900 318122 218952
rect 65978 218832 65984 218884
rect 66036 218872 66042 218884
rect 278866 218872 278872 218884
rect 66036 218844 278872 218872
rect 66036 218832 66042 218844
rect 278866 218832 278872 218844
rect 278924 218832 278930 218884
rect 48222 218764 48228 218816
rect 48280 218804 48286 218816
rect 343634 218804 343640 218816
rect 48280 218776 343640 218804
rect 48280 218764 48286 218776
rect 343634 218764 343640 218776
rect 343692 218764 343698 218816
rect 150342 218696 150348 218748
rect 150400 218736 150406 218748
rect 582466 218736 582472 218748
rect 150400 218708 582472 218736
rect 150400 218696 150406 218708
rect 582466 218696 582472 218708
rect 582524 218696 582530 218748
rect 145650 217540 145656 217592
rect 145708 217580 145714 217592
rect 266446 217580 266452 217592
rect 145708 217552 266452 217580
rect 145708 217540 145714 217552
rect 266446 217540 266452 217552
rect 266504 217540 266510 217592
rect 148594 217472 148600 217524
rect 148652 217512 148658 217524
rect 270494 217512 270500 217524
rect 148652 217484 270500 217512
rect 148652 217472 148658 217484
rect 270494 217472 270500 217484
rect 270552 217472 270558 217524
rect 138750 217404 138756 217456
rect 138808 217444 138814 217456
rect 274726 217444 274732 217456
rect 138808 217416 274732 217444
rect 138808 217404 138814 217416
rect 274726 217404 274732 217416
rect 274784 217404 274790 217456
rect 106918 217336 106924 217388
rect 106976 217376 106982 217388
rect 160738 217376 160744 217388
rect 106976 217348 160744 217376
rect 106976 217336 106982 217348
rect 160738 217336 160744 217348
rect 160796 217336 160802 217388
rect 160830 217336 160836 217388
rect 160888 217376 160894 217388
rect 356054 217376 356060 217388
rect 160888 217348 356060 217376
rect 160888 217336 160894 217348
rect 356054 217336 356060 217348
rect 356112 217336 356118 217388
rect 102226 217268 102232 217320
rect 102284 217308 102290 217320
rect 319530 217308 319536 217320
rect 102284 217280 319536 217308
rect 102284 217268 102290 217280
rect 319530 217268 319536 217280
rect 319588 217268 319594 217320
rect 100846 216112 100852 216164
rect 100904 216152 100910 216164
rect 255314 216152 255320 216164
rect 100904 216124 255320 216152
rect 100904 216112 100910 216124
rect 255314 216112 255320 216124
rect 255372 216112 255378 216164
rect 159542 216044 159548 216096
rect 159600 216084 159606 216096
rect 345106 216084 345112 216096
rect 159600 216056 345112 216084
rect 159600 216044 159606 216056
rect 345106 216044 345112 216056
rect 345164 216044 345170 216096
rect 116578 215976 116584 216028
rect 116636 216016 116642 216028
rect 315390 216016 315396 216028
rect 116636 215988 315396 216016
rect 116636 215976 116642 215988
rect 315390 215976 315396 215988
rect 315448 215976 315454 216028
rect 134794 215908 134800 215960
rect 134852 215948 134858 215960
rect 338114 215948 338120 215960
rect 134852 215920 338120 215948
rect 134852 215908 134858 215920
rect 338114 215908 338120 215920
rect 338172 215908 338178 215960
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 21358 215268 21364 215280
rect 3384 215240 21364 215268
rect 3384 215228 3390 215240
rect 21358 215228 21364 215240
rect 21416 215228 21422 215280
rect 258074 215024 258080 215076
rect 258132 215064 258138 215076
rect 264238 215064 264244 215076
rect 258132 215036 264244 215064
rect 258132 215024 258138 215036
rect 264238 215024 264244 215036
rect 264296 215024 264302 215076
rect 144270 214752 144276 214804
rect 144328 214792 144334 214804
rect 210418 214792 210424 214804
rect 144328 214764 210424 214792
rect 144328 214752 144334 214764
rect 210418 214752 210424 214764
rect 210476 214752 210482 214804
rect 163682 214684 163688 214736
rect 163740 214724 163746 214736
rect 276014 214724 276020 214736
rect 163740 214696 276020 214724
rect 163740 214684 163746 214696
rect 276014 214684 276020 214696
rect 276072 214684 276078 214736
rect 114554 214616 114560 214668
rect 114612 214656 114618 214668
rect 325694 214656 325700 214668
rect 114612 214628 325700 214656
rect 114612 214616 114618 214628
rect 325694 214616 325700 214628
rect 325752 214616 325758 214668
rect 46842 214548 46848 214600
rect 46900 214588 46906 214600
rect 311250 214588 311256 214600
rect 46900 214560 311256 214588
rect 46900 214548 46906 214560
rect 311250 214548 311256 214560
rect 311308 214548 311314 214600
rect 255958 213868 255964 213920
rect 256016 213908 256022 213920
rect 258718 213908 258724 213920
rect 256016 213880 258724 213908
rect 256016 213868 256022 213880
rect 258718 213868 258724 213880
rect 258776 213868 258782 213920
rect 152734 213392 152740 213444
rect 152792 213432 152798 213444
rect 236638 213432 236644 213444
rect 152792 213404 236644 213432
rect 152792 213392 152798 213404
rect 236638 213392 236644 213404
rect 236696 213392 236702 213444
rect 149698 213324 149704 213376
rect 149756 213364 149762 213376
rect 277394 213364 277400 213376
rect 149756 213336 277400 213364
rect 149756 213324 149762 213336
rect 277394 213324 277400 213336
rect 277452 213324 277458 213376
rect 99374 213256 99380 213308
rect 99432 213296 99438 213308
rect 325878 213296 325884 213308
rect 99432 213268 325884 213296
rect 99432 213256 99438 213268
rect 325878 213256 325884 213268
rect 325936 213256 325942 213308
rect 86954 213188 86960 213240
rect 87012 213228 87018 213240
rect 322934 213228 322940 213240
rect 87012 213200 322940 213228
rect 87012 213188 87018 213200
rect 322934 213188 322940 213200
rect 322992 213188 322998 213240
rect 124950 211896 124956 211948
rect 125008 211936 125014 211948
rect 273254 211936 273260 211948
rect 125008 211908 273260 211936
rect 125008 211896 125014 211908
rect 273254 211896 273260 211908
rect 273312 211896 273318 211948
rect 89806 211828 89812 211880
rect 89864 211868 89870 211880
rect 274818 211868 274824 211880
rect 89864 211840 274824 211868
rect 89864 211828 89870 211840
rect 274818 211828 274824 211840
rect 274876 211828 274882 211880
rect 61746 211760 61752 211812
rect 61804 211800 61810 211812
rect 259454 211800 259460 211812
rect 61804 211772 259460 211800
rect 61804 211760 61810 211772
rect 259454 211760 259460 211772
rect 259512 211760 259518 211812
rect 260098 211760 260104 211812
rect 260156 211800 260162 211812
rect 332594 211800 332600 211812
rect 260156 211772 332600 211800
rect 260156 211760 260162 211772
rect 332594 211760 332600 211772
rect 332652 211760 332658 211812
rect 231854 210604 231860 210656
rect 231912 210644 231918 210656
rect 282914 210644 282920 210656
rect 231912 210616 282920 210644
rect 231912 210604 231918 210616
rect 282914 210604 282920 210616
rect 282972 210604 282978 210656
rect 133230 210536 133236 210588
rect 133288 210576 133294 210588
rect 232498 210576 232504 210588
rect 133288 210548 232504 210576
rect 133288 210536 133294 210548
rect 232498 210536 232504 210548
rect 232556 210536 232562 210588
rect 4798 210468 4804 210520
rect 4856 210508 4862 210520
rect 83458 210508 83464 210520
rect 4856 210480 83464 210508
rect 4856 210468 4862 210480
rect 83458 210468 83464 210480
rect 83516 210468 83522 210520
rect 144546 210468 144552 210520
rect 144604 210508 144610 210520
rect 246390 210508 246396 210520
rect 144604 210480 246396 210508
rect 144604 210468 144610 210480
rect 246390 210468 246396 210480
rect 246448 210468 246454 210520
rect 74626 210400 74632 210452
rect 74684 210440 74690 210452
rect 246298 210440 246304 210452
rect 74684 210412 246304 210440
rect 74684 210400 74690 210412
rect 246298 210400 246304 210412
rect 246356 210400 246362 210452
rect 271874 210400 271880 210452
rect 271932 210440 271938 210452
rect 294046 210440 294052 210452
rect 271932 210412 294052 210440
rect 271932 210400 271938 210412
rect 294046 210400 294052 210412
rect 294104 210400 294110 210452
rect 138842 209176 138848 209228
rect 138900 209216 138906 209228
rect 258166 209216 258172 209228
rect 138900 209188 258172 209216
rect 138900 209176 138906 209188
rect 258166 209176 258172 209188
rect 258224 209176 258230 209228
rect 67450 209108 67456 209160
rect 67508 209148 67514 209160
rect 247770 209148 247776 209160
rect 67508 209120 247776 209148
rect 67508 209108 67514 209120
rect 247770 209108 247776 209120
rect 247828 209108 247834 209160
rect 103698 209040 103704 209092
rect 103756 209080 103762 209092
rect 327074 209080 327080 209092
rect 103756 209052 327080 209080
rect 103756 209040 103762 209052
rect 327074 209040 327080 209052
rect 327132 209040 327138 209092
rect 237374 207952 237380 208004
rect 237432 207992 237438 208004
rect 279418 207992 279424 208004
rect 237432 207964 279424 207992
rect 237432 207952 237438 207964
rect 279418 207952 279424 207964
rect 279476 207952 279482 208004
rect 197998 207884 198004 207936
rect 198056 207924 198062 207936
rect 305638 207924 305644 207936
rect 198056 207896 305644 207924
rect 198056 207884 198062 207896
rect 305638 207884 305644 207896
rect 305696 207884 305702 207936
rect 151170 207816 151176 207868
rect 151228 207856 151234 207868
rect 281626 207856 281632 207868
rect 151228 207828 281632 207856
rect 151228 207816 151234 207828
rect 281626 207816 281632 207828
rect 281684 207816 281690 207868
rect 55030 207748 55036 207800
rect 55088 207788 55094 207800
rect 239398 207788 239404 207800
rect 55088 207760 239404 207788
rect 55088 207748 55094 207760
rect 239398 207748 239404 207760
rect 239456 207748 239462 207800
rect 126422 207680 126428 207732
rect 126480 207720 126486 207732
rect 339678 207720 339684 207732
rect 126480 207692 339684 207720
rect 126480 207680 126486 207692
rect 339678 207680 339684 207692
rect 339736 207680 339742 207732
rect 53650 207612 53656 207664
rect 53708 207652 53714 207664
rect 271966 207652 271972 207664
rect 53708 207624 271972 207652
rect 53708 207612 53714 207624
rect 271966 207612 271972 207624
rect 272024 207612 272030 207664
rect 281534 207612 281540 207664
rect 281592 207652 281598 207664
rect 342254 207652 342260 207664
rect 281592 207624 342260 207652
rect 281592 207612 281598 207624
rect 342254 207612 342260 207624
rect 342312 207612 342318 207664
rect 45370 206388 45376 206440
rect 45428 206428 45434 206440
rect 228358 206428 228364 206440
rect 45428 206400 228364 206428
rect 45428 206388 45434 206400
rect 228358 206388 228364 206400
rect 228416 206388 228422 206440
rect 260834 206388 260840 206440
rect 260892 206428 260898 206440
rect 289078 206428 289084 206440
rect 260892 206400 289084 206428
rect 260892 206388 260898 206400
rect 289078 206388 289084 206400
rect 289136 206388 289142 206440
rect 160738 206320 160744 206372
rect 160796 206360 160802 206372
rect 347774 206360 347780 206372
rect 160796 206332 347780 206360
rect 160796 206320 160802 206332
rect 347774 206320 347780 206332
rect 347832 206320 347838 206372
rect 75914 206252 75920 206304
rect 75972 206292 75978 206304
rect 327166 206292 327172 206304
rect 75972 206264 327172 206292
rect 75972 206252 75978 206264
rect 327166 206252 327172 206264
rect 327224 206252 327230 206304
rect 94038 205164 94044 205216
rect 94096 205204 94102 205216
rect 189902 205204 189908 205216
rect 94096 205176 189908 205204
rect 94096 205164 94102 205176
rect 189902 205164 189908 205176
rect 189960 205164 189966 205216
rect 189718 205096 189724 205148
rect 189776 205136 189782 205148
rect 339494 205136 339500 205148
rect 189776 205108 339500 205136
rect 189776 205096 189782 205108
rect 339494 205096 339500 205108
rect 339552 205096 339558 205148
rect 70394 205028 70400 205080
rect 70452 205068 70458 205080
rect 252830 205068 252836 205080
rect 70452 205040 252836 205068
rect 70452 205028 70458 205040
rect 252830 205028 252836 205040
rect 252888 205028 252894 205080
rect 59170 204960 59176 205012
rect 59228 205000 59234 205012
rect 259546 205000 259552 205012
rect 59228 204972 259552 205000
rect 59228 204960 59234 204972
rect 259546 204960 259552 204972
rect 259604 204960 259610 205012
rect 118694 204892 118700 204944
rect 118752 204932 118758 204944
rect 328638 204932 328644 204944
rect 118752 204904 328644 204932
rect 118752 204892 118758 204904
rect 328638 204892 328644 204904
rect 328696 204892 328702 204944
rect 153838 203804 153844 203856
rect 153896 203844 153902 203856
rect 243538 203844 243544 203856
rect 153896 203816 243544 203844
rect 153896 203804 153902 203816
rect 243538 203804 243544 203816
rect 243596 203804 243602 203856
rect 248414 203804 248420 203856
rect 248472 203844 248478 203856
rect 291194 203844 291200 203856
rect 248472 203816 291200 203844
rect 248472 203804 248478 203816
rect 291194 203804 291200 203816
rect 291252 203804 291258 203856
rect 166534 203736 166540 203788
rect 166592 203776 166598 203788
rect 342438 203776 342444 203788
rect 166592 203748 342444 203776
rect 166592 203736 166598 203748
rect 342438 203736 342444 203748
rect 342496 203736 342502 203788
rect 122098 203668 122104 203720
rect 122156 203708 122162 203720
rect 325786 203708 325792 203720
rect 122156 203680 325792 203708
rect 122156 203668 122162 203680
rect 325786 203668 325792 203680
rect 325844 203668 325850 203720
rect 57698 203600 57704 203652
rect 57756 203640 57762 203652
rect 273438 203640 273444 203652
rect 57756 203612 273444 203640
rect 57756 203600 57762 203612
rect 273438 203600 273444 203612
rect 273496 203600 273502 203652
rect 71774 203532 71780 203584
rect 71832 203572 71838 203584
rect 327258 203572 327264 203584
rect 71832 203544 327264 203572
rect 71832 203532 71838 203544
rect 327258 203532 327264 203544
rect 327316 203532 327322 203584
rect 245654 202444 245660 202496
rect 245712 202484 245718 202496
rect 308582 202484 308588 202496
rect 245712 202456 308588 202484
rect 245712 202444 245718 202456
rect 308582 202444 308588 202456
rect 308640 202444 308646 202496
rect 146938 202376 146944 202428
rect 146996 202416 147002 202428
rect 281534 202416 281540 202428
rect 146996 202388 281540 202416
rect 146996 202376 147002 202388
rect 281534 202376 281540 202388
rect 281592 202376 281598 202428
rect 102134 202308 102140 202360
rect 102192 202348 102198 202360
rect 252646 202348 252652 202360
rect 102192 202320 252652 202348
rect 102192 202308 102198 202320
rect 252646 202308 252652 202320
rect 252704 202308 252710 202360
rect 160002 202240 160008 202292
rect 160060 202280 160066 202292
rect 354674 202280 354680 202292
rect 160060 202252 354680 202280
rect 160060 202240 160066 202252
rect 354674 202240 354680 202252
rect 354732 202240 354738 202292
rect 145558 202172 145564 202224
rect 145616 202212 145622 202224
rect 343726 202212 343732 202224
rect 145616 202184 343732 202212
rect 145616 202172 145622 202184
rect 343726 202172 343732 202184
rect 343784 202172 343790 202224
rect 60550 202104 60556 202156
rect 60608 202144 60614 202156
rect 276106 202144 276112 202156
rect 60608 202116 276112 202144
rect 60608 202104 60614 202116
rect 276106 202104 276112 202116
rect 276164 202104 276170 202156
rect 131758 200812 131764 200864
rect 131816 200852 131822 200864
rect 258258 200852 258264 200864
rect 131816 200824 258264 200852
rect 131816 200812 131822 200824
rect 258258 200812 258264 200824
rect 258316 200812 258322 200864
rect 56502 200744 56508 200796
rect 56560 200784 56566 200796
rect 231118 200784 231124 200796
rect 56560 200756 231124 200784
rect 56560 200744 56566 200756
rect 231118 200744 231124 200756
rect 231176 200744 231182 200796
rect 142890 199520 142896 199572
rect 142948 199560 142954 199572
rect 269114 199560 269120 199572
rect 142948 199532 269120 199560
rect 142948 199520 142954 199532
rect 269114 199520 269120 199532
rect 269172 199520 269178 199572
rect 162302 199452 162308 199504
rect 162360 199492 162366 199504
rect 342346 199492 342352 199504
rect 162360 199464 342352 199492
rect 162360 199452 162366 199464
rect 342346 199452 342352 199464
rect 342404 199452 342410 199504
rect 96522 199384 96528 199436
rect 96580 199424 96586 199436
rect 582374 199424 582380 199436
rect 96580 199396 582380 199424
rect 96580 199384 96586 199396
rect 582374 199384 582380 199396
rect 582432 199384 582438 199436
rect 126330 198160 126336 198212
rect 126388 198200 126394 198212
rect 239490 198200 239496 198212
rect 126388 198172 239496 198200
rect 126388 198160 126394 198172
rect 239490 198160 239496 198172
rect 239548 198160 239554 198212
rect 140314 198092 140320 198144
rect 140372 198132 140378 198144
rect 264974 198132 264980 198144
rect 140372 198104 264980 198132
rect 140372 198092 140378 198104
rect 264974 198092 264980 198104
rect 265032 198092 265038 198144
rect 115934 198024 115940 198076
rect 115992 198064 115998 198076
rect 260926 198064 260932 198076
rect 115992 198036 260932 198064
rect 115992 198024 115998 198036
rect 260926 198024 260932 198036
rect 260984 198024 260990 198076
rect 151078 197956 151084 198008
rect 151136 197996 151142 198008
rect 319622 197996 319628 198008
rect 151136 197968 319628 197996
rect 151136 197956 151142 197968
rect 319622 197956 319628 197968
rect 319680 197956 319686 198008
rect 130654 196936 130660 196988
rect 130712 196976 130718 196988
rect 250070 196976 250076 196988
rect 130712 196948 250076 196976
rect 130712 196936 130718 196948
rect 250070 196936 250076 196948
rect 250128 196936 250134 196988
rect 192478 196868 192484 196920
rect 192536 196908 192542 196920
rect 312538 196908 312544 196920
rect 192536 196880 312544 196908
rect 192536 196868 192542 196880
rect 312538 196868 312544 196880
rect 312596 196868 312602 196920
rect 66162 196800 66168 196852
rect 66220 196840 66226 196852
rect 251174 196840 251180 196852
rect 66220 196812 251180 196840
rect 66220 196800 66226 196812
rect 251174 196800 251180 196812
rect 251232 196800 251238 196852
rect 123478 196732 123484 196784
rect 123536 196772 123542 196784
rect 349338 196772 349344 196784
rect 123536 196744 349344 196772
rect 123536 196732 123542 196744
rect 349338 196732 349344 196744
rect 349396 196732 349402 196784
rect 69658 196664 69664 196716
rect 69716 196704 69722 196716
rect 320818 196704 320824 196716
rect 69716 196676 320824 196704
rect 69716 196664 69722 196676
rect 320818 196664 320824 196676
rect 320876 196664 320882 196716
rect 50890 196596 50896 196648
rect 50948 196636 50954 196648
rect 334158 196636 334164 196648
rect 50948 196608 334164 196636
rect 50948 196596 50954 196608
rect 334158 196596 334164 196608
rect 334216 196596 334222 196648
rect 134610 195508 134616 195560
rect 134668 195548 134674 195560
rect 267826 195548 267832 195560
rect 134668 195520 267832 195548
rect 134668 195508 134674 195520
rect 267826 195508 267832 195520
rect 267884 195508 267890 195560
rect 89714 195440 89720 195492
rect 89772 195480 89778 195492
rect 263594 195480 263600 195492
rect 89772 195452 263600 195480
rect 89772 195440 89778 195452
rect 263594 195440 263600 195452
rect 263652 195440 263658 195492
rect 158070 195372 158076 195424
rect 158128 195412 158134 195424
rect 347866 195412 347872 195424
rect 158128 195384 347872 195412
rect 158128 195372 158134 195384
rect 347866 195372 347872 195384
rect 347924 195372 347930 195424
rect 104894 195304 104900 195356
rect 104952 195344 104958 195356
rect 336826 195344 336832 195356
rect 104952 195316 336832 195344
rect 104952 195304 104958 195316
rect 336826 195304 336832 195316
rect 336884 195304 336890 195356
rect 92474 195236 92480 195288
rect 92532 195276 92538 195288
rect 328730 195276 328736 195288
rect 92532 195248 328736 195276
rect 92532 195236 92538 195248
rect 328730 195236 328736 195248
rect 328788 195236 328794 195288
rect 196710 194148 196716 194200
rect 196768 194188 196774 194200
rect 244918 194188 244924 194200
rect 196768 194160 244924 194188
rect 196768 194148 196774 194160
rect 244918 194148 244924 194160
rect 244976 194148 244982 194200
rect 253198 194148 253204 194200
rect 253256 194188 253262 194200
rect 329926 194188 329932 194200
rect 253256 194160 329932 194188
rect 253256 194148 253262 194160
rect 329926 194148 329932 194160
rect 329984 194148 329990 194200
rect 129182 194080 129188 194132
rect 129240 194120 129246 194132
rect 262398 194120 262404 194132
rect 129240 194092 262404 194120
rect 129240 194080 129246 194092
rect 262398 194080 262404 194092
rect 262456 194080 262462 194132
rect 167730 194012 167736 194064
rect 167788 194052 167794 194064
rect 318150 194052 318156 194064
rect 167788 194024 318156 194052
rect 167788 194012 167794 194024
rect 318150 194012 318156 194024
rect 318208 194012 318214 194064
rect 147122 193944 147128 193996
rect 147180 193984 147186 193996
rect 331306 193984 331312 193996
rect 147180 193956 331312 193984
rect 147180 193944 147186 193956
rect 331306 193944 331312 193956
rect 331364 193944 331370 193996
rect 44082 193876 44088 193928
rect 44140 193916 44146 193928
rect 270586 193916 270592 193928
rect 44140 193888 270592 193916
rect 44140 193876 44146 193888
rect 270586 193876 270592 193888
rect 270644 193876 270650 193928
rect 96614 193808 96620 193860
rect 96672 193848 96678 193860
rect 331214 193848 331220 193860
rect 96672 193820 331220 193848
rect 96672 193808 96678 193820
rect 331214 193808 331220 193820
rect 331272 193808 331278 193860
rect 127618 192584 127624 192636
rect 127676 192624 127682 192636
rect 272058 192624 272064 192636
rect 127676 192596 272064 192624
rect 127676 192584 127682 192596
rect 272058 192584 272064 192596
rect 272116 192584 272122 192636
rect 93946 192516 93952 192568
rect 94004 192556 94010 192568
rect 254118 192556 254124 192568
rect 94004 192528 254124 192556
rect 94004 192516 94010 192528
rect 254118 192516 254124 192528
rect 254176 192516 254182 192568
rect 133138 192448 133144 192500
rect 133196 192488 133202 192500
rect 341058 192488 341064 192500
rect 133196 192460 341064 192488
rect 133196 192448 133202 192460
rect 341058 192448 341064 192460
rect 341116 192448 341122 192500
rect 142982 191360 142988 191412
rect 143040 191400 143046 191412
rect 242250 191400 242256 191412
rect 143040 191372 242256 191400
rect 143040 191360 143046 191372
rect 242250 191360 242256 191372
rect 242308 191360 242314 191412
rect 149790 191292 149796 191344
rect 149848 191332 149854 191344
rect 260834 191332 260840 191344
rect 149848 191304 260840 191332
rect 149848 191292 149854 191304
rect 260834 191292 260840 191304
rect 260892 191292 260898 191344
rect 137278 191224 137284 191276
rect 137336 191264 137342 191276
rect 255498 191264 255504 191276
rect 137336 191236 255504 191264
rect 137336 191224 137342 191236
rect 255498 191224 255504 191236
rect 255556 191224 255562 191276
rect 264330 191224 264336 191276
rect 264388 191264 264394 191276
rect 338206 191264 338212 191276
rect 264388 191236 338212 191264
rect 264388 191224 264394 191236
rect 338206 191224 338212 191236
rect 338264 191224 338270 191276
rect 227714 191156 227720 191208
rect 227772 191196 227778 191208
rect 346394 191196 346400 191208
rect 227772 191168 346400 191196
rect 227772 191156 227778 191168
rect 346394 191156 346400 191168
rect 346452 191156 346458 191208
rect 135898 191088 135904 191140
rect 135956 191128 135962 191140
rect 343818 191128 343824 191140
rect 135956 191100 343824 191128
rect 135956 191088 135962 191100
rect 343818 191088 343824 191100
rect 343876 191088 343882 191140
rect 102042 190476 102048 190528
rect 102100 190516 102106 190528
rect 203610 190516 203616 190528
rect 102100 190488 203616 190516
rect 102100 190476 102106 190488
rect 203610 190476 203616 190488
rect 203668 190476 203674 190528
rect 211062 190068 211068 190120
rect 211120 190108 211126 190120
rect 244274 190108 244280 190120
rect 211120 190080 244280 190108
rect 211120 190068 211126 190080
rect 244274 190068 244280 190080
rect 244332 190068 244338 190120
rect 229094 190000 229100 190052
rect 229152 190040 229158 190052
rect 268378 190040 268384 190052
rect 229152 190012 268384 190040
rect 229152 190000 229158 190012
rect 268378 190000 268384 190012
rect 268436 190000 268442 190052
rect 144454 189932 144460 189984
rect 144512 189972 144518 189984
rect 261018 189972 261024 189984
rect 144512 189944 261024 189972
rect 144512 189932 144518 189944
rect 261018 189932 261024 189944
rect 261076 189932 261082 189984
rect 141418 189864 141424 189916
rect 141476 189904 141482 189916
rect 269206 189904 269212 189916
rect 141476 189876 269212 189904
rect 141476 189864 141482 189876
rect 269206 189864 269212 189876
rect 269264 189864 269270 189916
rect 21358 189796 21364 189848
rect 21416 189836 21422 189848
rect 111058 189836 111064 189848
rect 21416 189808 111064 189836
rect 21416 189796 21422 189808
rect 111058 189796 111064 189808
rect 111116 189796 111122 189848
rect 173250 189796 173256 189848
rect 173308 189836 173314 189848
rect 324498 189836 324504 189848
rect 173308 189808 324504 189836
rect 173308 189796 173314 189808
rect 324498 189796 324504 189808
rect 324556 189796 324562 189848
rect 84286 189728 84292 189780
rect 84344 189768 84350 189780
rect 254026 189768 254032 189780
rect 84344 189740 254032 189768
rect 84344 189728 84350 189740
rect 254026 189728 254032 189740
rect 254084 189728 254090 189780
rect 257338 189728 257344 189780
rect 257396 189768 257402 189780
rect 340966 189768 340972 189780
rect 257396 189740 340972 189768
rect 257396 189728 257402 189740
rect 340966 189728 340972 189740
rect 341024 189728 341030 189780
rect 107562 189184 107568 189236
rect 107620 189224 107626 189236
rect 171870 189224 171876 189236
rect 107620 189196 171876 189224
rect 107620 189184 107626 189196
rect 171870 189184 171876 189196
rect 171928 189184 171934 189236
rect 118602 189116 118608 189168
rect 118660 189156 118666 189168
rect 189810 189156 189816 189168
rect 118660 189128 189816 189156
rect 118660 189116 118666 189128
rect 189810 189116 189816 189128
rect 189868 189116 189874 189168
rect 133782 189048 133788 189100
rect 133840 189088 133846 189100
rect 214650 189088 214656 189100
rect 133840 189060 214656 189088
rect 133840 189048 133846 189060
rect 214650 189048 214656 189060
rect 214708 189048 214714 189100
rect 3142 188980 3148 189032
rect 3200 189020 3206 189032
rect 14458 189020 14464 189032
rect 3200 188992 14464 189020
rect 3200 188980 3206 188992
rect 14458 188980 14464 188992
rect 14516 188980 14522 189032
rect 206278 188572 206284 188624
rect 206336 188612 206342 188624
rect 263686 188612 263692 188624
rect 206336 188584 263692 188612
rect 206336 188572 206342 188584
rect 263686 188572 263692 188584
rect 263744 188572 263750 188624
rect 138658 188504 138664 188556
rect 138716 188544 138722 188556
rect 258074 188544 258080 188556
rect 138716 188516 258080 188544
rect 138716 188504 138722 188516
rect 258074 188504 258080 188516
rect 258132 188504 258138 188556
rect 258718 188504 258724 188556
rect 258776 188544 258782 188556
rect 339770 188544 339776 188556
rect 258776 188516 339776 188544
rect 258776 188504 258782 188516
rect 339770 188504 339776 188516
rect 339828 188504 339834 188556
rect 135990 188436 135996 188488
rect 136048 188476 136054 188488
rect 266538 188476 266544 188488
rect 136048 188448 266544 188476
rect 136048 188436 136054 188448
rect 266538 188436 266544 188448
rect 266596 188436 266602 188488
rect 18598 188368 18604 188420
rect 18656 188408 18662 188420
rect 109034 188408 109040 188420
rect 18656 188380 109040 188408
rect 18656 188368 18662 188380
rect 109034 188368 109040 188380
rect 109092 188368 109098 188420
rect 152458 188368 152464 188420
rect 152516 188408 152522 188420
rect 349430 188408 349436 188420
rect 152516 188380 349436 188408
rect 152516 188368 152522 188380
rect 349430 188368 349436 188380
rect 349488 188368 349494 188420
rect 80146 188300 80152 188352
rect 80204 188340 80210 188352
rect 327350 188340 327356 188352
rect 80204 188312 327356 188340
rect 80204 188300 80210 188312
rect 327350 188300 327356 188312
rect 327408 188300 327414 188352
rect 106182 187756 106188 187808
rect 106240 187796 106246 187808
rect 167730 187796 167736 187808
rect 106240 187768 167736 187796
rect 106240 187756 106246 187768
rect 167730 187756 167736 187768
rect 167788 187756 167794 187808
rect 100662 187688 100668 187740
rect 100720 187728 100726 187740
rect 170398 187728 170404 187740
rect 100720 187700 170404 187728
rect 100720 187688 100726 187700
rect 170398 187688 170404 187700
rect 170456 187688 170462 187740
rect 157242 187280 157248 187332
rect 157300 187320 157306 187332
rect 189718 187320 189724 187332
rect 157300 187292 189724 187320
rect 157300 187280 157306 187292
rect 189718 187280 189724 187292
rect 189776 187280 189782 187332
rect 148410 187212 148416 187264
rect 148468 187252 148474 187264
rect 252738 187252 252744 187264
rect 148468 187224 252744 187252
rect 148468 187212 148474 187224
rect 252738 187212 252744 187224
rect 252796 187212 252802 187264
rect 129090 187144 129096 187196
rect 129148 187184 129154 187196
rect 256694 187184 256700 187196
rect 129148 187156 256700 187184
rect 129148 187144 129154 187156
rect 256694 187144 256700 187156
rect 256752 187144 256758 187196
rect 63402 187076 63408 187128
rect 63460 187116 63466 187128
rect 249058 187116 249064 187128
rect 63460 187088 249064 187116
rect 63460 187076 63466 187088
rect 249058 187076 249064 187088
rect 249116 187076 249122 187128
rect 95326 187008 95332 187060
rect 95384 187048 95390 187060
rect 321278 187048 321284 187060
rect 95384 187020 321284 187048
rect 95384 187008 95390 187020
rect 321278 187008 321284 187020
rect 321336 187008 321342 187060
rect 73246 186940 73252 186992
rect 73304 186980 73310 186992
rect 320174 186980 320180 186992
rect 73304 186952 320180 186980
rect 73304 186940 73310 186952
rect 320174 186940 320180 186952
rect 320232 186940 320238 186992
rect 155310 185852 155316 185904
rect 155368 185892 155374 185904
rect 255590 185892 255596 185904
rect 155368 185864 255596 185892
rect 155368 185852 155374 185864
rect 255590 185852 255596 185864
rect 255648 185852 255654 185904
rect 107654 185784 107660 185836
rect 107712 185824 107718 185836
rect 346578 185824 346584 185836
rect 107712 185796 346584 185824
rect 107712 185784 107718 185796
rect 346578 185784 346584 185796
rect 346636 185784 346642 185836
rect 68922 185716 68928 185768
rect 68980 185756 68986 185768
rect 321738 185756 321744 185768
rect 68980 185728 321744 185756
rect 68980 185716 68986 185728
rect 321738 185716 321744 185728
rect 321796 185716 321802 185768
rect 69014 185648 69020 185700
rect 69072 185688 69078 185700
rect 323118 185688 323124 185700
rect 69072 185660 323124 185688
rect 69072 185648 69078 185660
rect 323118 185648 323124 185660
rect 323176 185648 323182 185700
rect 59262 185580 59268 185632
rect 59320 185620 59326 185632
rect 337010 185620 337016 185632
rect 59320 185592 337016 185620
rect 59320 185580 59326 185592
rect 337010 185580 337016 185592
rect 337068 185580 337074 185632
rect 134518 184900 134524 184952
rect 134576 184940 134582 184952
rect 210602 184940 210608 184952
rect 134576 184912 210608 184940
rect 134576 184900 134582 184912
rect 210602 184900 210608 184912
rect 210660 184900 210666 184952
rect 222838 184424 222844 184476
rect 222896 184464 222902 184476
rect 350626 184464 350632 184476
rect 222896 184436 350632 184464
rect 222896 184424 222902 184436
rect 350626 184424 350632 184436
rect 350684 184424 350690 184476
rect 163498 184356 163504 184408
rect 163556 184396 163562 184408
rect 334250 184396 334256 184408
rect 163556 184368 334256 184396
rect 163556 184356 163562 184368
rect 334250 184356 334256 184368
rect 334308 184356 334314 184408
rect 63310 184288 63316 184340
rect 63368 184328 63374 184340
rect 256786 184328 256792 184340
rect 63368 184300 256792 184328
rect 63368 184288 63374 184300
rect 256786 184288 256792 184300
rect 256844 184288 256850 184340
rect 84194 184220 84200 184272
rect 84252 184260 84258 184272
rect 325970 184260 325976 184272
rect 84252 184232 325976 184260
rect 84252 184220 84258 184232
rect 325970 184220 325976 184232
rect 326028 184220 326034 184272
rect 88334 184152 88340 184204
rect 88392 184192 88398 184204
rect 346670 184192 346676 184204
rect 88392 184164 346676 184192
rect 88392 184152 88398 184164
rect 346670 184152 346676 184164
rect 346728 184152 346734 184204
rect 114462 183608 114468 183660
rect 114520 183648 114526 183660
rect 169294 183648 169300 183660
rect 114520 183620 169300 183648
rect 114520 183608 114526 183620
rect 169294 183608 169300 183620
rect 169352 183608 169358 183660
rect 128262 183540 128268 183592
rect 128320 183580 128326 183592
rect 214742 183580 214748 183592
rect 128320 183552 214748 183580
rect 128320 183540 128326 183552
rect 214742 183540 214748 183552
rect 214800 183540 214806 183592
rect 220078 183132 220084 183184
rect 220136 183172 220142 183184
rect 258350 183172 258356 183184
rect 220136 183144 258356 183172
rect 220136 183132 220142 183144
rect 258350 183132 258356 183144
rect 258408 183132 258414 183184
rect 156690 183064 156696 183116
rect 156748 183104 156754 183116
rect 245654 183104 245660 183116
rect 156748 183076 245660 183104
rect 156748 183064 156754 183076
rect 245654 183064 245660 183076
rect 245712 183064 245718 183116
rect 172422 182996 172428 183048
rect 172480 183036 172486 183048
rect 282178 183036 282184 183048
rect 172480 183008 282184 183036
rect 172480 182996 172486 183008
rect 282178 182996 282184 183008
rect 282236 182996 282242 183048
rect 189902 182928 189908 182980
rect 189960 182968 189966 182980
rect 334066 182968 334072 182980
rect 189960 182940 334072 182968
rect 189960 182928 189966 182940
rect 334066 182928 334072 182940
rect 334124 182928 334130 182980
rect 148502 182860 148508 182912
rect 148560 182900 148566 182912
rect 338298 182900 338304 182912
rect 148560 182872 338304 182900
rect 148560 182860 148566 182872
rect 338298 182860 338304 182872
rect 338356 182860 338362 182912
rect 93854 182792 93860 182844
rect 93912 182832 93918 182844
rect 330110 182832 330116 182844
rect 93912 182804 330116 182832
rect 93912 182792 93918 182804
rect 330110 182792 330116 182804
rect 330168 182792 330174 182844
rect 127802 182180 127808 182232
rect 127860 182220 127866 182232
rect 206462 182220 206468 182232
rect 127860 182192 206468 182220
rect 127860 182180 127866 182192
rect 206462 182180 206468 182192
rect 206520 182180 206526 182232
rect 228358 181704 228364 181756
rect 228416 181744 228422 181756
rect 265066 181744 265072 181756
rect 228416 181716 265072 181744
rect 228416 181704 228422 181716
rect 265066 181704 265072 181716
rect 265124 181704 265130 181756
rect 140038 181636 140044 181688
rect 140096 181676 140102 181688
rect 249334 181676 249340 181688
rect 140096 181648 249340 181676
rect 140096 181636 140102 181648
rect 249334 181636 249340 181648
rect 249392 181636 249398 181688
rect 224218 181568 224224 181620
rect 224276 181608 224282 181620
rect 332778 181608 332784 181620
rect 224276 181580 332784 181608
rect 224276 181568 224282 181580
rect 332778 181568 332784 181580
rect 332836 181568 332842 181620
rect 156598 181500 156604 181552
rect 156656 181540 156662 181552
rect 341150 181540 341156 181552
rect 156656 181512 341156 181540
rect 156656 181500 156662 181512
rect 341150 181500 341156 181512
rect 341208 181500 341214 181552
rect 147030 181432 147036 181484
rect 147088 181472 147094 181484
rect 342530 181472 342536 181484
rect 147088 181444 342536 181472
rect 147088 181432 147094 181444
rect 342530 181432 342536 181444
rect 342588 181432 342594 181484
rect 116946 180956 116952 181008
rect 117004 180996 117010 181008
rect 166534 180996 166540 181008
rect 117004 180968 166540 180996
rect 117004 180956 117010 180968
rect 166534 180956 166540 180968
rect 166592 180956 166598 181008
rect 112990 180888 112996 180940
rect 113048 180928 113054 180940
rect 167822 180928 167828 180940
rect 113048 180900 167828 180928
rect 113048 180888 113054 180900
rect 167822 180888 167828 180900
rect 167880 180888 167886 180940
rect 129458 180820 129464 180872
rect 129516 180860 129522 180872
rect 206554 180860 206560 180872
rect 129516 180832 206560 180860
rect 129516 180820 129522 180832
rect 206554 180820 206560 180832
rect 206612 180820 206618 180872
rect 162762 180276 162768 180328
rect 162820 180316 162826 180328
rect 203518 180316 203524 180328
rect 162820 180288 203524 180316
rect 162820 180276 162826 180288
rect 203518 180276 203524 180288
rect 203576 180276 203582 180328
rect 231118 180276 231124 180328
rect 231176 180316 231182 180328
rect 262490 180316 262496 180328
rect 231176 180288 262496 180316
rect 231176 180276 231182 180288
rect 262490 180276 262496 180288
rect 262548 180276 262554 180328
rect 169110 180208 169116 180260
rect 169168 180248 169174 180260
rect 318334 180248 318340 180260
rect 169168 180220 318340 180248
rect 169168 180208 169174 180220
rect 318334 180208 318340 180220
rect 318392 180208 318398 180260
rect 64782 180140 64788 180192
rect 64840 180180 64846 180192
rect 251266 180180 251272 180192
rect 64840 180152 251272 180180
rect 64840 180140 64846 180152
rect 251266 180140 251272 180152
rect 251324 180140 251330 180192
rect 283558 180140 283564 180192
rect 283616 180180 283622 180192
rect 335446 180180 335452 180192
rect 283616 180152 335452 180180
rect 283616 180140 283622 180152
rect 335446 180140 335452 180152
rect 335504 180140 335510 180192
rect 157978 180072 157984 180124
rect 158036 180112 158042 180124
rect 345198 180112 345204 180124
rect 158036 180084 345204 180112
rect 158036 180072 158042 180084
rect 345198 180072 345204 180084
rect 345256 180072 345262 180124
rect 113910 179528 113916 179580
rect 113968 179568 113974 179580
rect 166350 179568 166356 179580
rect 113968 179540 166356 179568
rect 113968 179528 113974 179540
rect 166350 179528 166356 179540
rect 166408 179528 166414 179580
rect 110690 179460 110696 179512
rect 110748 179500 110754 179512
rect 166258 179500 166264 179512
rect 110748 179472 166264 179500
rect 110748 179460 110754 179472
rect 166258 179460 166264 179472
rect 166316 179460 166322 179512
rect 97810 179392 97816 179444
rect 97868 179432 97874 179444
rect 169202 179432 169208 179444
rect 97868 179404 169208 179432
rect 97868 179392 97874 179404
rect 169202 179392 169208 179404
rect 169260 179392 169266 179444
rect 373258 179324 373264 179376
rect 373316 179364 373322 179376
rect 580166 179364 580172 179376
rect 373316 179336 580172 179364
rect 373316 179324 373322 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 246390 178984 246396 179036
rect 246448 179024 246454 179036
rect 252554 179024 252560 179036
rect 246448 178996 252560 179024
rect 246448 178984 246454 178996
rect 252554 178984 252560 178996
rect 252612 178984 252618 179036
rect 240778 178916 240784 178968
rect 240836 178956 240842 178968
rect 256878 178956 256884 178968
rect 240836 178928 256884 178956
rect 240836 178916 240842 178928
rect 256878 178916 256884 178928
rect 256936 178916 256942 178968
rect 210418 178848 210424 178900
rect 210476 178888 210482 178900
rect 249978 178888 249984 178900
rect 210476 178860 249984 178888
rect 210476 178848 210482 178860
rect 249978 178848 249984 178860
rect 250036 178848 250042 178900
rect 312538 178848 312544 178900
rect 312596 178888 312602 178900
rect 339586 178888 339592 178900
rect 312596 178860 339592 178888
rect 312596 178848 312602 178860
rect 339586 178848 339592 178860
rect 339644 178848 339650 178900
rect 167638 178780 167644 178832
rect 167696 178820 167702 178832
rect 251450 178820 251456 178832
rect 167696 178792 251456 178820
rect 167696 178780 167702 178792
rect 251450 178780 251456 178792
rect 251508 178780 251514 178832
rect 305638 178780 305644 178832
rect 305696 178820 305702 178832
rect 335538 178820 335544 178832
rect 305696 178792 335544 178820
rect 305696 178780 305702 178792
rect 335538 178780 335544 178792
rect 335596 178780 335602 178832
rect 128998 178712 129004 178764
rect 129056 178752 129062 178764
rect 318702 178752 318708 178764
rect 129056 178724 318708 178752
rect 129056 178712 129062 178724
rect 318702 178712 318708 178724
rect 318760 178712 318766 178764
rect 78674 178644 78680 178696
rect 78732 178684 78738 178696
rect 343910 178684 343916 178696
rect 78732 178656 343916 178684
rect 78732 178644 78738 178656
rect 343910 178644 343916 178656
rect 343968 178644 343974 178696
rect 109862 178236 109868 178288
rect 109920 178276 109926 178288
rect 162762 178276 162768 178288
rect 109920 178248 162768 178276
rect 109920 178236 109926 178248
rect 162762 178236 162768 178248
rect 162820 178236 162826 178288
rect 148226 178168 148232 178220
rect 148284 178208 148290 178220
rect 206278 178208 206284 178220
rect 148284 178180 206284 178208
rect 148284 178168 148290 178180
rect 206278 178168 206284 178180
rect 206336 178168 206342 178220
rect 122006 178100 122012 178152
rect 122064 178140 122070 178152
rect 196710 178140 196716 178152
rect 122064 178112 196716 178140
rect 122064 178100 122070 178112
rect 196710 178100 196716 178112
rect 196768 178100 196774 178152
rect 124950 178032 124956 178084
rect 125008 178072 125014 178084
rect 214926 178072 214932 178084
rect 125008 178044 214932 178072
rect 125008 178032 125014 178044
rect 214926 178032 214932 178044
rect 214984 178032 214990 178084
rect 119706 177964 119712 178016
rect 119764 178004 119770 178016
rect 134518 178004 134524 178016
rect 119764 177976 134524 178004
rect 119764 177964 119770 177976
rect 134518 177964 134524 177976
rect 134576 177964 134582 178016
rect 217962 177964 217968 178016
rect 218020 178004 218026 178016
rect 220814 178004 220820 178016
rect 218020 177976 220820 178004
rect 218020 177964 218026 177976
rect 220814 177964 220820 177976
rect 220872 177964 220878 178016
rect 236638 177624 236644 177676
rect 236696 177664 236702 177676
rect 249242 177664 249248 177676
rect 236696 177636 249248 177664
rect 236696 177624 236702 177636
rect 249242 177624 249248 177636
rect 249300 177624 249306 177676
rect 242250 177556 242256 177608
rect 242308 177596 242314 177608
rect 256970 177596 256976 177608
rect 242308 177568 256976 177596
rect 242308 177556 242314 177568
rect 256970 177556 256976 177568
rect 257028 177556 257034 177608
rect 168282 177488 168288 177540
rect 168340 177528 168346 177540
rect 202138 177528 202144 177540
rect 168340 177500 202144 177528
rect 168340 177488 168346 177500
rect 202138 177488 202144 177500
rect 202196 177488 202202 177540
rect 216582 177488 216588 177540
rect 216640 177528 216646 177540
rect 224954 177528 224960 177540
rect 216640 177500 224960 177528
rect 216640 177488 216646 177500
rect 224954 177488 224960 177500
rect 225012 177488 225018 177540
rect 242158 177488 242164 177540
rect 242216 177528 242222 177540
rect 262306 177528 262312 177540
rect 242216 177500 262312 177528
rect 242216 177488 242222 177500
rect 262306 177488 262312 177500
rect 262364 177488 262370 177540
rect 318058 177488 318064 177540
rect 318116 177528 318122 177540
rect 318116 177500 325694 177528
rect 318116 177488 318122 177500
rect 169018 177420 169024 177472
rect 169076 177460 169082 177472
rect 251358 177460 251364 177472
rect 169076 177432 251364 177460
rect 169076 177420 169082 177432
rect 251358 177420 251364 177432
rect 251416 177420 251422 177472
rect 318334 177420 318340 177472
rect 318392 177460 318398 177472
rect 321830 177460 321836 177472
rect 318392 177432 321836 177460
rect 318392 177420 318398 177432
rect 321830 177420 321836 177432
rect 321888 177420 321894 177472
rect 325666 177460 325694 177500
rect 332870 177460 332876 177472
rect 325666 177432 332876 177460
rect 332870 177420 332876 177432
rect 332928 177420 332934 177472
rect 164878 177352 164884 177404
rect 164936 177392 164942 177404
rect 249150 177392 249156 177404
rect 164936 177364 249156 177392
rect 164936 177352 164942 177364
rect 249150 177352 249156 177364
rect 249208 177352 249214 177404
rect 315390 177352 315396 177404
rect 315448 177392 315454 177404
rect 331398 177392 331404 177404
rect 315448 177364 331404 177392
rect 315448 177352 315454 177364
rect 331398 177352 331404 177364
rect 331456 177352 331462 177404
rect 1302 177284 1308 177336
rect 1360 177324 1366 177336
rect 120074 177324 120080 177336
rect 1360 177296 120080 177324
rect 1360 177284 1366 177296
rect 120074 177284 120080 177296
rect 120132 177284 120138 177336
rect 166442 177284 166448 177336
rect 166500 177324 166506 177336
rect 330018 177324 330024 177336
rect 166500 177296 330024 177324
rect 166500 177284 166506 177296
rect 330018 177284 330024 177296
rect 330076 177284 330082 177336
rect 108114 177012 108120 177064
rect 108172 177052 108178 177064
rect 165246 177052 165252 177064
rect 108172 177024 165252 177052
rect 108172 177012 108178 177024
rect 165246 177012 165252 177024
rect 165304 177012 165310 177064
rect 132034 176944 132040 176996
rect 132092 176984 132098 176996
rect 165430 176984 165436 176996
rect 132092 176956 165436 176984
rect 132092 176944 132098 176956
rect 165430 176944 165436 176956
rect 165488 176944 165494 176996
rect 123018 176876 123024 176928
rect 123076 176916 123082 176928
rect 165522 176916 165528 176928
rect 123076 176888 165528 176916
rect 123076 176876 123082 176888
rect 165522 176876 165528 176888
rect 165580 176876 165586 176928
rect 125870 176808 125876 176860
rect 125928 176848 125934 176860
rect 167914 176848 167920 176860
rect 125928 176820 167920 176848
rect 125928 176808 125934 176820
rect 167914 176808 167920 176820
rect 167972 176808 167978 176860
rect 158990 176740 158996 176792
rect 159048 176780 159054 176792
rect 187050 176780 187056 176792
rect 159048 176752 187056 176780
rect 159048 176740 159054 176752
rect 187050 176740 187056 176752
rect 187108 176740 187114 176792
rect 134426 176672 134432 176724
rect 134484 176712 134490 176724
rect 195974 176712 195980 176724
rect 134484 176684 195980 176712
rect 134484 176672 134490 176684
rect 195974 176672 195980 176684
rect 196032 176672 196038 176724
rect 318150 176672 318156 176724
rect 318208 176712 318214 176724
rect 321554 176712 321560 176724
rect 318208 176684 321560 176712
rect 318208 176672 318214 176684
rect 321554 176672 321560 176684
rect 321612 176672 321618 176724
rect 135714 176604 135720 176656
rect 135772 176644 135778 176656
rect 213914 176644 213920 176656
rect 135772 176616 213920 176644
rect 135772 176604 135778 176616
rect 213914 176604 213920 176616
rect 213972 176604 213978 176656
rect 245654 176604 245660 176656
rect 245712 176644 245718 176656
rect 249886 176644 249892 176656
rect 245712 176616 249892 176644
rect 245712 176604 245718 176616
rect 249886 176604 249892 176616
rect 249944 176604 249950 176656
rect 311250 176604 311256 176656
rect 311308 176644 311314 176656
rect 321462 176644 321468 176656
rect 311308 176616 321468 176644
rect 311308 176604 311314 176616
rect 321462 176604 321468 176616
rect 321520 176604 321526 176656
rect 162762 176196 162768 176248
rect 162820 176236 162826 176248
rect 206370 176236 206376 176248
rect 162820 176208 206376 176236
rect 162820 176196 162826 176208
rect 206370 176196 206376 176208
rect 206428 176196 206434 176248
rect 120810 176128 120816 176180
rect 120868 176168 120874 176180
rect 167638 176168 167644 176180
rect 120868 176140 167644 176168
rect 120868 176128 120874 176140
rect 167638 176128 167644 176140
rect 167696 176128 167702 176180
rect 115750 176060 115756 176112
rect 115808 176100 115814 176112
rect 166442 176100 166448 176112
rect 115808 176072 166448 176100
rect 115808 176060 115814 176072
rect 166442 176060 166448 176072
rect 166500 176060 166506 176112
rect 249058 176060 249064 176112
rect 249116 176100 249122 176112
rect 253934 176100 253940 176112
rect 249116 176072 253940 176100
rect 249116 176060 249122 176072
rect 253934 176060 253940 176072
rect 253992 176060 253998 176112
rect 104618 175992 104624 176044
rect 104676 176032 104682 176044
rect 169018 176032 169024 176044
rect 104676 176004 169024 176032
rect 104676 175992 104682 176004
rect 169018 175992 169024 176004
rect 169076 175992 169082 176044
rect 246298 175992 246304 176044
rect 246356 176032 246362 176044
rect 255406 176032 255412 176044
rect 246356 176004 255412 176032
rect 246356 175992 246362 176004
rect 255406 175992 255412 176004
rect 255464 175992 255470 176044
rect 305638 175992 305644 176044
rect 305696 176032 305702 176044
rect 306374 176032 306380 176044
rect 305696 176004 306380 176032
rect 305696 175992 305702 176004
rect 306374 175992 306380 176004
rect 306432 176032 306438 176044
rect 307570 176032 307576 176044
rect 306432 176004 307576 176032
rect 306432 175992 306438 176004
rect 307570 175992 307576 176004
rect 307628 175992 307634 176044
rect 319622 175992 319628 176044
rect 319680 176032 319686 176044
rect 326062 176032 326068 176044
rect 319680 176004 326068 176032
rect 319680 175992 319686 176004
rect 326062 175992 326068 176004
rect 326120 175992 326126 176044
rect 130746 175924 130752 175976
rect 130804 175964 130810 175976
rect 214006 175964 214012 175976
rect 130804 175936 214012 175964
rect 130804 175924 130810 175936
rect 214006 175924 214012 175936
rect 214064 175924 214070 175976
rect 247678 175924 247684 175976
rect 247736 175964 247742 175976
rect 259638 175964 259644 175976
rect 247736 175936 259644 175964
rect 247736 175924 247742 175936
rect 259638 175924 259644 175936
rect 259696 175924 259702 175976
rect 319530 175924 319536 175976
rect 319588 175964 319594 175976
rect 335630 175964 335636 175976
rect 319588 175936 335636 175964
rect 319588 175924 319594 175936
rect 335630 175924 335636 175936
rect 335688 175924 335694 175976
rect 318702 175856 318708 175908
rect 318760 175896 318766 175908
rect 321922 175896 321928 175908
rect 318760 175868 321928 175896
rect 318760 175856 318766 175868
rect 321922 175856 321928 175868
rect 321980 175856 321986 175908
rect 243538 175788 243544 175840
rect 243596 175828 243602 175840
rect 248046 175828 248052 175840
rect 243596 175800 248052 175828
rect 243596 175788 243602 175800
rect 248046 175788 248052 175800
rect 248104 175788 248110 175840
rect 195974 175176 195980 175228
rect 196032 175216 196038 175228
rect 213914 175216 213920 175228
rect 196032 175188 213920 175216
rect 196032 175176 196038 175188
rect 213914 175176 213920 175188
rect 213972 175176 213978 175228
rect 3510 150356 3516 150408
rect 3568 150396 3574 150408
rect 26878 150396 26884 150408
rect 3568 150368 26884 150396
rect 3568 150356 3574 150368
rect 26878 150356 26884 150368
rect 26936 150356 26942 150408
rect 3510 137912 3516 137964
rect 3568 137952 3574 137964
rect 13078 137952 13084 137964
rect 3568 137924 13084 137952
rect 3568 137912 3574 137924
rect 13078 137912 13084 137924
rect 13136 137912 13142 137964
rect 59262 125604 59268 125656
rect 59320 125644 59326 125656
rect 66162 125644 66168 125656
rect 59320 125616 66168 125644
rect 59320 125604 59326 125616
rect 66162 125604 66168 125616
rect 66220 125604 66226 125656
rect 63310 124176 63316 124228
rect 63368 124216 63374 124228
rect 65518 124216 65524 124228
rect 63368 124188 65524 124216
rect 63368 124176 63374 124188
rect 65518 124176 65524 124188
rect 65576 124176 65582 124228
rect 62022 122816 62028 122868
rect 62080 122856 62086 122868
rect 66070 122856 66076 122868
rect 62080 122828 66076 122856
rect 62080 122816 62086 122828
rect 66070 122816 66076 122828
rect 66128 122816 66134 122868
rect 63402 121456 63408 121508
rect 63460 121496 63466 121508
rect 66070 121496 66076 121508
rect 63460 121468 66076 121496
rect 63460 121456 63466 121468
rect 66070 121456 66076 121468
rect 66128 121456 66134 121508
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 21358 111772 21364 111784
rect 3200 111744 21364 111772
rect 3200 111732 3206 111744
rect 21358 111732 21364 111744
rect 21416 111732 21422 111784
rect 2774 97724 2780 97776
rect 2832 97764 2838 97776
rect 4798 97764 4804 97776
rect 2832 97736 4804 97764
rect 2832 97724 2838 97736
rect 4798 97724 4804 97736
rect 4856 97724 4862 97776
rect 165430 174496 165436 174548
rect 165488 174536 165494 174548
rect 213914 174536 213920 174548
rect 165488 174508 213920 174536
rect 165488 174496 165494 174508
rect 213914 174496 213920 174508
rect 213972 174496 213978 174548
rect 288066 174020 288072 174072
rect 288124 174060 288130 174072
rect 307662 174060 307668 174072
rect 288124 174032 307668 174060
rect 288124 174020 288130 174032
rect 307662 174020 307668 174032
rect 307720 174020 307726 174072
rect 282270 173952 282276 174004
rect 282328 173992 282334 174004
rect 306742 173992 306748 174004
rect 282328 173964 306748 173992
rect 282328 173952 282334 173964
rect 306742 173952 306748 173964
rect 306800 173952 306806 174004
rect 264422 173884 264428 173936
rect 264480 173924 264486 173936
rect 307570 173924 307576 173936
rect 264480 173896 307576 173924
rect 264480 173884 264486 173896
rect 307570 173884 307576 173896
rect 307628 173884 307634 173936
rect 324314 173816 324320 173868
rect 324372 173856 324378 173868
rect 326062 173856 326068 173868
rect 324372 173828 326068 173856
rect 324372 173816 324378 173828
rect 326062 173816 326068 173828
rect 326120 173816 326126 173868
rect 252094 173680 252100 173732
rect 252152 173720 252158 173732
rect 256694 173720 256700 173732
rect 252152 173692 256700 173720
rect 252152 173680 252158 173692
rect 256694 173680 256700 173692
rect 256752 173680 256758 173732
rect 165246 173136 165252 173188
rect 165304 173176 165310 173188
rect 214282 173176 214288 173188
rect 165304 173148 214288 173176
rect 165304 173136 165310 173148
rect 214282 173136 214288 173148
rect 214340 173136 214346 173188
rect 271230 172592 271236 172644
rect 271288 172632 271294 172644
rect 307294 172632 307300 172644
rect 271288 172604 307300 172632
rect 271288 172592 271294 172604
rect 307294 172592 307300 172604
rect 307352 172592 307358 172644
rect 269850 172524 269856 172576
rect 269908 172564 269914 172576
rect 306926 172564 306932 172576
rect 269908 172536 306932 172564
rect 269908 172524 269914 172536
rect 306926 172524 306932 172536
rect 306984 172524 306990 172576
rect 206554 172456 206560 172508
rect 206612 172496 206618 172508
rect 213914 172496 213920 172508
rect 206612 172468 213920 172496
rect 206612 172456 206618 172468
rect 213914 172456 213920 172468
rect 213972 172456 213978 172508
rect 252462 171504 252468 171556
rect 252520 171544 252526 171556
rect 258166 171544 258172 171556
rect 252520 171516 258172 171544
rect 252520 171504 252526 171516
rect 258166 171504 258172 171516
rect 258224 171504 258230 171556
rect 280798 171232 280804 171284
rect 280856 171272 280862 171284
rect 306926 171272 306932 171284
rect 280856 171244 306932 171272
rect 280856 171232 280862 171244
rect 306926 171232 306932 171244
rect 306984 171232 306990 171284
rect 265618 171164 265624 171216
rect 265676 171204 265682 171216
rect 307662 171204 307668 171216
rect 265676 171176 307668 171204
rect 265676 171164 265682 171176
rect 307662 171164 307668 171176
rect 307720 171164 307726 171216
rect 168006 171096 168012 171148
rect 168064 171136 168070 171148
rect 210510 171136 210516 171148
rect 168064 171108 210516 171136
rect 168064 171096 168070 171108
rect 210510 171096 210516 171108
rect 210568 171096 210574 171148
rect 261662 171096 261668 171148
rect 261720 171136 261726 171148
rect 307570 171136 307576 171148
rect 261720 171108 307576 171136
rect 261720 171096 261726 171108
rect 307570 171096 307576 171108
rect 307628 171096 307634 171148
rect 167914 171028 167920 171080
rect 167972 171068 167978 171080
rect 214006 171068 214012 171080
rect 167972 171040 214012 171068
rect 167972 171028 167978 171040
rect 214006 171028 214012 171040
rect 214064 171028 214070 171080
rect 206462 170960 206468 171012
rect 206520 171000 206526 171012
rect 213914 171000 213920 171012
rect 206520 170972 213920 171000
rect 206520 170960 206526 170972
rect 213914 170960 213920 170972
rect 213972 170960 213978 171012
rect 251358 170892 251364 170944
rect 251416 170932 251422 170944
rect 251542 170932 251548 170944
rect 251416 170904 251548 170932
rect 251416 170892 251422 170904
rect 251542 170892 251548 170904
rect 251600 170892 251606 170944
rect 251726 170892 251732 170944
rect 251784 170932 251790 170944
rect 255498 170932 255504 170944
rect 251784 170904 255504 170932
rect 251784 170892 251790 170904
rect 255498 170892 255504 170904
rect 255556 170892 255562 170944
rect 294598 170348 294604 170400
rect 294656 170388 294662 170400
rect 306558 170388 306564 170400
rect 294656 170360 306564 170388
rect 294656 170348 294662 170360
rect 306558 170348 306564 170360
rect 306616 170348 306622 170400
rect 251358 170280 251364 170332
rect 251416 170320 251422 170332
rect 253934 170320 253940 170332
rect 251416 170292 253940 170320
rect 251416 170280 251422 170292
rect 253934 170280 253940 170292
rect 253992 170280 253998 170332
rect 251818 169804 251824 169856
rect 251876 169844 251882 169856
rect 259546 169844 259552 169856
rect 251876 169816 259552 169844
rect 251876 169804 251882 169816
rect 259546 169804 259552 169816
rect 259604 169804 259610 169856
rect 267090 169804 267096 169856
rect 267148 169844 267154 169856
rect 307662 169844 307668 169856
rect 267148 169816 307668 169844
rect 267148 169804 267154 169816
rect 307662 169804 307668 169816
rect 307720 169804 307726 169856
rect 260374 169736 260380 169788
rect 260432 169776 260438 169788
rect 306742 169776 306748 169788
rect 260432 169748 306748 169776
rect 260432 169736 260438 169748
rect 306742 169736 306748 169748
rect 306800 169736 306806 169788
rect 252278 169668 252284 169720
rect 252336 169708 252342 169720
rect 262398 169708 262404 169720
rect 252336 169680 262404 169708
rect 252336 169668 252342 169680
rect 262398 169668 262404 169680
rect 262456 169668 262462 169720
rect 324314 169668 324320 169720
rect 324372 169708 324378 169720
rect 337010 169708 337016 169720
rect 324372 169680 337016 169708
rect 324372 169668 324378 169680
rect 337010 169668 337016 169680
rect 337068 169668 337074 169720
rect 169110 168988 169116 169040
rect 169168 169028 169174 169040
rect 214650 169028 214656 169040
rect 169168 169000 214656 169028
rect 169168 168988 169174 169000
rect 214650 168988 214656 169000
rect 214708 168988 214714 169040
rect 283558 168512 283564 168564
rect 283616 168552 283622 168564
rect 307662 168552 307668 168564
rect 283616 168524 307668 168552
rect 283616 168512 283622 168524
rect 307662 168512 307668 168524
rect 307720 168512 307726 168564
rect 273898 168444 273904 168496
rect 273956 168484 273962 168496
rect 307478 168484 307484 168496
rect 273956 168456 307484 168484
rect 273956 168444 273962 168456
rect 307478 168444 307484 168456
rect 307536 168444 307542 168496
rect 262858 168376 262864 168428
rect 262916 168416 262922 168428
rect 307570 168416 307576 168428
rect 262916 168388 307576 168416
rect 262916 168376 262922 168388
rect 307570 168376 307576 168388
rect 307628 168376 307634 168428
rect 167638 168308 167644 168360
rect 167696 168348 167702 168360
rect 214006 168348 214012 168360
rect 167696 168320 214012 168348
rect 167696 168308 167702 168320
rect 214006 168308 214012 168320
rect 214064 168308 214070 168360
rect 251910 168308 251916 168360
rect 251968 168348 251974 168360
rect 255590 168348 255596 168360
rect 251968 168320 255596 168348
rect 251968 168308 251974 168320
rect 255590 168308 255596 168320
rect 255648 168308 255654 168360
rect 324314 168308 324320 168360
rect 324372 168348 324378 168360
rect 334158 168348 334164 168360
rect 324372 168320 334164 168348
rect 324372 168308 324378 168320
rect 334158 168308 334164 168320
rect 334216 168308 334222 168360
rect 196710 168240 196716 168292
rect 196768 168280 196774 168292
rect 213914 168280 213920 168292
rect 196768 168252 213920 168280
rect 196768 168240 196774 168252
rect 213914 168240 213920 168252
rect 213972 168240 213978 168292
rect 252462 167220 252468 167272
rect 252520 167260 252526 167272
rect 258258 167260 258264 167272
rect 252520 167232 258264 167260
rect 252520 167220 252526 167232
rect 258258 167220 258264 167232
rect 258316 167220 258322 167272
rect 291930 167152 291936 167204
rect 291988 167192 291994 167204
rect 307294 167192 307300 167204
rect 291988 167164 307300 167192
rect 291988 167152 291994 167164
rect 307294 167152 307300 167164
rect 307352 167152 307358 167204
rect 278222 167084 278228 167136
rect 278280 167124 278286 167136
rect 307662 167124 307668 167136
rect 278280 167096 307668 167124
rect 278280 167084 278286 167096
rect 307662 167084 307668 167096
rect 307720 167084 307726 167136
rect 275278 167016 275284 167068
rect 275336 167056 275342 167068
rect 307478 167056 307484 167068
rect 275336 167028 307484 167056
rect 275336 167016 275342 167028
rect 307478 167016 307484 167028
rect 307536 167016 307542 167068
rect 166534 166948 166540 167000
rect 166592 166988 166598 167000
rect 214006 166988 214012 167000
rect 166592 166960 214012 166988
rect 166592 166948 166598 166960
rect 214006 166948 214012 166960
rect 214064 166948 214070 167000
rect 252094 166948 252100 167000
rect 252152 166988 252158 167000
rect 261018 166988 261024 167000
rect 252152 166960 261024 166988
rect 252152 166948 252158 166960
rect 261018 166948 261024 166960
rect 261076 166948 261082 167000
rect 189810 166880 189816 166932
rect 189868 166920 189874 166932
rect 213914 166920 213920 166932
rect 189868 166892 213920 166920
rect 189868 166880 189874 166892
rect 213914 166880 213920 166892
rect 213972 166880 213978 166932
rect 210602 166812 210608 166864
rect 210660 166852 210666 166864
rect 214098 166852 214104 166864
rect 210660 166824 214104 166852
rect 210660 166812 210666 166824
rect 214098 166812 214104 166824
rect 214156 166812 214162 166864
rect 252370 166744 252376 166796
rect 252428 166784 252434 166796
rect 256878 166784 256884 166796
rect 252428 166756 256884 166784
rect 252428 166744 252434 166756
rect 256878 166744 256884 166756
rect 256936 166744 256942 166796
rect 252462 166472 252468 166524
rect 252520 166512 252526 166524
rect 258350 166512 258356 166524
rect 252520 166484 258356 166512
rect 252520 166472 252526 166484
rect 258350 166472 258356 166484
rect 258408 166472 258414 166524
rect 269942 165656 269948 165708
rect 270000 165696 270006 165708
rect 307570 165696 307576 165708
rect 270000 165668 307576 165696
rect 270000 165656 270006 165668
rect 307570 165656 307576 165668
rect 307628 165656 307634 165708
rect 259086 165588 259092 165640
rect 259144 165628 259150 165640
rect 307662 165628 307668 165640
rect 259144 165600 307668 165628
rect 259144 165588 259150 165600
rect 307662 165588 307668 165600
rect 307720 165588 307726 165640
rect 166442 165520 166448 165572
rect 166500 165560 166506 165572
rect 213914 165560 213920 165572
rect 166500 165532 213920 165560
rect 166500 165520 166506 165532
rect 213914 165520 213920 165532
rect 213972 165520 213978 165572
rect 252462 165520 252468 165572
rect 252520 165560 252526 165572
rect 266538 165560 266544 165572
rect 252520 165532 266544 165560
rect 252520 165520 252526 165532
rect 266538 165520 266544 165532
rect 266596 165520 266602 165572
rect 324314 165520 324320 165572
rect 324372 165560 324378 165572
rect 335630 165560 335636 165572
rect 324372 165532 335636 165560
rect 324372 165520 324378 165532
rect 335630 165520 335636 165532
rect 335688 165520 335694 165572
rect 169294 165452 169300 165504
rect 169352 165492 169358 165504
rect 214006 165492 214012 165504
rect 169352 165464 214012 165492
rect 169352 165452 169358 165464
rect 214006 165452 214012 165464
rect 214064 165452 214070 165504
rect 252094 165452 252100 165504
rect 252152 165492 252158 165504
rect 263594 165492 263600 165504
rect 252152 165464 263600 165492
rect 252152 165452 252158 165464
rect 263594 165452 263600 165464
rect 263652 165452 263658 165504
rect 251726 165384 251732 165436
rect 251784 165424 251790 165436
rect 262490 165424 262496 165436
rect 251784 165396 262496 165424
rect 251784 165384 251790 165396
rect 262490 165384 262496 165396
rect 262548 165384 262554 165436
rect 271322 164908 271328 164960
rect 271380 164948 271386 164960
rect 306926 164948 306932 164960
rect 271380 164920 306932 164948
rect 271380 164908 271386 164920
rect 306926 164908 306932 164920
rect 306984 164908 306990 164960
rect 257430 164840 257436 164892
rect 257488 164880 257494 164892
rect 307478 164880 307484 164892
rect 257488 164852 307484 164880
rect 257488 164840 257494 164852
rect 307478 164840 307484 164852
rect 307536 164840 307542 164892
rect 300118 164296 300124 164348
rect 300176 164336 300182 164348
rect 307662 164336 307668 164348
rect 300176 164308 307668 164336
rect 300176 164296 300182 164308
rect 307662 164296 307668 164308
rect 307720 164296 307726 164348
rect 287790 164228 287796 164280
rect 287848 164268 287854 164280
rect 307294 164268 307300 164280
rect 287848 164240 307300 164268
rect 287848 164228 287854 164240
rect 307294 164228 307300 164240
rect 307352 164228 307358 164280
rect 166350 164160 166356 164212
rect 166408 164200 166414 164212
rect 213914 164200 213920 164212
rect 166408 164172 213920 164200
rect 166408 164160 166414 164172
rect 213914 164160 213920 164172
rect 213972 164160 213978 164212
rect 252186 164160 252192 164212
rect 252244 164200 252250 164212
rect 270494 164200 270500 164212
rect 252244 164172 270500 164200
rect 252244 164160 252250 164172
rect 270494 164160 270500 164172
rect 270552 164160 270558 164212
rect 324406 164160 324412 164212
rect 324464 164200 324470 164212
rect 331398 164200 331404 164212
rect 324464 164172 331404 164200
rect 324464 164160 324470 164172
rect 331398 164160 331404 164172
rect 331456 164160 331462 164212
rect 167822 164092 167828 164144
rect 167880 164132 167886 164144
rect 214006 164132 214012 164144
rect 167880 164104 214012 164132
rect 167880 164092 167886 164104
rect 214006 164092 214012 164104
rect 214064 164092 214070 164144
rect 324314 164092 324320 164144
rect 324372 164132 324378 164144
rect 329926 164132 329932 164144
rect 324372 164104 329932 164132
rect 324372 164092 324378 164104
rect 329926 164092 329932 164104
rect 329984 164092 329990 164144
rect 290458 163004 290464 163056
rect 290516 163044 290522 163056
rect 307294 163044 307300 163056
rect 290516 163016 307300 163044
rect 290516 163004 290522 163016
rect 307294 163004 307300 163016
rect 307352 163004 307358 163056
rect 272518 162936 272524 162988
rect 272576 162976 272582 162988
rect 306742 162976 306748 162988
rect 272576 162948 306748 162976
rect 272576 162936 272582 162948
rect 306742 162936 306748 162948
rect 306800 162936 306806 162988
rect 265710 162868 265716 162920
rect 265768 162908 265774 162920
rect 307662 162908 307668 162920
rect 265768 162880 307668 162908
rect 265768 162868 265774 162880
rect 307662 162868 307668 162880
rect 307720 162868 307726 162920
rect 166258 162800 166264 162852
rect 166316 162840 166322 162852
rect 213914 162840 213920 162852
rect 166316 162812 213920 162840
rect 166316 162800 166322 162812
rect 213914 162800 213920 162812
rect 213972 162800 213978 162852
rect 252462 162800 252468 162852
rect 252520 162840 252526 162852
rect 263686 162840 263692 162852
rect 252520 162812 263692 162840
rect 252520 162800 252526 162812
rect 263686 162800 263692 162812
rect 263744 162800 263750 162852
rect 324406 162800 324412 162852
rect 324464 162840 324470 162852
rect 342530 162840 342536 162852
rect 324464 162812 342536 162840
rect 324464 162800 324470 162812
rect 342530 162800 342536 162812
rect 342588 162800 342594 162852
rect 206370 162732 206376 162784
rect 206428 162772 206434 162784
rect 214006 162772 214012 162784
rect 206428 162744 214012 162772
rect 206428 162732 206434 162744
rect 214006 162732 214012 162744
rect 214064 162732 214070 162784
rect 324314 162732 324320 162784
rect 324372 162772 324378 162784
rect 332870 162772 332876 162784
rect 324372 162744 332876 162772
rect 324372 162732 324378 162744
rect 332870 162732 332876 162744
rect 332928 162732 332934 162784
rect 262950 162120 262956 162172
rect 263008 162160 263014 162172
rect 307110 162160 307116 162172
rect 263008 162132 307116 162160
rect 263008 162120 263014 162132
rect 307110 162120 307116 162132
rect 307168 162120 307174 162172
rect 289262 161508 289268 161560
rect 289320 161548 289326 161560
rect 307478 161548 307484 161560
rect 289320 161520 307484 161548
rect 289320 161508 289326 161520
rect 307478 161508 307484 161520
rect 307536 161508 307542 161560
rect 279602 161440 279608 161492
rect 279660 161480 279666 161492
rect 307662 161480 307668 161492
rect 279660 161452 307668 161480
rect 279660 161440 279666 161452
rect 307662 161440 307668 161452
rect 307720 161440 307726 161492
rect 171870 161372 171876 161424
rect 171928 161412 171934 161424
rect 213914 161412 213920 161424
rect 171928 161384 213920 161412
rect 171928 161372 171934 161384
rect 213914 161372 213920 161384
rect 213972 161372 213978 161424
rect 252462 161372 252468 161424
rect 252520 161412 252526 161424
rect 260926 161412 260932 161424
rect 252520 161384 260932 161412
rect 252520 161372 252526 161384
rect 260926 161372 260932 161384
rect 260984 161372 260990 161424
rect 324314 161372 324320 161424
rect 324372 161412 324378 161424
rect 346486 161412 346492 161424
rect 324372 161384 346492 161412
rect 324372 161372 324378 161384
rect 346486 161372 346492 161384
rect 346544 161372 346550 161424
rect 324406 161304 324412 161356
rect 324464 161344 324470 161356
rect 332778 161344 332784 161356
rect 324464 161316 332784 161344
rect 324464 161304 324470 161316
rect 332778 161304 332784 161316
rect 332836 161304 332842 161356
rect 260098 160760 260104 160812
rect 260156 160800 260162 160812
rect 306466 160800 306472 160812
rect 260156 160772 306472 160800
rect 260156 160760 260162 160772
rect 306466 160760 306472 160772
rect 306524 160760 306530 160812
rect 254854 160692 254860 160744
rect 254912 160732 254918 160744
rect 307202 160732 307208 160744
rect 254912 160704 307208 160732
rect 254912 160692 254918 160704
rect 307202 160692 307208 160704
rect 307260 160692 307266 160744
rect 303062 160148 303068 160200
rect 303120 160188 303126 160200
rect 307662 160188 307668 160200
rect 303120 160160 307668 160188
rect 303120 160148 303126 160160
rect 307662 160148 307668 160160
rect 307720 160148 307726 160200
rect 276842 160080 276848 160132
rect 276900 160120 276906 160132
rect 307570 160120 307576 160132
rect 276900 160092 307576 160120
rect 276900 160080 276906 160092
rect 307570 160080 307576 160092
rect 307628 160080 307634 160132
rect 167730 160012 167736 160064
rect 167788 160052 167794 160064
rect 213914 160052 213920 160064
rect 167788 160024 213920 160052
rect 167788 160012 167794 160024
rect 213914 160012 213920 160024
rect 213972 160012 213978 160064
rect 324314 160012 324320 160064
rect 324372 160052 324378 160064
rect 331306 160052 331312 160064
rect 324372 160024 331312 160052
rect 324372 160012 324378 160024
rect 331306 160012 331312 160024
rect 331364 160012 331370 160064
rect 169018 159944 169024 159996
rect 169076 159984 169082 159996
rect 214006 159984 214012 159996
rect 169076 159956 214012 159984
rect 169076 159944 169082 159956
rect 214006 159944 214012 159956
rect 214064 159944 214070 159996
rect 251082 159332 251088 159384
rect 251140 159372 251146 159384
rect 259638 159372 259644 159384
rect 251140 159344 259644 159372
rect 251140 159332 251146 159344
rect 259638 159332 259644 159344
rect 259696 159332 259702 159384
rect 278314 159332 278320 159384
rect 278372 159372 278378 159384
rect 307386 159372 307392 159384
rect 278372 159344 307392 159372
rect 278372 159332 278378 159344
rect 307386 159332 307392 159344
rect 307444 159332 307450 159384
rect 264330 158788 264336 158840
rect 264388 158828 264394 158840
rect 306926 158828 306932 158840
rect 264388 158800 306932 158828
rect 264388 158788 264394 158800
rect 306926 158788 306932 158800
rect 306984 158788 306990 158840
rect 261754 158720 261760 158772
rect 261812 158760 261818 158772
rect 307662 158760 307668 158772
rect 261812 158732 307668 158760
rect 261812 158720 261818 158732
rect 307662 158720 307668 158732
rect 307720 158720 307726 158772
rect 203610 158652 203616 158704
rect 203668 158692 203674 158704
rect 213914 158692 213920 158704
rect 203668 158664 213920 158692
rect 203668 158652 203674 158664
rect 213914 158652 213920 158664
rect 213972 158652 213978 158704
rect 251910 158652 251916 158704
rect 251968 158692 251974 158704
rect 256786 158692 256792 158704
rect 251968 158664 256792 158692
rect 251968 158652 251974 158664
rect 256786 158652 256792 158664
rect 256844 158652 256850 158704
rect 324406 158652 324412 158704
rect 324464 158692 324470 158704
rect 341150 158692 341156 158704
rect 324464 158664 341156 158692
rect 324464 158652 324470 158664
rect 341150 158652 341156 158664
rect 341208 158652 341214 158704
rect 324314 158584 324320 158636
rect 324372 158624 324378 158636
rect 334250 158624 334256 158636
rect 324372 158596 334256 158624
rect 324372 158584 324378 158596
rect 334250 158584 334256 158596
rect 334308 158584 334314 158636
rect 287974 157496 287980 157548
rect 288032 157536 288038 157548
rect 307662 157536 307668 157548
rect 288032 157508 307668 157536
rect 288032 157496 288038 157508
rect 307662 157496 307668 157508
rect 307720 157496 307726 157548
rect 260190 157428 260196 157480
rect 260248 157468 260254 157480
rect 307478 157468 307484 157480
rect 260248 157440 307484 157468
rect 260248 157428 260254 157440
rect 307478 157428 307484 157440
rect 307536 157428 307542 157480
rect 257338 157360 257344 157412
rect 257396 157400 257402 157412
rect 306926 157400 306932 157412
rect 257396 157372 306932 157400
rect 257396 157360 257402 157372
rect 306926 157360 306932 157372
rect 306984 157360 306990 157412
rect 170398 157292 170404 157344
rect 170456 157332 170462 157344
rect 213914 157332 213920 157344
rect 170456 157304 213920 157332
rect 170456 157292 170462 157304
rect 213914 157292 213920 157304
rect 213972 157292 213978 157344
rect 252462 157292 252468 157344
rect 252520 157332 252526 157344
rect 272058 157332 272064 157344
rect 252520 157304 272064 157332
rect 252520 157292 252526 157304
rect 272058 157292 272064 157304
rect 272116 157292 272122 157344
rect 252370 157224 252376 157276
rect 252428 157264 252434 157276
rect 265066 157264 265072 157276
rect 252428 157236 265072 157264
rect 252428 157224 252434 157236
rect 265066 157224 265072 157236
rect 265124 157224 265130 157276
rect 324314 157224 324320 157276
rect 324372 157264 324378 157276
rect 339770 157264 339776 157276
rect 324372 157236 339776 157264
rect 324372 157224 324378 157236
rect 339770 157224 339776 157236
rect 339828 157224 339834 157276
rect 285122 156068 285128 156120
rect 285180 156108 285186 156120
rect 307478 156108 307484 156120
rect 285180 156080 307484 156108
rect 285180 156068 285186 156080
rect 307478 156068 307484 156080
rect 307536 156068 307542 156120
rect 258718 156000 258724 156052
rect 258776 156040 258782 156052
rect 307570 156040 307576 156052
rect 258776 156012 307576 156040
rect 258776 156000 258782 156012
rect 307570 156000 307576 156012
rect 307628 156000 307634 156052
rect 254670 155932 254676 155984
rect 254728 155972 254734 155984
rect 307662 155972 307668 155984
rect 254728 155944 307668 155972
rect 254728 155932 254734 155944
rect 307662 155932 307668 155944
rect 307720 155932 307726 155984
rect 169202 155864 169208 155916
rect 169260 155904 169266 155916
rect 214006 155904 214012 155916
rect 169260 155876 214012 155904
rect 169260 155864 169266 155876
rect 214006 155864 214012 155876
rect 214064 155864 214070 155916
rect 251910 155864 251916 155916
rect 251968 155904 251974 155916
rect 255314 155904 255320 155916
rect 251968 155876 255320 155904
rect 251968 155864 251974 155876
rect 255314 155864 255320 155876
rect 255372 155864 255378 155916
rect 324314 155864 324320 155916
rect 324372 155904 324378 155916
rect 338390 155904 338396 155916
rect 324372 155876 338396 155904
rect 324372 155864 324378 155876
rect 338390 155864 338396 155876
rect 338448 155864 338454 155916
rect 170490 155796 170496 155848
rect 170548 155836 170554 155848
rect 213914 155836 213920 155848
rect 170548 155808 213920 155836
rect 170548 155796 170554 155808
rect 213914 155796 213920 155808
rect 213972 155796 213978 155848
rect 251174 155796 251180 155848
rect 251232 155836 251238 155848
rect 254026 155836 254032 155848
rect 251232 155808 254032 155836
rect 251232 155796 251238 155808
rect 254026 155796 254032 155808
rect 254084 155796 254090 155848
rect 324406 155796 324412 155848
rect 324464 155836 324470 155848
rect 328546 155836 328552 155848
rect 324464 155808 328552 155836
rect 324464 155796 324470 155808
rect 328546 155796 328552 155808
rect 328604 155796 328610 155848
rect 252462 155728 252468 155780
rect 252520 155768 252526 155780
rect 269114 155768 269120 155780
rect 252520 155740 269120 155768
rect 252520 155728 252526 155740
rect 269114 155728 269120 155740
rect 269172 155728 269178 155780
rect 295978 154640 295984 154692
rect 296036 154680 296042 154692
rect 307662 154680 307668 154692
rect 296036 154652 307668 154680
rect 296036 154640 296042 154652
rect 307662 154640 307668 154652
rect 307720 154640 307726 154692
rect 261478 154572 261484 154624
rect 261536 154612 261542 154624
rect 307478 154612 307484 154624
rect 261536 154584 307484 154612
rect 261536 154572 261542 154584
rect 307478 154572 307484 154584
rect 307536 154572 307542 154624
rect 251634 154504 251640 154556
rect 251692 154544 251698 154556
rect 270586 154544 270592 154556
rect 251692 154516 270592 154544
rect 251692 154504 251698 154516
rect 270586 154504 270592 154516
rect 270644 154504 270650 154556
rect 324314 154504 324320 154556
rect 324372 154544 324378 154556
rect 346670 154544 346676 154556
rect 324372 154516 346676 154544
rect 324372 154504 324378 154516
rect 346670 154504 346676 154516
rect 346728 154504 346734 154556
rect 283742 153348 283748 153400
rect 283800 153388 283806 153400
rect 307570 153388 307576 153400
rect 283800 153360 307576 153388
rect 283800 153348 283806 153360
rect 307570 153348 307576 153360
rect 307628 153348 307634 153400
rect 184198 153280 184204 153332
rect 184256 153320 184262 153332
rect 214006 153320 214012 153332
rect 184256 153292 214012 153320
rect 184256 153280 184262 153292
rect 214006 153280 214012 153292
rect 214064 153280 214070 153332
rect 263042 153280 263048 153332
rect 263100 153320 263106 153332
rect 307662 153320 307668 153332
rect 263100 153292 307668 153320
rect 263100 153280 263106 153292
rect 307662 153280 307668 153292
rect 307720 153280 307726 153332
rect 324314 153280 324320 153332
rect 324372 153320 324378 153332
rect 327350 153320 327356 153332
rect 324372 153292 327356 153320
rect 324372 153280 324378 153292
rect 327350 153280 327356 153292
rect 327408 153280 327414 153332
rect 171870 153212 171876 153264
rect 171928 153252 171934 153264
rect 213914 153252 213920 153264
rect 171928 153224 213920 153252
rect 171928 153212 171934 153224
rect 213914 153212 213920 153224
rect 213972 153212 213978 153264
rect 255958 153212 255964 153264
rect 256016 153252 256022 153264
rect 307478 153252 307484 153264
rect 256016 153224 307484 153252
rect 256016 153212 256022 153224
rect 307478 153212 307484 153224
rect 307536 153212 307542 153264
rect 251910 153144 251916 153196
rect 251968 153184 251974 153196
rect 281626 153184 281632 153196
rect 251968 153156 281632 153184
rect 251968 153144 251974 153156
rect 281626 153144 281632 153156
rect 281684 153144 281690 153196
rect 252370 153076 252376 153128
rect 252428 153116 252434 153128
rect 271966 153116 271972 153128
rect 252428 153088 271972 153116
rect 252428 153076 252434 153088
rect 271966 153076 271972 153088
rect 272024 153076 272030 153128
rect 252462 153008 252468 153060
rect 252520 153048 252526 153060
rect 269206 153048 269212 153060
rect 252520 153020 269212 153048
rect 252520 153008 252526 153020
rect 269206 153008 269212 153020
rect 269264 153008 269270 153060
rect 258902 152464 258908 152516
rect 258960 152504 258966 152516
rect 306558 152504 306564 152516
rect 258960 152476 306564 152504
rect 258960 152464 258966 152476
rect 306558 152464 306564 152476
rect 306616 152464 306622 152516
rect 203610 151852 203616 151904
rect 203668 151892 203674 151904
rect 213914 151892 213920 151904
rect 203668 151864 213920 151892
rect 203668 151852 203674 151864
rect 213914 151852 213920 151864
rect 213972 151852 213978 151904
rect 300762 151852 300768 151904
rect 300820 151892 300826 151904
rect 307570 151892 307576 151904
rect 300820 151864 307576 151892
rect 300820 151852 300826 151864
rect 307570 151852 307576 151864
rect 307628 151852 307634 151904
rect 191098 151784 191104 151836
rect 191156 151824 191162 151836
rect 214006 151824 214012 151836
rect 191156 151796 214012 151824
rect 191156 151784 191162 151796
rect 214006 151784 214012 151796
rect 214064 151784 214070 151836
rect 253474 151784 253480 151836
rect 253532 151824 253538 151836
rect 307662 151824 307668 151836
rect 253532 151796 307668 151824
rect 253532 151784 253538 151796
rect 307662 151784 307668 151796
rect 307720 151784 307726 151836
rect 251910 151716 251916 151768
rect 251968 151756 251974 151768
rect 276014 151756 276020 151768
rect 251968 151728 276020 151756
rect 251968 151716 251974 151728
rect 276014 151716 276020 151728
rect 276072 151716 276078 151768
rect 324314 151716 324320 151768
rect 324372 151756 324378 151768
rect 346578 151756 346584 151768
rect 324372 151728 346584 151756
rect 324372 151716 324378 151728
rect 346578 151716 346584 151728
rect 346636 151716 346642 151768
rect 252370 151648 252376 151700
rect 252428 151688 252434 151700
rect 274818 151688 274824 151700
rect 252428 151660 274824 151688
rect 252428 151648 252434 151660
rect 274818 151648 274824 151660
rect 274876 151648 274882 151700
rect 252462 151580 252468 151632
rect 252520 151620 252526 151632
rect 267734 151620 267740 151632
rect 252520 151592 267740 151620
rect 252520 151580 252526 151592
rect 267734 151580 267740 151592
rect 267792 151580 267798 151632
rect 177666 151036 177672 151088
rect 177724 151076 177730 151088
rect 210418 151076 210424 151088
rect 177724 151048 210424 151076
rect 177724 151036 177730 151048
rect 210418 151036 210424 151048
rect 210476 151036 210482 151088
rect 298922 150560 298928 150612
rect 298980 150600 298986 150612
rect 307662 150600 307668 150612
rect 298980 150572 307668 150600
rect 298980 150560 298986 150572
rect 307662 150560 307668 150572
rect 307720 150560 307726 150612
rect 211798 150492 211804 150544
rect 211856 150532 211862 150544
rect 214006 150532 214012 150544
rect 211856 150504 214012 150532
rect 211856 150492 211862 150504
rect 214006 150492 214012 150504
rect 214064 150492 214070 150544
rect 268562 150492 268568 150544
rect 268620 150532 268626 150544
rect 307478 150532 307484 150544
rect 268620 150504 307484 150532
rect 268620 150492 268626 150504
rect 307478 150492 307484 150504
rect 307536 150492 307542 150544
rect 207658 150424 207664 150476
rect 207716 150464 207722 150476
rect 213914 150464 213920 150476
rect 207716 150436 213920 150464
rect 207716 150424 207722 150436
rect 213914 150424 213920 150436
rect 213972 150424 213978 150476
rect 254578 150424 254584 150476
rect 254636 150464 254642 150476
rect 306742 150464 306748 150476
rect 254636 150436 306748 150464
rect 254636 150424 254642 150436
rect 306742 150424 306748 150436
rect 306800 150424 306806 150476
rect 206278 150356 206284 150408
rect 206336 150396 206342 150408
rect 214006 150396 214012 150408
rect 206336 150368 214012 150396
rect 206336 150356 206342 150368
rect 214006 150356 214012 150368
rect 214064 150356 214070 150408
rect 251174 150356 251180 150408
rect 251232 150396 251238 150408
rect 254118 150396 254124 150408
rect 251232 150368 254124 150396
rect 251232 150356 251238 150368
rect 254118 150356 254124 150368
rect 254176 150356 254182 150408
rect 324314 150356 324320 150408
rect 324372 150396 324378 150408
rect 330018 150396 330024 150408
rect 324372 150368 330024 150396
rect 324372 150356 324378 150368
rect 330018 150356 330024 150368
rect 330076 150356 330082 150408
rect 210510 150288 210516 150340
rect 210568 150328 210574 150340
rect 213914 150328 213920 150340
rect 210568 150300 213920 150328
rect 210568 150288 210574 150300
rect 213914 150288 213920 150300
rect 213972 150288 213978 150340
rect 252002 150288 252008 150340
rect 252060 150328 252066 150340
rect 273346 150328 273352 150340
rect 252060 150300 273352 150328
rect 252060 150288 252066 150300
rect 273346 150288 273352 150300
rect 273404 150288 273410 150340
rect 252462 150220 252468 150272
rect 252520 150260 252526 150272
rect 274726 150260 274732 150272
rect 252520 150232 274732 150260
rect 252520 150220 252526 150232
rect 274726 150220 274732 150232
rect 274784 150220 274790 150272
rect 296070 149676 296076 149728
rect 296128 149716 296134 149728
rect 307110 149716 307116 149728
rect 296128 149688 307116 149716
rect 296128 149676 296134 149688
rect 307110 149676 307116 149688
rect 307168 149676 307174 149728
rect 300302 149200 300308 149252
rect 300360 149240 300366 149252
rect 306742 149240 306748 149252
rect 300360 149212 306748 149240
rect 300360 149200 300366 149212
rect 306742 149200 306748 149212
rect 306800 149200 306806 149252
rect 301774 149132 301780 149184
rect 301832 149172 301838 149184
rect 307662 149172 307668 149184
rect 301832 149144 307668 149172
rect 301832 149132 301838 149144
rect 307662 149132 307668 149144
rect 307720 149132 307726 149184
rect 253198 149064 253204 149116
rect 253256 149104 253262 149116
rect 307570 149104 307576 149116
rect 253256 149076 307576 149104
rect 253256 149064 253262 149076
rect 307570 149064 307576 149076
rect 307628 149064 307634 149116
rect 187050 148996 187056 149048
rect 187108 149036 187114 149048
rect 213914 149036 213920 149048
rect 187108 149008 213920 149036
rect 187108 148996 187114 149008
rect 213914 148996 213920 149008
rect 213972 148996 213978 149048
rect 252462 148996 252468 149048
rect 252520 149036 252526 149048
rect 266446 149036 266452 149048
rect 252520 149008 266452 149036
rect 252520 148996 252526 149008
rect 266446 148996 266452 149008
rect 266504 148996 266510 149048
rect 324314 148928 324320 148980
rect 324372 148968 324378 148980
rect 349430 148968 349436 148980
rect 324372 148940 349436 148968
rect 324372 148928 324378 148940
rect 349430 148928 349436 148940
rect 349488 148928 349494 148980
rect 251910 148860 251916 148912
rect 251968 148900 251974 148912
rect 255406 148900 255412 148912
rect 251968 148872 255412 148900
rect 251968 148860 251974 148872
rect 255406 148860 255412 148872
rect 255464 148860 255470 148912
rect 324406 148792 324412 148844
rect 324464 148832 324470 148844
rect 325970 148832 325976 148844
rect 324464 148804 325976 148832
rect 324464 148792 324470 148804
rect 325970 148792 325976 148804
rect 326028 148792 326034 148844
rect 252278 148588 252284 148640
rect 252336 148628 252342 148640
rect 259454 148628 259460 148640
rect 252336 148600 259460 148628
rect 252336 148588 252342 148600
rect 259454 148588 259460 148600
rect 259512 148588 259518 148640
rect 269758 147704 269764 147756
rect 269816 147744 269822 147756
rect 307570 147744 307576 147756
rect 269816 147716 307576 147744
rect 269816 147704 269822 147716
rect 307570 147704 307576 147716
rect 307628 147704 307634 147756
rect 198090 147636 198096 147688
rect 198148 147676 198154 147688
rect 213914 147676 213920 147688
rect 198148 147648 213920 147676
rect 198148 147636 198154 147648
rect 213914 147636 213920 147648
rect 213972 147636 213978 147688
rect 254762 147636 254768 147688
rect 254820 147676 254826 147688
rect 307662 147676 307668 147688
rect 254820 147648 307668 147676
rect 254820 147636 254826 147648
rect 307662 147636 307668 147648
rect 307720 147636 307726 147688
rect 252462 147568 252468 147620
rect 252520 147608 252526 147620
rect 277394 147608 277400 147620
rect 252520 147580 277400 147608
rect 252520 147568 252526 147580
rect 277394 147568 277400 147580
rect 277452 147568 277458 147620
rect 324314 147568 324320 147620
rect 324372 147608 324378 147620
rect 343818 147608 343824 147620
rect 324372 147580 343824 147608
rect 324372 147568 324378 147580
rect 343818 147568 343824 147580
rect 343876 147568 343882 147620
rect 252370 147500 252376 147552
rect 252428 147540 252434 147552
rect 276106 147540 276112 147552
rect 252428 147512 276112 147540
rect 252428 147500 252434 147512
rect 276106 147500 276112 147512
rect 276164 147500 276170 147552
rect 251910 146888 251916 146940
rect 251968 146928 251974 146940
rect 273898 146928 273904 146940
rect 251968 146900 273904 146928
rect 251968 146888 251974 146900
rect 273898 146888 273904 146900
rect 273956 146888 273962 146940
rect 276750 146888 276756 146940
rect 276808 146928 276814 146940
rect 307386 146928 307392 146940
rect 276808 146900 307392 146928
rect 276808 146888 276814 146900
rect 307386 146888 307392 146900
rect 307444 146888 307450 146940
rect 304350 146412 304356 146464
rect 304408 146452 304414 146464
rect 307662 146452 307668 146464
rect 304408 146424 307668 146452
rect 304408 146412 304414 146424
rect 307662 146412 307668 146424
rect 307720 146412 307726 146464
rect 182818 146344 182824 146396
rect 182876 146384 182882 146396
rect 213914 146384 213920 146396
rect 182876 146356 213920 146384
rect 182876 146344 182882 146356
rect 213914 146344 213920 146356
rect 213972 146344 213978 146396
rect 274174 146344 274180 146396
rect 274232 146384 274238 146396
rect 307570 146384 307576 146396
rect 274232 146356 307576 146384
rect 274232 146344 274238 146356
rect 307570 146344 307576 146356
rect 307628 146344 307634 146396
rect 167638 146276 167644 146328
rect 167696 146316 167702 146328
rect 214006 146316 214012 146328
rect 167696 146288 214012 146316
rect 167696 146276 167702 146288
rect 214006 146276 214012 146288
rect 214064 146276 214070 146328
rect 256142 146276 256148 146328
rect 256200 146316 256206 146328
rect 307478 146316 307484 146328
rect 256200 146288 307484 146316
rect 256200 146276 256206 146288
rect 307478 146276 307484 146288
rect 307536 146276 307542 146328
rect 252462 146208 252468 146260
rect 252520 146248 252526 146260
rect 273438 146248 273444 146260
rect 252520 146220 273444 146248
rect 252520 146208 252526 146220
rect 273438 146208 273444 146220
rect 273496 146208 273502 146260
rect 252094 146140 252100 146192
rect 252152 146180 252158 146192
rect 262306 146180 262312 146192
rect 252152 146152 262312 146180
rect 252152 146140 252158 146152
rect 262306 146140 262312 146152
rect 262364 146140 262370 146192
rect 251818 146072 251824 146124
rect 251876 146112 251882 146124
rect 258074 146112 258080 146124
rect 251876 146084 258080 146112
rect 251876 146072 251882 146084
rect 258074 146072 258080 146084
rect 258132 146072 258138 146124
rect 282454 145732 282460 145784
rect 282512 145772 282518 145784
rect 303614 145772 303620 145784
rect 282512 145744 303620 145772
rect 282512 145732 282518 145744
rect 303614 145732 303620 145744
rect 303672 145732 303678 145784
rect 265066 145664 265072 145716
rect 265124 145704 265130 145716
rect 293034 145704 293040 145716
rect 265124 145676 293040 145704
rect 265124 145664 265130 145676
rect 293034 145664 293040 145676
rect 293092 145664 293098 145716
rect 256234 145596 256240 145648
rect 256292 145636 256298 145648
rect 306650 145636 306656 145648
rect 256292 145608 306656 145636
rect 256292 145596 256298 145608
rect 306650 145596 306656 145608
rect 306708 145596 306714 145648
rect 196802 145528 196808 145580
rect 196860 145568 196866 145580
rect 214374 145568 214380 145580
rect 196860 145540 214380 145568
rect 196860 145528 196866 145540
rect 214374 145528 214380 145540
rect 214432 145528 214438 145580
rect 253382 145528 253388 145580
rect 253440 145568 253446 145580
rect 307294 145568 307300 145580
rect 253440 145540 307300 145568
rect 253440 145528 253446 145540
rect 307294 145528 307300 145540
rect 307352 145528 307358 145580
rect 252278 145460 252284 145512
rect 252336 145500 252342 145512
rect 256970 145500 256976 145512
rect 252336 145472 256976 145500
rect 252336 145460 252342 145472
rect 256970 145460 256976 145472
rect 257028 145460 257034 145512
rect 193950 144984 193956 145036
rect 194008 145024 194014 145036
rect 213914 145024 213920 145036
rect 194008 144996 213920 145024
rect 194008 144984 194014 144996
rect 213914 144984 213920 144996
rect 213972 144984 213978 145036
rect 304442 144984 304448 145036
rect 304500 145024 304506 145036
rect 307662 145024 307668 145036
rect 304500 144996 307668 145024
rect 304500 144984 304506 144996
rect 307662 144984 307668 144996
rect 307720 144984 307726 145036
rect 171962 144916 171968 144968
rect 172020 144956 172026 144968
rect 214006 144956 214012 144968
rect 172020 144928 214012 144956
rect 172020 144916 172026 144928
rect 214006 144916 214012 144928
rect 214064 144916 214070 144968
rect 293402 144916 293408 144968
rect 293460 144956 293466 144968
rect 307478 144956 307484 144968
rect 293460 144928 307484 144956
rect 293460 144916 293466 144928
rect 307478 144916 307484 144928
rect 307536 144916 307542 144968
rect 252094 144848 252100 144900
rect 252152 144888 252158 144900
rect 264974 144888 264980 144900
rect 252152 144860 264980 144888
rect 252152 144848 252158 144860
rect 264974 144848 264980 144860
rect 265032 144848 265038 144900
rect 324314 144848 324320 144900
rect 324372 144888 324378 144900
rect 342438 144888 342444 144900
rect 324372 144860 342444 144888
rect 324372 144848 324378 144860
rect 342438 144848 342444 144860
rect 342496 144848 342502 144900
rect 252462 144780 252468 144832
rect 252520 144820 252526 144832
rect 260834 144820 260840 144832
rect 252520 144792 260840 144820
rect 252520 144780 252526 144792
rect 260834 144780 260840 144792
rect 260892 144780 260898 144832
rect 204990 143624 204996 143676
rect 205048 143664 205054 143676
rect 214006 143664 214012 143676
rect 205048 143636 214012 143664
rect 205048 143624 205054 143636
rect 214006 143624 214012 143636
rect 214064 143624 214070 143676
rect 188338 143556 188344 143608
rect 188396 143596 188402 143608
rect 213914 143596 213920 143608
rect 188396 143568 213920 143596
rect 188396 143556 188402 143568
rect 213914 143556 213920 143568
rect 213972 143556 213978 143608
rect 274082 143556 274088 143608
rect 274140 143596 274146 143608
rect 307662 143596 307668 143608
rect 274140 143568 307668 143596
rect 274140 143556 274146 143568
rect 307662 143556 307668 143568
rect 307720 143556 307726 143608
rect 323578 143488 323584 143540
rect 323636 143528 323642 143540
rect 324498 143528 324504 143540
rect 323636 143500 324504 143528
rect 323636 143488 323642 143500
rect 324498 143488 324504 143500
rect 324556 143488 324562 143540
rect 324590 143488 324596 143540
rect 324648 143528 324654 143540
rect 343726 143528 343732 143540
rect 324648 143500 343732 143528
rect 324648 143488 324654 143500
rect 343726 143488 343732 143500
rect 343784 143488 343790 143540
rect 324314 143420 324320 143472
rect 324372 143460 324378 143472
rect 336918 143460 336924 143472
rect 324372 143432 336924 143460
rect 324372 143420 324378 143432
rect 336918 143420 336924 143432
rect 336976 143420 336982 143472
rect 250622 142808 250628 142860
rect 250680 142848 250686 142860
rect 305086 142848 305092 142860
rect 250680 142820 305092 142848
rect 250680 142808 250686 142820
rect 305086 142808 305092 142820
rect 305144 142808 305150 142860
rect 256050 142264 256056 142316
rect 256108 142304 256114 142316
rect 307662 142304 307668 142316
rect 256108 142276 307668 142304
rect 256108 142264 256114 142276
rect 307662 142264 307668 142276
rect 307720 142264 307726 142316
rect 272610 142196 272616 142248
rect 272668 142236 272674 142248
rect 307570 142236 307576 142248
rect 272668 142208 307576 142236
rect 272668 142196 272674 142208
rect 307570 142196 307576 142208
rect 307628 142196 307634 142248
rect 195238 142128 195244 142180
rect 195296 142168 195302 142180
rect 213914 142168 213920 142180
rect 195296 142140 213920 142168
rect 195296 142128 195302 142140
rect 213914 142128 213920 142140
rect 213972 142128 213978 142180
rect 324590 142060 324596 142112
rect 324648 142100 324654 142112
rect 345198 142100 345204 142112
rect 324648 142072 345204 142100
rect 324648 142060 324654 142072
rect 345198 142060 345204 142072
rect 345256 142060 345262 142112
rect 324314 141992 324320 142044
rect 324372 142032 324378 142044
rect 336734 142032 336740 142044
rect 324372 142004 336740 142032
rect 324372 141992 324378 142004
rect 336734 141992 336740 142004
rect 336792 141992 336798 142044
rect 171778 141380 171784 141432
rect 171836 141420 171842 141432
rect 209038 141420 209044 141432
rect 171836 141392 209044 141420
rect 171836 141380 171842 141392
rect 209038 141380 209044 141392
rect 209096 141380 209102 141432
rect 253290 141380 253296 141432
rect 253348 141420 253354 141432
rect 307018 141420 307024 141432
rect 253348 141392 307024 141420
rect 253348 141380 253354 141392
rect 307018 141380 307024 141392
rect 307076 141380 307082 141432
rect 210510 140836 210516 140888
rect 210568 140876 210574 140888
rect 214006 140876 214012 140888
rect 210568 140848 214012 140876
rect 210568 140836 210574 140848
rect 214006 140836 214012 140848
rect 214064 140836 214070 140888
rect 280982 140836 280988 140888
rect 281040 140876 281046 140888
rect 306926 140876 306932 140888
rect 281040 140848 306932 140876
rect 281040 140836 281046 140848
rect 306926 140836 306932 140848
rect 306984 140836 306990 140888
rect 206278 140768 206284 140820
rect 206336 140808 206342 140820
rect 213914 140808 213920 140820
rect 206336 140780 213920 140808
rect 206336 140768 206342 140780
rect 213914 140768 213920 140780
rect 213972 140768 213978 140820
rect 252094 140700 252100 140752
rect 252152 140740 252158 140752
rect 281534 140740 281540 140752
rect 252152 140712 281540 140740
rect 252152 140700 252158 140712
rect 281534 140700 281540 140712
rect 281592 140700 281598 140752
rect 324314 140700 324320 140752
rect 324372 140740 324378 140752
rect 338298 140740 338304 140752
rect 324372 140712 338304 140740
rect 324372 140700 324378 140712
rect 338298 140700 338304 140712
rect 338356 140700 338362 140752
rect 177758 140020 177764 140072
rect 177816 140060 177822 140072
rect 216030 140060 216036 140072
rect 177816 140032 216036 140060
rect 177816 140020 177822 140032
rect 216030 140020 216036 140032
rect 216088 140020 216094 140072
rect 252278 139816 252284 139868
rect 252336 139856 252342 139868
rect 260374 139856 260380 139868
rect 252336 139828 260380 139856
rect 252336 139816 252342 139828
rect 260374 139816 260380 139828
rect 260432 139816 260438 139868
rect 286318 139544 286324 139596
rect 286376 139584 286382 139596
rect 307662 139584 307668 139596
rect 286376 139556 307668 139584
rect 286376 139544 286382 139556
rect 307662 139544 307668 139556
rect 307720 139544 307726 139596
rect 271138 139476 271144 139528
rect 271196 139516 271202 139528
rect 307570 139516 307576 139528
rect 271196 139488 307576 139516
rect 271196 139476 271202 139488
rect 307570 139476 307576 139488
rect 307628 139476 307634 139528
rect 206370 139408 206376 139460
rect 206428 139448 206434 139460
rect 213914 139448 213920 139460
rect 206428 139420 213920 139448
rect 206428 139408 206434 139420
rect 213914 139408 213920 139420
rect 213972 139408 213978 139460
rect 260282 139408 260288 139460
rect 260340 139448 260346 139460
rect 307478 139448 307484 139460
rect 260340 139420 307484 139448
rect 260340 139408 260346 139420
rect 307478 139408 307484 139420
rect 307536 139408 307542 139460
rect 324314 139340 324320 139392
rect 324372 139380 324378 139392
rect 339678 139380 339684 139392
rect 324372 139352 339684 139380
rect 324372 139340 324378 139352
rect 339678 139340 339684 139352
rect 339736 139340 339742 139392
rect 472618 139340 472624 139392
rect 472676 139380 472682 139392
rect 580166 139380 580172 139392
rect 472676 139352 580172 139380
rect 472676 139340 472682 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 287882 138116 287888 138168
rect 287940 138156 287946 138168
rect 307662 138156 307668 138168
rect 287940 138128 307668 138156
rect 287940 138116 287946 138128
rect 307662 138116 307668 138128
rect 307720 138116 307726 138168
rect 170490 138048 170496 138100
rect 170548 138088 170554 138100
rect 213914 138088 213920 138100
rect 170548 138060 213920 138088
rect 170548 138048 170554 138060
rect 213914 138048 213920 138060
rect 213972 138048 213978 138100
rect 261570 138048 261576 138100
rect 261628 138088 261634 138100
rect 307570 138088 307576 138100
rect 261628 138060 307576 138088
rect 261628 138048 261634 138060
rect 307570 138048 307576 138060
rect 307628 138048 307634 138100
rect 166258 137980 166264 138032
rect 166316 138020 166322 138032
rect 214006 138020 214012 138032
rect 166316 137992 214012 138020
rect 166316 137980 166322 137992
rect 214006 137980 214012 137992
rect 214064 137980 214070 138032
rect 250438 137980 250444 138032
rect 250496 138020 250502 138032
rect 307478 138020 307484 138032
rect 250496 137992 307484 138020
rect 250496 137980 250502 137992
rect 307478 137980 307484 137992
rect 307536 137980 307542 138032
rect 252370 137912 252376 137964
rect 252428 137952 252434 137964
rect 278866 137952 278872 137964
rect 252428 137924 278872 137952
rect 252428 137912 252434 137924
rect 278866 137912 278872 137924
rect 278924 137912 278930 137964
rect 324406 137912 324412 137964
rect 324464 137952 324470 137964
rect 343910 137952 343916 137964
rect 324464 137924 343916 137952
rect 324464 137912 324470 137924
rect 343910 137912 343916 137924
rect 343968 137912 343974 137964
rect 252094 137844 252100 137896
rect 252152 137884 252158 137896
rect 273254 137884 273260 137896
rect 252152 137856 273260 137884
rect 252152 137844 252158 137856
rect 273254 137844 273260 137856
rect 273312 137844 273318 137896
rect 324314 137844 324320 137896
rect 324372 137884 324378 137896
rect 335538 137884 335544 137896
rect 324372 137856 335544 137884
rect 324372 137844 324378 137856
rect 335538 137844 335544 137856
rect 335596 137844 335602 137896
rect 252462 137776 252468 137828
rect 252520 137816 252526 137828
rect 267826 137816 267832 137828
rect 252520 137788 267832 137816
rect 252520 137776 252526 137788
rect 267826 137776 267832 137788
rect 267884 137776 267890 137828
rect 167730 137232 167736 137284
rect 167788 137272 167794 137284
rect 211798 137272 211804 137284
rect 167788 137244 211804 137272
rect 167788 137232 167794 137244
rect 211798 137232 211804 137244
rect 211856 137232 211862 137284
rect 252186 137096 252192 137148
rect 252244 137136 252250 137148
rect 259086 137136 259092 137148
rect 252244 137108 259092 137136
rect 252244 137096 252250 137108
rect 259086 137096 259092 137108
rect 259144 137096 259150 137148
rect 280890 136756 280896 136808
rect 280948 136796 280954 136808
rect 307570 136796 307576 136808
rect 280948 136768 307576 136796
rect 280948 136756 280954 136768
rect 307570 136756 307576 136768
rect 307628 136756 307634 136808
rect 258810 136688 258816 136740
rect 258868 136728 258874 136740
rect 306558 136728 306564 136740
rect 258868 136700 306564 136728
rect 258868 136688 258874 136700
rect 306558 136688 306564 136700
rect 306616 136688 306622 136740
rect 177298 136620 177304 136672
rect 177356 136660 177362 136672
rect 213914 136660 213920 136672
rect 177356 136632 213920 136660
rect 177356 136620 177362 136632
rect 213914 136620 213920 136632
rect 213972 136620 213978 136672
rect 249058 136620 249064 136672
rect 249116 136660 249122 136672
rect 307662 136660 307668 136672
rect 249116 136632 307668 136660
rect 249116 136620 249122 136632
rect 307662 136620 307668 136632
rect 307720 136620 307726 136672
rect 252370 136552 252376 136604
rect 252428 136592 252434 136604
rect 288066 136592 288072 136604
rect 252428 136564 288072 136592
rect 252428 136552 252434 136564
rect 288066 136552 288072 136564
rect 288124 136552 288130 136604
rect 324406 136552 324412 136604
rect 324464 136592 324470 136604
rect 341058 136592 341064 136604
rect 324464 136564 341064 136592
rect 324464 136552 324470 136564
rect 341058 136552 341064 136564
rect 341116 136552 341122 136604
rect 252094 136484 252100 136536
rect 252152 136524 252158 136536
rect 282270 136524 282276 136536
rect 252152 136496 282276 136524
rect 252152 136484 252158 136496
rect 282270 136484 282276 136496
rect 282328 136484 282334 136536
rect 252462 136416 252468 136468
rect 252520 136456 252526 136468
rect 264422 136456 264428 136468
rect 252520 136428 264428 136456
rect 252520 136416 252526 136428
rect 264422 136416 264428 136428
rect 264480 136416 264486 136468
rect 324314 136348 324320 136400
rect 324372 136388 324378 136400
rect 327258 136388 327264 136400
rect 324372 136360 327264 136388
rect 324372 136348 324378 136360
rect 327258 136348 327264 136360
rect 327316 136348 327322 136400
rect 251910 135872 251916 135924
rect 251968 135912 251974 135924
rect 290458 135912 290464 135924
rect 251968 135884 290464 135912
rect 251968 135872 251974 135884
rect 290458 135872 290464 135884
rect 290516 135872 290522 135924
rect 282362 135464 282368 135516
rect 282420 135504 282426 135516
rect 307478 135504 307484 135516
rect 282420 135476 307484 135504
rect 282420 135464 282426 135476
rect 307478 135464 307484 135476
rect 307536 135464 307542 135516
rect 297450 135396 297456 135448
rect 297508 135436 297514 135448
rect 307662 135436 307668 135448
rect 297508 135408 307668 135436
rect 297508 135396 297514 135408
rect 307662 135396 307668 135408
rect 307720 135396 307726 135448
rect 193858 135328 193864 135380
rect 193916 135368 193922 135380
rect 214006 135368 214012 135380
rect 193916 135340 214012 135368
rect 193916 135328 193922 135340
rect 214006 135328 214012 135340
rect 214064 135328 214070 135380
rect 290550 135328 290556 135380
rect 290608 135368 290614 135380
rect 307570 135368 307576 135380
rect 290608 135340 307576 135368
rect 290608 135328 290614 135340
rect 307570 135328 307576 135340
rect 307628 135328 307634 135380
rect 169018 135260 169024 135312
rect 169076 135300 169082 135312
rect 213914 135300 213920 135312
rect 169076 135272 213920 135300
rect 169076 135260 169082 135272
rect 213914 135260 213920 135272
rect 213972 135260 213978 135312
rect 304258 135260 304264 135312
rect 304316 135300 304322 135312
rect 307662 135300 307668 135312
rect 304316 135272 307668 135300
rect 304316 135260 304322 135272
rect 307662 135260 307668 135272
rect 307720 135260 307726 135312
rect 251634 135192 251640 135244
rect 251692 135232 251698 135244
rect 294598 135232 294604 135244
rect 251692 135204 294604 135232
rect 251692 135192 251698 135204
rect 294598 135192 294604 135204
rect 294656 135192 294662 135244
rect 252462 135124 252468 135176
rect 252520 135164 252526 135176
rect 269850 135164 269856 135176
rect 252520 135136 269856 135164
rect 252520 135124 252526 135136
rect 269850 135124 269856 135136
rect 269908 135124 269914 135176
rect 294690 134036 294696 134088
rect 294748 134076 294754 134088
rect 307662 134076 307668 134088
rect 294748 134048 307668 134076
rect 294748 134036 294754 134048
rect 307662 134036 307668 134048
rect 307720 134036 307726 134088
rect 289354 133968 289360 134020
rect 289412 134008 289418 134020
rect 307478 134008 307484 134020
rect 289412 133980 307484 134008
rect 289412 133968 289418 133980
rect 307478 133968 307484 133980
rect 307536 133968 307542 134020
rect 189810 133900 189816 133952
rect 189868 133940 189874 133952
rect 213914 133940 213920 133952
rect 189868 133912 213920 133940
rect 189868 133900 189874 133912
rect 213914 133900 213920 133912
rect 213972 133900 213978 133952
rect 270034 133900 270040 133952
rect 270092 133940 270098 133952
rect 307570 133940 307576 133952
rect 270092 133912 307576 133940
rect 270092 133900 270098 133912
rect 307570 133900 307576 133912
rect 307628 133900 307634 133952
rect 251450 133832 251456 133884
rect 251508 133872 251514 133884
rect 280798 133872 280804 133884
rect 251508 133844 280804 133872
rect 251508 133832 251514 133844
rect 280798 133832 280804 133844
rect 280856 133832 280862 133884
rect 252462 133764 252468 133816
rect 252520 133804 252526 133816
rect 271230 133804 271236 133816
rect 252520 133776 271236 133804
rect 252520 133764 252526 133776
rect 271230 133764 271236 133776
rect 271288 133764 271294 133816
rect 252002 133696 252008 133748
rect 252060 133736 252066 133748
rect 261662 133736 261668 133748
rect 252060 133708 261668 133736
rect 252060 133696 252066 133708
rect 261662 133696 261668 133708
rect 261720 133696 261726 133748
rect 271414 133152 271420 133204
rect 271472 133192 271478 133204
rect 307110 133192 307116 133204
rect 271472 133164 307116 133192
rect 271472 133152 271478 133164
rect 307110 133152 307116 133164
rect 307168 133152 307174 133204
rect 302970 132608 302976 132660
rect 303028 132648 303034 132660
rect 307570 132648 307576 132660
rect 303028 132620 307576 132648
rect 303028 132608 303034 132620
rect 307570 132608 307576 132620
rect 307628 132608 307634 132660
rect 293218 132540 293224 132592
rect 293276 132580 293282 132592
rect 307662 132580 307668 132592
rect 293276 132552 307668 132580
rect 293276 132540 293282 132552
rect 307662 132540 307668 132552
rect 307720 132540 307726 132592
rect 173250 132472 173256 132524
rect 173308 132512 173314 132524
rect 213914 132512 213920 132524
rect 173308 132484 213920 132512
rect 173308 132472 173314 132484
rect 213914 132472 213920 132484
rect 213972 132472 213978 132524
rect 282270 132472 282276 132524
rect 282328 132512 282334 132524
rect 307386 132512 307392 132524
rect 282328 132484 307392 132512
rect 282328 132472 282334 132484
rect 307386 132472 307392 132484
rect 307444 132472 307450 132524
rect 252462 132404 252468 132456
rect 252520 132444 252526 132456
rect 265618 132444 265624 132456
rect 252520 132416 265624 132444
rect 252520 132404 252526 132416
rect 265618 132404 265624 132416
rect 265676 132404 265682 132456
rect 324314 132404 324320 132456
rect 324372 132444 324378 132456
rect 347866 132444 347872 132456
rect 324372 132416 347872 132444
rect 324372 132404 324378 132416
rect 347866 132404 347872 132416
rect 347924 132404 347930 132456
rect 251542 132132 251548 132184
rect 251600 132172 251606 132184
rect 254854 132172 254860 132184
rect 251600 132144 254860 132172
rect 251600 132132 251606 132144
rect 254854 132132 254860 132144
rect 254912 132132 254918 132184
rect 202230 131112 202236 131164
rect 202288 131152 202294 131164
rect 213914 131152 213920 131164
rect 202288 131124 213920 131152
rect 202288 131112 202294 131124
rect 213914 131112 213920 131124
rect 213972 131112 213978 131164
rect 266998 131112 267004 131164
rect 267056 131152 267062 131164
rect 307662 131152 307668 131164
rect 267056 131124 307668 131152
rect 267056 131112 267062 131124
rect 307662 131112 307668 131124
rect 307720 131112 307726 131164
rect 252462 131044 252468 131096
rect 252520 131084 252526 131096
rect 271322 131084 271328 131096
rect 252520 131056 271328 131084
rect 252520 131044 252526 131056
rect 271322 131044 271328 131056
rect 271380 131044 271386 131096
rect 324314 131044 324320 131096
rect 324372 131084 324378 131096
rect 350626 131084 350632 131096
rect 324372 131056 350632 131084
rect 324372 131044 324378 131056
rect 350626 131044 350632 131056
rect 350684 131044 350690 131096
rect 251542 130976 251548 131028
rect 251600 131016 251606 131028
rect 267090 131016 267096 131028
rect 251600 130988 267096 131016
rect 251600 130976 251606 130988
rect 267090 130976 267096 130988
rect 267148 130976 267154 131028
rect 324406 130976 324412 131028
rect 324464 131016 324470 131028
rect 328730 131016 328736 131028
rect 324464 130988 328736 131016
rect 324464 130976 324470 130988
rect 328730 130976 328736 130988
rect 328788 130976 328794 131028
rect 183002 130364 183008 130416
rect 183060 130404 183066 130416
rect 214742 130404 214748 130416
rect 183060 130376 214748 130404
rect 183060 130364 183066 130376
rect 214742 130364 214748 130376
rect 214800 130364 214806 130416
rect 283650 129888 283656 129940
rect 283708 129928 283714 129940
rect 307662 129928 307668 129940
rect 283708 129900 307668 129928
rect 283708 129888 283714 129900
rect 307662 129888 307668 129900
rect 307720 129888 307726 129940
rect 273898 129820 273904 129872
rect 273956 129860 273962 129872
rect 307570 129860 307576 129872
rect 273956 129832 307576 129860
rect 273956 129820 273962 129832
rect 307570 129820 307576 129832
rect 307628 129820 307634 129872
rect 171778 129752 171784 129804
rect 171836 129792 171842 129804
rect 213914 129792 213920 129804
rect 171836 129764 213920 129792
rect 171836 129752 171842 129764
rect 213914 129752 213920 129764
rect 213972 129752 213978 129804
rect 268470 129752 268476 129804
rect 268528 129792 268534 129804
rect 306742 129792 306748 129804
rect 268528 129764 306748 129792
rect 268528 129752 268534 129764
rect 306742 129752 306748 129764
rect 306800 129752 306806 129804
rect 251726 129684 251732 129736
rect 251784 129724 251790 129736
rect 283558 129724 283564 129736
rect 251784 129696 283564 129724
rect 251784 129684 251790 129696
rect 283558 129684 283564 129696
rect 283616 129684 283622 129736
rect 324314 129684 324320 129736
rect 324372 129724 324378 129736
rect 351914 129724 351920 129736
rect 324372 129696 351920 129724
rect 324372 129684 324378 129696
rect 351914 129684 351920 129696
rect 351972 129684 351978 129736
rect 252002 129616 252008 129668
rect 252060 129656 252066 129668
rect 275278 129656 275284 129668
rect 252060 129628 275284 129656
rect 252060 129616 252066 129628
rect 275278 129616 275284 129628
rect 275336 129616 275342 129668
rect 324406 129616 324412 129668
rect 324464 129656 324470 129668
rect 328638 129656 328644 129668
rect 324464 129628 328644 129656
rect 324464 129616 324470 129628
rect 328638 129616 328644 129628
rect 328696 129616 328702 129668
rect 252462 129548 252468 129600
rect 252520 129588 252526 129600
rect 262858 129588 262864 129600
rect 252520 129560 262864 129588
rect 252520 129548 252526 129560
rect 262858 129548 262864 129560
rect 262916 129548 262922 129600
rect 297358 128460 297364 128512
rect 297416 128500 297422 128512
rect 307662 128500 307668 128512
rect 297416 128472 307668 128500
rect 297416 128460 297422 128472
rect 307662 128460 307668 128472
rect 307720 128460 307726 128512
rect 276658 128392 276664 128444
rect 276716 128432 276722 128444
rect 307386 128432 307392 128444
rect 276716 128404 307392 128432
rect 276716 128392 276722 128404
rect 307386 128392 307392 128404
rect 307444 128392 307450 128444
rect 174538 128324 174544 128376
rect 174596 128364 174602 128376
rect 213914 128364 213920 128376
rect 174596 128336 213920 128364
rect 174596 128324 174602 128336
rect 213914 128324 213920 128336
rect 213972 128324 213978 128376
rect 275370 128324 275376 128376
rect 275428 128364 275434 128376
rect 307570 128364 307576 128376
rect 275428 128336 307576 128364
rect 275428 128324 275434 128336
rect 307570 128324 307576 128336
rect 307628 128324 307634 128376
rect 252370 128256 252376 128308
rect 252428 128296 252434 128308
rect 291930 128296 291936 128308
rect 252428 128268 291936 128296
rect 252428 128256 252434 128268
rect 291930 128256 291936 128268
rect 291988 128256 291994 128308
rect 324314 128256 324320 128308
rect 324372 128296 324378 128308
rect 328454 128296 328460 128308
rect 324372 128268 328460 128296
rect 324372 128256 324378 128268
rect 328454 128256 328460 128268
rect 328512 128256 328518 128308
rect 252462 128188 252468 128240
rect 252520 128228 252526 128240
rect 278222 128228 278228 128240
rect 252520 128200 278228 128228
rect 252520 128188 252526 128200
rect 278222 128188 278228 128200
rect 278280 128188 278286 128240
rect 252002 128120 252008 128172
rect 252060 128160 252066 128172
rect 269942 128160 269948 128172
rect 252060 128132 269948 128160
rect 252060 128120 252066 128132
rect 269942 128120 269948 128132
rect 270000 128120 270006 128172
rect 324406 127916 324412 127968
rect 324464 127956 324470 127968
rect 327166 127956 327172 127968
rect 324464 127928 327172 127956
rect 324464 127916 324470 127928
rect 327166 127916 327172 127928
rect 327224 127916 327230 127968
rect 251818 127576 251824 127628
rect 251876 127616 251882 127628
rect 261754 127616 261760 127628
rect 251876 127588 261760 127616
rect 251876 127576 251882 127588
rect 261754 127576 261760 127588
rect 261812 127576 261818 127628
rect 279510 127100 279516 127152
rect 279568 127140 279574 127152
rect 307110 127140 307116 127152
rect 279568 127112 307116 127140
rect 279568 127100 279574 127112
rect 307110 127100 307116 127112
rect 307168 127100 307174 127152
rect 188430 127032 188436 127084
rect 188488 127072 188494 127084
rect 213914 127072 213920 127084
rect 188488 127044 213920 127072
rect 188488 127032 188494 127044
rect 213914 127032 213920 127044
rect 213972 127032 213978 127084
rect 278130 127032 278136 127084
rect 278188 127072 278194 127084
rect 307662 127072 307668 127084
rect 278188 127044 307668 127072
rect 278188 127032 278194 127044
rect 307662 127032 307668 127044
rect 307720 127032 307726 127084
rect 170398 126964 170404 127016
rect 170456 127004 170462 127016
rect 214006 127004 214012 127016
rect 170456 126976 214012 127004
rect 170456 126964 170462 126976
rect 214006 126964 214012 126976
rect 214064 126964 214070 127016
rect 269850 126964 269856 127016
rect 269908 127004 269914 127016
rect 306742 127004 306748 127016
rect 269908 126976 306748 127004
rect 269908 126964 269914 126976
rect 306742 126964 306748 126976
rect 306800 126964 306806 127016
rect 252186 126896 252192 126948
rect 252244 126936 252250 126948
rect 278314 126936 278320 126948
rect 252244 126908 278320 126936
rect 252244 126896 252250 126908
rect 278314 126896 278320 126908
rect 278372 126896 278378 126948
rect 449158 126896 449164 126948
rect 449216 126936 449222 126948
rect 580166 126936 580172 126948
rect 449216 126908 580172 126936
rect 449216 126896 449222 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 252462 126692 252468 126744
rect 252520 126732 252526 126744
rect 257430 126732 257436 126744
rect 252520 126704 257436 126732
rect 252520 126692 252526 126704
rect 257430 126692 257436 126704
rect 257488 126692 257494 126744
rect 251266 126216 251272 126268
rect 251324 126256 251330 126268
rect 300118 126256 300124 126268
rect 251324 126228 300124 126256
rect 251324 126216 251330 126228
rect 300118 126216 300124 126228
rect 300176 126216 300182 126268
rect 211890 125672 211896 125724
rect 211948 125712 211954 125724
rect 214466 125712 214472 125724
rect 211948 125684 214472 125712
rect 211948 125672 211954 125684
rect 214466 125672 214472 125684
rect 214524 125672 214530 125724
rect 290458 125672 290464 125724
rect 290516 125712 290522 125724
rect 307662 125712 307668 125724
rect 290516 125684 307668 125712
rect 290516 125672 290522 125684
rect 307662 125672 307668 125684
rect 307720 125672 307726 125724
rect 166442 125604 166448 125656
rect 166500 125644 166506 125656
rect 213914 125644 213920 125656
rect 166500 125616 213920 125644
rect 166500 125604 166506 125616
rect 213914 125604 213920 125616
rect 213972 125604 213978 125656
rect 271322 125604 271328 125656
rect 271380 125644 271386 125656
rect 306742 125644 306748 125656
rect 271380 125616 306748 125644
rect 271380 125604 271386 125616
rect 306742 125604 306748 125616
rect 306800 125604 306806 125656
rect 252186 125536 252192 125588
rect 252244 125576 252250 125588
rect 287790 125576 287796 125588
rect 252244 125548 287796 125576
rect 252244 125536 252250 125548
rect 287790 125536 287796 125548
rect 287848 125536 287854 125588
rect 324314 125536 324320 125588
rect 324372 125576 324378 125588
rect 342346 125576 342352 125588
rect 324372 125548 342352 125576
rect 324372 125536 324378 125548
rect 342346 125536 342352 125548
rect 342404 125536 342410 125588
rect 251174 125332 251180 125384
rect 251232 125372 251238 125384
rect 253290 125372 253296 125384
rect 251232 125344 253296 125372
rect 251232 125332 251238 125344
rect 253290 125332 253296 125344
rect 253348 125332 253354 125384
rect 252094 124856 252100 124908
rect 252152 124896 252158 124908
rect 265710 124896 265716 124908
rect 252152 124868 265716 124896
rect 252152 124856 252158 124868
rect 265710 124856 265716 124868
rect 265768 124856 265774 124908
rect 301498 124380 301504 124432
rect 301556 124420 301562 124432
rect 307662 124420 307668 124432
rect 301556 124392 307668 124420
rect 301556 124380 301562 124392
rect 307662 124380 307668 124392
rect 307720 124380 307726 124432
rect 287698 124312 287704 124364
rect 287756 124352 287762 124364
rect 306742 124352 306748 124364
rect 287756 124324 306748 124352
rect 287756 124312 287762 124324
rect 306742 124312 306748 124324
rect 306800 124312 306806 124364
rect 180058 124244 180064 124296
rect 180116 124284 180122 124296
rect 214006 124284 214012 124296
rect 180116 124256 214012 124284
rect 180116 124244 180122 124256
rect 214006 124244 214012 124256
rect 214064 124244 214070 124296
rect 265618 124244 265624 124296
rect 265676 124284 265682 124296
rect 307110 124284 307116 124296
rect 265676 124256 307116 124284
rect 265676 124244 265682 124256
rect 307110 124244 307116 124256
rect 307168 124244 307174 124296
rect 166350 124176 166356 124228
rect 166408 124216 166414 124228
rect 213914 124216 213920 124228
rect 166408 124188 213920 124216
rect 166408 124176 166414 124188
rect 213914 124176 213920 124188
rect 213972 124176 213978 124228
rect 260374 124176 260380 124228
rect 260432 124216 260438 124228
rect 307570 124216 307576 124228
rect 260432 124188 307576 124216
rect 260432 124176 260438 124188
rect 307570 124176 307576 124188
rect 307628 124176 307634 124228
rect 252462 124108 252468 124160
rect 252520 124148 252526 124160
rect 272518 124148 272524 124160
rect 252520 124120 272524 124148
rect 252520 124108 252526 124120
rect 272518 124108 272524 124120
rect 272576 124108 272582 124160
rect 324314 124108 324320 124160
rect 324372 124148 324378 124160
rect 340966 124148 340972 124160
rect 324372 124120 340972 124148
rect 324372 124108 324378 124120
rect 340966 124108 340972 124120
rect 341024 124108 341030 124160
rect 252002 123428 252008 123480
rect 252060 123468 252066 123480
rect 283742 123468 283748 123480
rect 252060 123440 283748 123468
rect 252060 123428 252066 123440
rect 283742 123428 283748 123440
rect 283800 123428 283806 123480
rect 211982 123360 211988 123412
rect 212040 123400 212046 123412
rect 214006 123400 214012 123412
rect 212040 123372 214012 123400
rect 212040 123360 212046 123372
rect 214006 123360 214012 123372
rect 214064 123360 214070 123412
rect 289170 122952 289176 123004
rect 289228 122992 289234 123004
rect 306558 122992 306564 123004
rect 289228 122964 306564 122992
rect 289228 122952 289234 122964
rect 306558 122952 306564 122964
rect 306616 122952 306622 123004
rect 283558 122884 283564 122936
rect 283616 122924 283622 122936
rect 307662 122924 307668 122936
rect 283616 122896 307668 122924
rect 283616 122884 283622 122896
rect 307662 122884 307668 122896
rect 307720 122884 307726 122936
rect 185578 122816 185584 122868
rect 185636 122856 185642 122868
rect 213914 122856 213920 122868
rect 185636 122828 213920 122856
rect 185636 122816 185642 122828
rect 213914 122816 213920 122828
rect 213972 122816 213978 122868
rect 252278 122816 252284 122868
rect 252336 122856 252342 122868
rect 258718 122856 258724 122868
rect 252336 122828 258724 122856
rect 252336 122816 252342 122828
rect 258718 122816 258724 122828
rect 258776 122816 258782 122868
rect 275278 122816 275284 122868
rect 275336 122856 275342 122868
rect 307570 122856 307576 122868
rect 275336 122828 307576 122856
rect 275336 122816 275342 122828
rect 307570 122816 307576 122828
rect 307628 122816 307634 122868
rect 252462 122748 252468 122800
rect 252520 122788 252526 122800
rect 289262 122788 289268 122800
rect 252520 122760 289268 122788
rect 252520 122748 252526 122760
rect 289262 122748 289268 122760
rect 289320 122748 289326 122800
rect 324314 122748 324320 122800
rect 324372 122788 324378 122800
rect 349338 122788 349344 122800
rect 324372 122760 349344 122788
rect 324372 122748 324378 122760
rect 349338 122748 349344 122760
rect 349396 122748 349402 122800
rect 252370 122680 252376 122732
rect 252428 122720 252434 122732
rect 279602 122720 279608 122732
rect 252428 122692 279608 122720
rect 252428 122680 252434 122692
rect 279602 122680 279608 122692
rect 279660 122680 279666 122732
rect 291930 121592 291936 121644
rect 291988 121632 291994 121644
rect 307570 121632 307576 121644
rect 291988 121604 307576 121632
rect 291988 121592 291994 121604
rect 307570 121592 307576 121604
rect 307628 121592 307634 121644
rect 186958 121524 186964 121576
rect 187016 121564 187022 121576
rect 213914 121564 213920 121576
rect 187016 121536 213920 121564
rect 187016 121524 187022 121536
rect 213914 121524 213920 121536
rect 213972 121524 213978 121576
rect 252462 121524 252468 121576
rect 252520 121564 252526 121576
rect 260098 121564 260104 121576
rect 252520 121536 260104 121564
rect 252520 121524 252526 121536
rect 260098 121524 260104 121536
rect 260156 121524 260162 121576
rect 284938 121524 284944 121576
rect 284996 121564 285002 121576
rect 307662 121564 307668 121576
rect 284996 121536 307668 121564
rect 284996 121524 285002 121536
rect 307662 121524 307668 121536
rect 307720 121524 307726 121576
rect 178770 121456 178776 121508
rect 178828 121496 178834 121508
rect 214006 121496 214012 121508
rect 178828 121468 214012 121496
rect 178828 121456 178834 121468
rect 214006 121456 214012 121468
rect 214064 121456 214070 121508
rect 278222 121456 278228 121508
rect 278280 121496 278286 121508
rect 306742 121496 306748 121508
rect 278280 121468 306748 121496
rect 278280 121456 278286 121468
rect 306742 121456 306748 121468
rect 306800 121456 306806 121508
rect 251910 121388 251916 121440
rect 251968 121428 251974 121440
rect 303062 121428 303068 121440
rect 251968 121400 303068 121428
rect 251968 121388 251974 121400
rect 303062 121388 303068 121400
rect 303120 121388 303126 121440
rect 324406 121388 324412 121440
rect 324464 121428 324470 121440
rect 345014 121428 345020 121440
rect 324464 121400 345020 121428
rect 324464 121388 324470 121400
rect 345014 121388 345020 121400
rect 345072 121388 345078 121440
rect 252462 121320 252468 121372
rect 252520 121360 252526 121372
rect 276842 121360 276848 121372
rect 252520 121332 276848 121360
rect 252520 121320 252526 121332
rect 276842 121320 276848 121332
rect 276900 121320 276906 121372
rect 324314 121320 324320 121372
rect 324372 121360 324378 121372
rect 330110 121360 330116 121372
rect 324372 121332 330116 121360
rect 324372 121320 324378 121332
rect 330110 121320 330116 121332
rect 330168 121320 330174 121372
rect 252094 121252 252100 121304
rect 252152 121292 252158 121304
rect 258902 121292 258908 121304
rect 252152 121264 258908 121292
rect 252152 121252 252158 121264
rect 258902 121252 258908 121264
rect 258960 121252 258966 121304
rect 302878 120232 302884 120284
rect 302936 120272 302942 120284
rect 306742 120272 306748 120284
rect 302936 120244 306748 120272
rect 302936 120232 302942 120244
rect 306742 120232 306748 120244
rect 306800 120232 306806 120284
rect 196710 120164 196716 120216
rect 196768 120204 196774 120216
rect 214006 120204 214012 120216
rect 196768 120176 214012 120204
rect 196768 120164 196774 120176
rect 214006 120164 214012 120176
rect 214064 120164 214070 120216
rect 280798 120164 280804 120216
rect 280856 120204 280862 120216
rect 307570 120204 307576 120216
rect 280856 120176 307576 120204
rect 280856 120164 280862 120176
rect 307570 120164 307576 120176
rect 307628 120164 307634 120216
rect 169110 120096 169116 120148
rect 169168 120136 169174 120148
rect 213914 120136 213920 120148
rect 169168 120108 213920 120136
rect 169168 120096 169174 120108
rect 213914 120096 213920 120108
rect 213972 120096 213978 120148
rect 273990 120096 273996 120148
rect 274048 120136 274054 120148
rect 307662 120136 307668 120148
rect 274048 120108 307668 120136
rect 274048 120096 274054 120108
rect 307662 120096 307668 120108
rect 307720 120096 307726 120148
rect 252370 120028 252376 120080
rect 252428 120068 252434 120080
rect 296070 120068 296076 120080
rect 252428 120040 296076 120068
rect 252428 120028 252434 120040
rect 296070 120028 296076 120040
rect 296128 120028 296134 120080
rect 324314 120028 324320 120080
rect 324372 120068 324378 120080
rect 338206 120068 338212 120080
rect 324372 120040 338212 120068
rect 324372 120028 324378 120040
rect 338206 120028 338212 120040
rect 338264 120028 338270 120080
rect 252462 119960 252468 120012
rect 252520 120000 252526 120012
rect 264330 120000 264336 120012
rect 252520 119972 264336 120000
rect 252520 119960 252526 119972
rect 264330 119960 264336 119972
rect 264388 119960 264394 120012
rect 261754 119348 261760 119400
rect 261812 119388 261818 119400
rect 307478 119388 307484 119400
rect 261812 119360 307484 119388
rect 261812 119348 261818 119360
rect 307478 119348 307484 119360
rect 307536 119348 307542 119400
rect 192570 118804 192576 118856
rect 192628 118844 192634 118856
rect 213914 118844 213920 118856
rect 192628 118816 213920 118844
rect 192628 118804 192634 118816
rect 213914 118804 213920 118816
rect 213972 118804 213978 118856
rect 173342 118736 173348 118788
rect 173400 118776 173406 118788
rect 214006 118776 214012 118788
rect 173400 118748 214012 118776
rect 173400 118736 173406 118748
rect 214006 118736 214012 118748
rect 214064 118736 214070 118788
rect 296162 118736 296168 118788
rect 296220 118776 296226 118788
rect 307662 118776 307668 118788
rect 296220 118748 307668 118776
rect 296220 118736 296226 118748
rect 307662 118736 307668 118748
rect 307720 118736 307726 118788
rect 167822 118668 167828 118720
rect 167880 118708 167886 118720
rect 214098 118708 214104 118720
rect 167880 118680 214104 118708
rect 167880 118668 167886 118680
rect 214098 118668 214104 118680
rect 214156 118668 214162 118720
rect 252462 118668 252468 118720
rect 252520 118708 252526 118720
rect 260190 118708 260196 118720
rect 252520 118680 260196 118708
rect 252520 118668 252526 118680
rect 260190 118668 260196 118680
rect 260248 118668 260254 118720
rect 294598 118668 294604 118720
rect 294656 118708 294662 118720
rect 306742 118708 306748 118720
rect 294656 118680 306748 118708
rect 294656 118668 294662 118680
rect 306742 118668 306748 118680
rect 306800 118668 306806 118720
rect 252094 118600 252100 118652
rect 252152 118640 252158 118652
rect 287974 118640 287980 118652
rect 252152 118612 287980 118640
rect 252152 118600 252158 118612
rect 287974 118600 287980 118612
rect 288032 118600 288038 118652
rect 324314 118600 324320 118652
rect 324372 118640 324378 118652
rect 336826 118640 336832 118652
rect 324372 118612 336832 118640
rect 324372 118600 324378 118612
rect 336826 118600 336832 118612
rect 336884 118600 336890 118652
rect 324406 118532 324412 118584
rect 324464 118572 324470 118584
rect 334066 118572 334072 118584
rect 324464 118544 334072 118572
rect 324464 118532 324470 118544
rect 334066 118532 334072 118544
rect 334124 118532 334130 118584
rect 251542 118396 251548 118448
rect 251600 118436 251606 118448
rect 257338 118436 257344 118448
rect 251600 118408 257344 118436
rect 251600 118396 251606 118408
rect 257338 118396 257344 118408
rect 257396 118396 257402 118448
rect 251818 117920 251824 117972
rect 251876 117960 251882 117972
rect 304350 117960 304356 117972
rect 251876 117932 304356 117960
rect 251876 117920 251882 117932
rect 304350 117920 304356 117932
rect 304408 117920 304414 117972
rect 203702 117376 203708 117428
rect 203760 117416 203766 117428
rect 214006 117416 214012 117428
rect 203760 117388 214012 117416
rect 203760 117376 203766 117388
rect 214006 117376 214012 117388
rect 214064 117376 214070 117428
rect 301682 117376 301688 117428
rect 301740 117416 301746 117428
rect 307662 117416 307668 117428
rect 301740 117388 307668 117416
rect 301740 117376 301746 117388
rect 307662 117376 307668 117388
rect 307720 117376 307726 117428
rect 167914 117308 167920 117360
rect 167972 117348 167978 117360
rect 213914 117348 213920 117360
rect 167972 117320 213920 117348
rect 167972 117308 167978 117320
rect 213914 117308 213920 117320
rect 213972 117308 213978 117360
rect 287790 117308 287796 117360
rect 287848 117348 287854 117360
rect 307478 117348 307484 117360
rect 287848 117320 307484 117348
rect 287848 117308 287854 117320
rect 307478 117308 307484 117320
rect 307536 117308 307542 117360
rect 252370 117240 252376 117292
rect 252428 117280 252434 117292
rect 285122 117280 285128 117292
rect 252428 117252 285128 117280
rect 252428 117240 252434 117252
rect 285122 117240 285128 117252
rect 285180 117240 285186 117292
rect 324314 117240 324320 117292
rect 324372 117280 324378 117292
rect 343634 117280 343640 117292
rect 324372 117252 343640 117280
rect 324372 117240 324378 117252
rect 343634 117240 343640 117252
rect 343692 117240 343698 117292
rect 324406 117172 324412 117224
rect 324464 117212 324470 117224
rect 335446 117212 335452 117224
rect 324464 117184 335452 117212
rect 324464 117172 324470 117184
rect 335446 117172 335452 117184
rect 335504 117172 335510 117224
rect 251542 116900 251548 116952
rect 251600 116940 251606 116952
rect 257522 116940 257528 116952
rect 251600 116912 257528 116940
rect 251600 116900 251606 116912
rect 257522 116900 257528 116912
rect 257580 116900 257586 116952
rect 251910 116560 251916 116612
rect 251968 116600 251974 116612
rect 263042 116600 263048 116612
rect 251968 116572 263048 116600
rect 251968 116560 251974 116572
rect 263042 116560 263048 116572
rect 263100 116560 263106 116612
rect 296070 116560 296076 116612
rect 296128 116600 296134 116612
rect 307202 116600 307208 116612
rect 296128 116572 307208 116600
rect 296128 116560 296134 116572
rect 307202 116560 307208 116572
rect 307260 116560 307266 116612
rect 189902 116016 189908 116068
rect 189960 116056 189966 116068
rect 214006 116056 214012 116068
rect 189960 116028 214012 116056
rect 189960 116016 189966 116028
rect 214006 116016 214012 116028
rect 214064 116016 214070 116068
rect 285030 116016 285036 116068
rect 285088 116056 285094 116068
rect 307478 116056 307484 116068
rect 285088 116028 307484 116056
rect 285088 116016 285094 116028
rect 307478 116016 307484 116028
rect 307536 116016 307542 116068
rect 187050 115948 187056 116000
rect 187108 115988 187114 116000
rect 213914 115988 213920 116000
rect 187108 115960 213920 115988
rect 187108 115948 187114 115960
rect 213914 115948 213920 115960
rect 213972 115948 213978 116000
rect 262858 115948 262864 116000
rect 262916 115988 262922 116000
rect 307662 115988 307668 116000
rect 262916 115960 307668 115988
rect 262916 115948 262922 115960
rect 307662 115948 307668 115960
rect 307720 115948 307726 116000
rect 252370 115880 252376 115932
rect 252428 115920 252434 115932
rect 295978 115920 295984 115932
rect 252428 115892 295984 115920
rect 252428 115880 252434 115892
rect 295978 115880 295984 115892
rect 296036 115880 296042 115932
rect 324314 115880 324320 115932
rect 324372 115920 324378 115932
rect 345106 115920 345112 115932
rect 324372 115892 345112 115920
rect 324372 115880 324378 115892
rect 345106 115880 345112 115892
rect 345164 115880 345170 115932
rect 251634 115812 251640 115864
rect 251692 115852 251698 115864
rect 254670 115852 254676 115864
rect 251692 115824 254676 115852
rect 251692 115812 251698 115824
rect 254670 115812 254676 115824
rect 254728 115812 254734 115864
rect 298830 114656 298836 114708
rect 298888 114696 298894 114708
rect 307570 114696 307576 114708
rect 298888 114668 307576 114696
rect 298888 114656 298894 114668
rect 307570 114656 307576 114668
rect 307628 114656 307634 114708
rect 185670 114588 185676 114640
rect 185728 114628 185734 114640
rect 213914 114628 213920 114640
rect 185728 114600 213920 114628
rect 185728 114588 185734 114600
rect 213914 114588 213920 114600
rect 213972 114588 213978 114640
rect 287974 114588 287980 114640
rect 288032 114628 288038 114640
rect 307662 114628 307668 114640
rect 288032 114600 307668 114628
rect 288032 114588 288038 114600
rect 307662 114588 307668 114600
rect 307720 114588 307726 114640
rect 182910 114520 182916 114572
rect 182968 114560 182974 114572
rect 214006 114560 214012 114572
rect 182968 114532 214012 114560
rect 182968 114520 182974 114532
rect 214006 114520 214012 114532
rect 214064 114520 214070 114572
rect 253290 114520 253296 114572
rect 253348 114560 253354 114572
rect 307478 114560 307484 114572
rect 253348 114532 307484 114560
rect 253348 114520 253354 114532
rect 307478 114520 307484 114532
rect 307536 114520 307542 114572
rect 252462 114452 252468 114504
rect 252520 114492 252526 114504
rect 261478 114492 261484 114504
rect 252520 114464 261484 114492
rect 252520 114452 252526 114464
rect 261478 114452 261484 114464
rect 261536 114452 261542 114504
rect 324406 114452 324412 114504
rect 324464 114492 324470 114504
rect 332686 114492 332692 114504
rect 324464 114464 332692 114492
rect 324464 114452 324470 114464
rect 332686 114452 332692 114464
rect 332744 114452 332750 114504
rect 324314 114384 324320 114436
rect 324372 114424 324378 114436
rect 331214 114424 331220 114436
rect 324372 114396 331220 114424
rect 324372 114384 324378 114396
rect 331214 114384 331220 114396
rect 331272 114384 331278 114436
rect 252462 113704 252468 113756
rect 252520 113744 252526 113756
rect 258994 113744 259000 113756
rect 252520 113716 259000 113744
rect 252520 113704 252526 113716
rect 258994 113704 259000 113716
rect 259052 113704 259058 113756
rect 251726 113364 251732 113416
rect 251784 113404 251790 113416
rect 253474 113404 253480 113416
rect 251784 113376 253480 113404
rect 251784 113364 251790 113376
rect 253474 113364 253480 113376
rect 253532 113364 253538 113416
rect 181438 113228 181444 113280
rect 181496 113268 181502 113280
rect 214006 113268 214012 113280
rect 181496 113240 214012 113268
rect 181496 113228 181502 113240
rect 214006 113228 214012 113240
rect 214064 113228 214070 113280
rect 264330 113228 264336 113280
rect 264388 113268 264394 113280
rect 307570 113268 307576 113280
rect 264388 113240 307576 113268
rect 264388 113228 264394 113240
rect 307570 113228 307576 113240
rect 307628 113228 307634 113280
rect 172054 113160 172060 113212
rect 172112 113200 172118 113212
rect 213914 113200 213920 113212
rect 172112 113172 213920 113200
rect 172112 113160 172118 113172
rect 213914 113160 213920 113172
rect 213972 113160 213978 113212
rect 260098 113160 260104 113212
rect 260156 113200 260162 113212
rect 307662 113200 307668 113212
rect 260156 113172 307668 113200
rect 260156 113160 260162 113172
rect 307662 113160 307668 113172
rect 307720 113160 307726 113212
rect 252094 113092 252100 113144
rect 252152 113132 252158 113144
rect 296070 113132 296076 113144
rect 252152 113104 296076 113132
rect 252152 113092 252158 113104
rect 296070 113092 296076 113104
rect 296128 113092 296134 113144
rect 324314 113092 324320 113144
rect 324372 113132 324378 113144
rect 338114 113132 338120 113144
rect 324372 113104 338120 113132
rect 324372 113092 324378 113104
rect 338114 113092 338120 113104
rect 338172 113092 338178 113144
rect 468478 113092 468484 113144
rect 468536 113132 468542 113144
rect 579798 113132 579804 113144
rect 468536 113104 579804 113132
rect 468536 113092 468542 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 252186 113024 252192 113076
rect 252244 113064 252250 113076
rect 255958 113064 255964 113076
rect 252244 113036 255964 113064
rect 252244 113024 252250 113036
rect 255958 113024 255964 113036
rect 256016 113024 256022 113076
rect 174630 112412 174636 112464
rect 174688 112452 174694 112464
rect 214926 112452 214932 112464
rect 174688 112424 214932 112452
rect 174688 112412 174694 112424
rect 214926 112412 214932 112424
rect 214984 112412 214990 112464
rect 252002 112412 252008 112464
rect 252060 112452 252066 112464
rect 304442 112452 304448 112464
rect 252060 112424 304448 112452
rect 252060 112412 252066 112424
rect 304442 112412 304448 112424
rect 304500 112412 304506 112464
rect 303062 111936 303068 111988
rect 303120 111976 303126 111988
rect 307294 111976 307300 111988
rect 303120 111948 307300 111976
rect 303120 111936 303126 111948
rect 307294 111936 307300 111948
rect 307352 111936 307358 111988
rect 167546 111868 167552 111920
rect 167604 111908 167610 111920
rect 167730 111908 167736 111920
rect 167604 111880 167736 111908
rect 167604 111868 167610 111880
rect 167730 111868 167736 111880
rect 167788 111868 167794 111920
rect 304350 111868 304356 111920
rect 304408 111908 304414 111920
rect 307662 111908 307668 111920
rect 304408 111880 307668 111908
rect 304408 111868 304414 111880
rect 307662 111868 307668 111880
rect 307720 111868 307726 111920
rect 177390 111800 177396 111852
rect 177448 111840 177454 111852
rect 213914 111840 213920 111852
rect 177448 111812 213920 111840
rect 177448 111800 177454 111812
rect 213914 111800 213920 111812
rect 213972 111800 213978 111852
rect 293310 111800 293316 111852
rect 293368 111840 293374 111852
rect 306558 111840 306564 111852
rect 293368 111812 306564 111840
rect 293368 111800 293374 111812
rect 306558 111800 306564 111812
rect 306616 111800 306622 111852
rect 167730 111732 167736 111784
rect 167788 111772 167794 111784
rect 207658 111772 207664 111784
rect 167788 111744 207664 111772
rect 167788 111732 167794 111744
rect 207658 111732 207664 111744
rect 207716 111732 207722 111784
rect 252370 111732 252376 111784
rect 252428 111772 252434 111784
rect 256234 111772 256240 111784
rect 252428 111744 256240 111772
rect 252428 111732 252434 111744
rect 256234 111732 256240 111744
rect 256292 111732 256298 111784
rect 324314 111732 324320 111784
rect 324372 111772 324378 111784
rect 339494 111772 339500 111784
rect 324372 111744 339500 111772
rect 324372 111732 324378 111744
rect 339494 111732 339500 111744
rect 339552 111732 339558 111784
rect 252278 111188 252284 111240
rect 252336 111228 252342 111240
rect 274174 111228 274180 111240
rect 252336 111200 274180 111228
rect 252336 111188 252342 111200
rect 274174 111188 274180 111200
rect 274232 111188 274238 111240
rect 256602 111120 256608 111172
rect 256660 111160 256666 111172
rect 282454 111160 282460 111172
rect 256660 111132 282460 111160
rect 256660 111120 256666 111132
rect 282454 111120 282460 111132
rect 282512 111120 282518 111172
rect 251910 111052 251916 111104
rect 251968 111092 251974 111104
rect 301774 111092 301780 111104
rect 251968 111064 301780 111092
rect 251968 111052 251974 111064
rect 301774 111052 301780 111064
rect 301832 111052 301838 111104
rect 300118 110576 300124 110628
rect 300176 110616 300182 110628
rect 306558 110616 306564 110628
rect 300176 110588 306564 110616
rect 300176 110576 300182 110588
rect 306558 110576 306564 110588
rect 306616 110576 306622 110628
rect 192662 110508 192668 110560
rect 192720 110548 192726 110560
rect 214006 110548 214012 110560
rect 192720 110520 214012 110548
rect 192720 110508 192726 110520
rect 214006 110508 214012 110520
rect 214064 110508 214070 110560
rect 295978 110508 295984 110560
rect 296036 110548 296042 110560
rect 307294 110548 307300 110560
rect 296036 110520 307300 110548
rect 296036 110508 296042 110520
rect 307294 110508 307300 110520
rect 307352 110508 307358 110560
rect 169202 110440 169208 110492
rect 169260 110480 169266 110492
rect 213914 110480 213920 110492
rect 169260 110452 213920 110480
rect 169260 110440 169266 110452
rect 213914 110440 213920 110452
rect 213972 110440 213978 110492
rect 283742 110440 283748 110492
rect 283800 110480 283806 110492
rect 306742 110480 306748 110492
rect 283800 110452 306748 110480
rect 283800 110440 283806 110452
rect 306742 110440 306748 110452
rect 306800 110440 306806 110492
rect 251450 110372 251456 110424
rect 251508 110412 251514 110424
rect 254578 110412 254584 110424
rect 251508 110384 254584 110412
rect 251508 110372 251514 110384
rect 254578 110372 254584 110384
rect 254636 110372 254642 110424
rect 324314 110372 324320 110424
rect 324372 110412 324378 110424
rect 332594 110412 332600 110424
rect 324372 110384 332600 110412
rect 324372 110372 324378 110384
rect 332594 110372 332600 110384
rect 332652 110372 332658 110424
rect 251542 110304 251548 110356
rect 251600 110344 251606 110356
rect 268562 110344 268568 110356
rect 251600 110316 268568 110344
rect 251600 110304 251606 110316
rect 268562 110304 268568 110316
rect 268620 110304 268626 110356
rect 252462 110236 252468 110288
rect 252520 110276 252526 110288
rect 298922 110276 298928 110288
rect 252520 110248 298928 110276
rect 252520 110236 252526 110248
rect 298922 110236 298928 110248
rect 298980 110236 298986 110288
rect 303154 109148 303160 109200
rect 303212 109188 303218 109200
rect 306742 109188 306748 109200
rect 303212 109160 306748 109188
rect 303212 109148 303218 109160
rect 306742 109148 306748 109160
rect 306800 109148 306806 109200
rect 296070 109080 296076 109132
rect 296128 109120 296134 109132
rect 307662 109120 307668 109132
rect 296128 109092 307668 109120
rect 296128 109080 296134 109092
rect 307662 109080 307668 109092
rect 307720 109080 307726 109132
rect 170582 109012 170588 109064
rect 170640 109052 170646 109064
rect 213914 109052 213920 109064
rect 170640 109024 213920 109052
rect 170640 109012 170646 109024
rect 213914 109012 213920 109024
rect 213972 109012 213978 109064
rect 272518 109012 272524 109064
rect 272576 109052 272582 109064
rect 307570 109052 307576 109064
rect 272576 109024 307576 109052
rect 272576 109012 272582 109024
rect 307570 109012 307576 109024
rect 307628 109012 307634 109064
rect 167730 108944 167736 108996
rect 167788 108984 167794 108996
rect 196802 108984 196808 108996
rect 167788 108956 196808 108984
rect 167788 108944 167794 108956
rect 196802 108944 196808 108956
rect 196860 108944 196866 108996
rect 251818 108944 251824 108996
rect 251876 108984 251882 108996
rect 300302 108984 300308 108996
rect 251876 108956 300308 108984
rect 251876 108944 251882 108956
rect 300302 108944 300308 108956
rect 300360 108944 300366 108996
rect 251174 108876 251180 108928
rect 251232 108916 251238 108928
rect 253198 108916 253204 108928
rect 251232 108888 253204 108916
rect 251232 108876 251238 108888
rect 253198 108876 253204 108888
rect 253256 108876 253262 108928
rect 324314 108876 324320 108928
rect 324372 108916 324378 108928
rect 339586 108916 339592 108928
rect 324372 108888 339592 108916
rect 324372 108876 324378 108888
rect 339586 108876 339592 108888
rect 339644 108876 339650 108928
rect 252554 108264 252560 108316
rect 252612 108304 252618 108316
rect 291838 108304 291844 108316
rect 252612 108276 291844 108304
rect 252612 108264 252618 108276
rect 291838 108264 291844 108276
rect 291896 108264 291902 108316
rect 255958 107856 255964 107908
rect 256016 107896 256022 107908
rect 307662 107896 307668 107908
rect 256016 107868 307668 107896
rect 256016 107856 256022 107868
rect 307662 107856 307668 107868
rect 307720 107856 307726 107908
rect 207658 107720 207664 107772
rect 207716 107760 207722 107772
rect 214006 107760 214012 107772
rect 207716 107732 214012 107760
rect 207716 107720 207722 107732
rect 214006 107720 214012 107732
rect 214064 107720 214070 107772
rect 300210 107720 300216 107772
rect 300268 107760 300274 107772
rect 307294 107760 307300 107772
rect 300268 107732 307300 107760
rect 300268 107720 300274 107732
rect 307294 107720 307300 107732
rect 307352 107720 307358 107772
rect 199378 107652 199384 107704
rect 199436 107692 199442 107704
rect 213914 107692 213920 107704
rect 199436 107664 213920 107692
rect 199436 107652 199442 107664
rect 213914 107652 213920 107664
rect 213972 107652 213978 107704
rect 301774 107652 301780 107704
rect 301832 107692 301838 107704
rect 307478 107692 307484 107704
rect 301832 107664 307484 107692
rect 301832 107652 301838 107664
rect 307478 107652 307484 107664
rect 307536 107652 307542 107704
rect 252370 107584 252376 107636
rect 252428 107624 252434 107636
rect 276750 107624 276756 107636
rect 252428 107596 276756 107624
rect 252428 107584 252434 107596
rect 276750 107584 276756 107596
rect 276808 107584 276814 107636
rect 252462 107516 252468 107568
rect 252520 107556 252526 107568
rect 269758 107556 269764 107568
rect 252520 107528 269764 107556
rect 252520 107516 252526 107528
rect 269758 107516 269764 107528
rect 269816 107516 269822 107568
rect 251542 107380 251548 107432
rect 251600 107420 251606 107432
rect 254762 107420 254768 107432
rect 251600 107392 254768 107420
rect 251600 107380 251606 107392
rect 254762 107380 254768 107392
rect 254820 107380 254826 107432
rect 292022 106972 292028 107024
rect 292080 107012 292086 107024
rect 307202 107012 307208 107024
rect 292080 106984 307208 107012
rect 292080 106972 292086 106984
rect 307202 106972 307208 106984
rect 307260 106972 307266 107024
rect 276106 106904 276112 106956
rect 276164 106944 276170 106956
rect 295334 106944 295340 106956
rect 276164 106916 295340 106944
rect 276164 106904 276170 106916
rect 295334 106904 295340 106916
rect 295392 106904 295398 106956
rect 304442 106428 304448 106480
rect 304500 106468 304506 106480
rect 307662 106468 307668 106480
rect 304500 106440 307668 106468
rect 304500 106428 304506 106440
rect 307662 106428 307668 106440
rect 307720 106428 307726 106480
rect 211798 106360 211804 106412
rect 211856 106400 211862 106412
rect 214466 106400 214472 106412
rect 211856 106372 214472 106400
rect 211856 106360 211862 106372
rect 214466 106360 214472 106372
rect 214524 106360 214530 106412
rect 298922 106360 298928 106412
rect 298980 106400 298986 106412
rect 307478 106400 307484 106412
rect 298980 106372 307484 106400
rect 298980 106360 298986 106372
rect 307478 106360 307484 106372
rect 307536 106360 307542 106412
rect 167730 106292 167736 106344
rect 167788 106332 167794 106344
rect 213914 106332 213920 106344
rect 167788 106304 213920 106332
rect 167788 106292 167794 106304
rect 213914 106292 213920 106304
rect 213972 106292 213978 106344
rect 261478 106292 261484 106344
rect 261536 106332 261542 106344
rect 307294 106332 307300 106344
rect 261536 106304 307300 106332
rect 261536 106292 261542 106304
rect 307294 106292 307300 106304
rect 307352 106292 307358 106344
rect 324314 106224 324320 106276
rect 324372 106264 324378 106276
rect 347774 106264 347780 106276
rect 324372 106236 347780 106264
rect 324372 106224 324378 106236
rect 347774 106224 347780 106236
rect 347832 106224 347838 106276
rect 251174 106156 251180 106208
rect 251232 106196 251238 106208
rect 253382 106196 253388 106208
rect 251232 106168 253388 106196
rect 251232 106156 251238 106168
rect 253382 106156 253388 106168
rect 253440 106156 253446 106208
rect 252370 105680 252376 105732
rect 252428 105720 252434 105732
rect 256142 105720 256148 105732
rect 252428 105692 256148 105720
rect 252428 105680 252434 105692
rect 256142 105680 256148 105692
rect 256200 105680 256206 105732
rect 252186 105612 252192 105664
rect 252244 105652 252250 105664
rect 306006 105652 306012 105664
rect 252244 105624 306012 105652
rect 252244 105612 252250 105624
rect 306006 105612 306012 105624
rect 306064 105612 306070 105664
rect 251634 105544 251640 105596
rect 251692 105584 251698 105596
rect 306098 105584 306104 105596
rect 251692 105556 306104 105584
rect 251692 105544 251698 105556
rect 306098 105544 306104 105556
rect 306156 105544 306162 105596
rect 293494 105000 293500 105052
rect 293552 105040 293558 105052
rect 307662 105040 307668 105052
rect 293552 105012 307668 105040
rect 293552 105000 293558 105012
rect 307662 105000 307668 105012
rect 307720 105000 307726 105052
rect 196894 104932 196900 104984
rect 196952 104972 196958 104984
rect 213914 104972 213920 104984
rect 196952 104944 213920 104972
rect 196952 104932 196958 104944
rect 213914 104932 213920 104944
rect 213972 104932 213978 104984
rect 194042 104864 194048 104916
rect 194100 104904 194106 104916
rect 214006 104904 214012 104916
rect 194100 104876 214012 104904
rect 194100 104864 194106 104876
rect 214006 104864 214012 104876
rect 214064 104864 214070 104916
rect 252462 104796 252468 104848
rect 252520 104836 252526 104848
rect 293402 104836 293408 104848
rect 252520 104808 293408 104836
rect 252520 104796 252526 104808
rect 293402 104796 293408 104808
rect 293460 104796 293466 104848
rect 324314 104796 324320 104848
rect 324372 104836 324378 104848
rect 356054 104836 356060 104848
rect 324372 104808 356060 104836
rect 324372 104796 324378 104808
rect 356054 104796 356060 104808
rect 356112 104796 356118 104848
rect 324314 104660 324320 104712
rect 324372 104700 324378 104712
rect 327074 104700 327080 104712
rect 324372 104672 327080 104700
rect 324372 104660 324378 104672
rect 327074 104660 327080 104672
rect 327132 104660 327138 104712
rect 252278 104116 252284 104168
rect 252336 104156 252342 104168
rect 305730 104156 305736 104168
rect 252336 104128 305736 104156
rect 252336 104116 252342 104128
rect 305730 104116 305736 104128
rect 305788 104116 305794 104168
rect 304534 103640 304540 103692
rect 304592 103680 304598 103692
rect 307662 103680 307668 103692
rect 304592 103652 307668 103680
rect 304592 103640 304598 103652
rect 307662 103640 307668 103652
rect 307720 103640 307726 103692
rect 202322 103572 202328 103624
rect 202380 103612 202386 103624
rect 213914 103612 213920 103624
rect 202380 103584 213920 103612
rect 202380 103572 202386 103584
rect 213914 103572 213920 103584
rect 213972 103572 213978 103624
rect 296254 103572 296260 103624
rect 296312 103612 296318 103624
rect 307478 103612 307484 103624
rect 296312 103584 307484 103612
rect 296312 103572 296318 103584
rect 307478 103572 307484 103584
rect 307536 103572 307542 103624
rect 199470 103504 199476 103556
rect 199528 103544 199534 103556
rect 214006 103544 214012 103556
rect 199528 103516 214012 103544
rect 199528 103504 199534 103516
rect 214006 103504 214012 103516
rect 214064 103504 214070 103556
rect 278314 103504 278320 103556
rect 278372 103544 278378 103556
rect 307570 103544 307576 103556
rect 278372 103516 307576 103544
rect 278372 103504 278378 103516
rect 307570 103504 307576 103516
rect 307628 103504 307634 103556
rect 252370 103436 252376 103488
rect 252428 103476 252434 103488
rect 274082 103476 274088 103488
rect 252428 103448 274088 103476
rect 252428 103436 252434 103448
rect 274082 103436 274088 103448
rect 274140 103436 274146 103488
rect 252462 103368 252468 103420
rect 252520 103408 252526 103420
rect 271414 103408 271420 103420
rect 252520 103380 271420 103408
rect 252520 103368 252526 103380
rect 271414 103368 271420 103380
rect 271472 103368 271478 103420
rect 299014 102280 299020 102332
rect 299072 102320 299078 102332
rect 306558 102320 306564 102332
rect 299072 102292 306564 102320
rect 299072 102280 299078 102292
rect 306558 102280 306564 102292
rect 306616 102280 306622 102332
rect 207750 102212 207756 102264
rect 207808 102252 207814 102264
rect 214006 102252 214012 102264
rect 207808 102224 214012 102252
rect 207808 102212 207814 102224
rect 214006 102212 214012 102224
rect 214064 102212 214070 102264
rect 274174 102212 274180 102264
rect 274232 102252 274238 102264
rect 307570 102252 307576 102264
rect 274232 102224 307576 102252
rect 274232 102212 274238 102224
rect 307570 102212 307576 102224
rect 307628 102212 307634 102264
rect 191190 102144 191196 102196
rect 191248 102184 191254 102196
rect 213914 102184 213920 102196
rect 191248 102156 213920 102184
rect 191248 102144 191254 102156
rect 213914 102144 213920 102156
rect 213972 102144 213978 102196
rect 271230 102144 271236 102196
rect 271288 102184 271294 102196
rect 307662 102184 307668 102196
rect 271288 102156 307668 102184
rect 271288 102144 271294 102156
rect 307662 102144 307668 102156
rect 307720 102144 307726 102196
rect 252462 102076 252468 102128
rect 252520 102116 252526 102128
rect 272610 102116 272616 102128
rect 252520 102088 272616 102116
rect 252520 102076 252526 102088
rect 272610 102076 272616 102088
rect 272668 102076 272674 102128
rect 252002 101192 252008 101244
rect 252060 101232 252066 101244
rect 256050 101232 256056 101244
rect 252060 101204 256056 101232
rect 252060 101192 252066 101204
rect 256050 101192 256056 101204
rect 256108 101192 256114 101244
rect 254578 100920 254584 100972
rect 254636 100960 254642 100972
rect 307662 100960 307668 100972
rect 254636 100932 307668 100960
rect 254636 100920 254642 100932
rect 307662 100920 307668 100932
rect 307720 100920 307726 100972
rect 297542 100852 297548 100904
rect 297600 100892 297606 100904
rect 306558 100892 306564 100904
rect 297600 100864 306564 100892
rect 297600 100852 297606 100864
rect 306558 100852 306564 100864
rect 306616 100852 306622 100904
rect 260190 100784 260196 100836
rect 260248 100824 260254 100836
rect 307662 100824 307668 100836
rect 260248 100796 307668 100824
rect 260248 100784 260254 100796
rect 307662 100784 307668 100796
rect 307720 100784 307726 100836
rect 206462 100716 206468 100768
rect 206520 100756 206526 100768
rect 213914 100756 213920 100768
rect 206520 100728 213920 100756
rect 206520 100716 206526 100728
rect 213914 100716 213920 100728
rect 213972 100716 213978 100768
rect 252094 100648 252100 100700
rect 252152 100688 252158 100700
rect 292022 100688 292028 100700
rect 252152 100660 292028 100688
rect 252152 100648 252158 100660
rect 292022 100648 292028 100660
rect 292080 100648 292086 100700
rect 467098 100648 467104 100700
rect 467156 100688 467162 100700
rect 580166 100688 580172 100700
rect 467156 100660 580172 100688
rect 467156 100648 467162 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 252462 100580 252468 100632
rect 252520 100620 252526 100632
rect 280982 100620 280988 100632
rect 252520 100592 280988 100620
rect 252520 100580 252526 100592
rect 280982 100580 280988 100592
rect 281040 100580 281046 100632
rect 170674 99968 170680 100020
rect 170732 100008 170738 100020
rect 214650 100008 214656 100020
rect 170732 99980 214656 100008
rect 170732 99968 170738 99980
rect 214650 99968 214656 99980
rect 214708 99968 214714 100020
rect 294782 99492 294788 99544
rect 294840 99532 294846 99544
rect 306558 99532 306564 99544
rect 294840 99504 306564 99532
rect 294840 99492 294846 99504
rect 306558 99492 306564 99504
rect 306616 99492 306622 99544
rect 291838 99424 291844 99476
rect 291896 99464 291902 99476
rect 306742 99464 306748 99476
rect 291896 99436 306748 99464
rect 291896 99424 291902 99436
rect 306742 99424 306748 99436
rect 306800 99424 306806 99476
rect 198182 99356 198188 99408
rect 198240 99396 198246 99408
rect 213914 99396 213920 99408
rect 198240 99368 213920 99396
rect 198240 99356 198246 99368
rect 213914 99356 213920 99368
rect 213972 99356 213978 99408
rect 258718 99356 258724 99408
rect 258776 99396 258782 99408
rect 307662 99396 307668 99408
rect 258776 99368 307668 99396
rect 258776 99356 258782 99368
rect 307662 99356 307668 99368
rect 307720 99356 307726 99408
rect 252462 99288 252468 99340
rect 252520 99328 252526 99340
rect 262950 99328 262956 99340
rect 252520 99300 262956 99328
rect 252520 99288 252526 99300
rect 262950 99288 262956 99300
rect 263008 99288 263014 99340
rect 252370 99220 252376 99272
rect 252428 99260 252434 99272
rect 261754 99260 261760 99272
rect 252428 99232 261760 99260
rect 252428 99220 252434 99232
rect 261754 99220 261760 99232
rect 261812 99220 261818 99272
rect 252462 98132 252468 98184
rect 252520 98172 252526 98184
rect 260282 98172 260288 98184
rect 252520 98144 260288 98172
rect 252520 98132 252526 98144
rect 260282 98132 260288 98144
rect 260340 98132 260346 98184
rect 196802 98064 196808 98116
rect 196860 98104 196866 98116
rect 213914 98104 213920 98116
rect 196860 98076 213920 98104
rect 196860 98064 196866 98076
rect 213914 98064 213920 98076
rect 213972 98064 213978 98116
rect 269758 98064 269764 98116
rect 269816 98104 269822 98116
rect 306742 98104 306748 98116
rect 269816 98076 306748 98104
rect 269816 98064 269822 98076
rect 306742 98064 306748 98076
rect 306800 98064 306806 98116
rect 166534 97996 166540 98048
rect 166592 98036 166598 98048
rect 214006 98036 214012 98048
rect 166592 98008 214012 98036
rect 166592 97996 166598 98008
rect 214006 97996 214012 98008
rect 214064 97996 214070 98048
rect 261662 97996 261668 98048
rect 261720 98036 261726 98048
rect 307662 98036 307668 98048
rect 261720 98008 307668 98036
rect 261720 97996 261726 98008
rect 307662 97996 307668 98008
rect 307720 97996 307726 98048
rect 169294 97248 169300 97300
rect 169352 97288 169358 97300
rect 214558 97288 214564 97300
rect 169352 97260 214564 97288
rect 169352 97248 169358 97260
rect 214558 97248 214564 97260
rect 214616 97248 214622 97300
rect 289262 96772 289268 96824
rect 289320 96812 289326 96824
rect 307662 96812 307668 96824
rect 289320 96784 307668 96812
rect 289320 96772 289326 96784
rect 307662 96772 307668 96784
rect 307720 96772 307726 96824
rect 253198 96704 253204 96756
rect 253256 96744 253262 96756
rect 307570 96744 307576 96756
rect 253256 96716 307576 96744
rect 253256 96704 253262 96716
rect 307570 96704 307576 96716
rect 307628 96704 307634 96756
rect 207842 96636 207848 96688
rect 207900 96676 207906 96688
rect 213914 96676 213920 96688
rect 207900 96648 213920 96676
rect 207900 96636 207906 96648
rect 213914 96636 213920 96648
rect 213972 96636 213978 96688
rect 250530 96636 250536 96688
rect 250588 96676 250594 96688
rect 307662 96676 307668 96688
rect 250588 96648 307668 96676
rect 250588 96636 250594 96648
rect 307662 96636 307668 96648
rect 307720 96636 307726 96688
rect 165522 95888 165528 95940
rect 165580 95928 165586 95940
rect 214098 95928 214104 95940
rect 165580 95900 214104 95928
rect 165580 95888 165586 95900
rect 214098 95888 214104 95900
rect 214156 95888 214162 95940
rect 251818 95208 251824 95260
rect 251876 95248 251882 95260
rect 306926 95248 306932 95260
rect 251876 95220 306932 95248
rect 251876 95208 251882 95220
rect 306926 95208 306932 95220
rect 306984 95208 306990 95260
rect 178678 95140 178684 95192
rect 178736 95180 178742 95192
rect 321462 95180 321468 95192
rect 178736 95152 321468 95180
rect 178736 95140 178742 95152
rect 321462 95140 321468 95152
rect 321520 95140 321526 95192
rect 59262 95004 59268 95056
rect 59320 95044 59326 95056
rect 199470 95044 199476 95056
rect 59320 95016 199476 95044
rect 59320 95004 59326 95016
rect 199470 95004 199476 95016
rect 199528 95004 199534 95056
rect 246942 94460 246948 94512
rect 247000 94500 247006 94512
rect 299566 94500 299572 94512
rect 247000 94472 299572 94500
rect 247000 94460 247006 94472
rect 299566 94460 299572 94472
rect 299624 94460 299630 94512
rect 133138 94052 133144 94104
rect 133196 94092 133202 94104
rect 182818 94092 182824 94104
rect 133196 94064 182824 94092
rect 133196 94052 133202 94064
rect 182818 94052 182824 94064
rect 182876 94052 182882 94104
rect 113726 93984 113732 94036
rect 113784 94024 113790 94036
rect 173342 94024 173348 94036
rect 113784 93996 173348 94024
rect 113784 93984 113790 93996
rect 173342 93984 173348 93996
rect 173400 93984 173406 94036
rect 115474 93916 115480 93968
rect 115532 93956 115538 93968
rect 177298 93956 177304 93968
rect 115532 93928 177304 93956
rect 115532 93916 115538 93928
rect 177298 93916 177304 93928
rect 177356 93916 177362 93968
rect 102042 93848 102048 93900
rect 102100 93888 102106 93900
rect 171778 93888 171784 93900
rect 102100 93860 171784 93888
rect 102100 93848 102106 93860
rect 171778 93848 171784 93860
rect 171836 93848 171842 93900
rect 62022 93780 62028 93832
rect 62080 93820 62086 93832
rect 207750 93820 207756 93832
rect 62080 93792 207756 93820
rect 62080 93780 62086 93792
rect 207750 93780 207756 93792
rect 207808 93780 207814 93832
rect 209038 93780 209044 93832
rect 209096 93820 209102 93832
rect 321646 93820 321652 93832
rect 209096 93792 321652 93820
rect 209096 93780 209102 93792
rect 321646 93780 321652 93792
rect 321704 93780 321710 93832
rect 151722 93372 151728 93424
rect 151780 93412 151786 93424
rect 171870 93412 171876 93424
rect 151780 93384 171876 93412
rect 151780 93372 151786 93384
rect 171870 93372 171876 93384
rect 171928 93372 171934 93424
rect 134426 93304 134432 93356
rect 134484 93344 134490 93356
rect 167638 93344 167644 93356
rect 134484 93316 167644 93344
rect 134484 93304 134490 93316
rect 167638 93304 167644 93316
rect 167696 93304 167702 93356
rect 118050 93236 118056 93288
rect 118108 93276 118114 93288
rect 170490 93276 170496 93288
rect 118108 93248 170496 93276
rect 118108 93236 118114 93248
rect 170490 93236 170496 93248
rect 170548 93236 170554 93288
rect 110138 93168 110144 93220
rect 110196 93208 110202 93220
rect 167914 93208 167920 93220
rect 110196 93180 167920 93208
rect 110196 93168 110202 93180
rect 167914 93168 167920 93180
rect 167972 93168 167978 93220
rect 119522 93100 119528 93152
rect 119580 93140 119586 93152
rect 178770 93140 178776 93152
rect 119580 93112 178776 93140
rect 119580 93100 119586 93112
rect 178770 93100 178776 93112
rect 178828 93100 178834 93152
rect 238754 93100 238760 93152
rect 238812 93140 238818 93152
rect 250622 93140 250628 93152
rect 238812 93112 250628 93140
rect 238812 93100 238818 93112
rect 250622 93100 250628 93112
rect 250680 93100 250686 93152
rect 88978 92420 88984 92472
rect 89036 92460 89042 92472
rect 165522 92460 165528 92472
rect 89036 92432 165528 92460
rect 89036 92420 89042 92432
rect 165522 92420 165528 92432
rect 165580 92420 165586 92472
rect 173158 92420 173164 92472
rect 173216 92460 173222 92472
rect 324590 92460 324596 92472
rect 173216 92432 324596 92460
rect 173216 92420 173222 92432
rect 324590 92420 324596 92432
rect 324648 92420 324654 92472
rect 130746 92352 130752 92404
rect 130804 92392 130810 92404
rect 193950 92392 193956 92404
rect 130804 92364 193956 92392
rect 130804 92352 130810 92364
rect 193950 92352 193956 92364
rect 194008 92352 194014 92404
rect 125870 92284 125876 92336
rect 125928 92324 125934 92336
rect 183002 92324 183008 92336
rect 125928 92296 183008 92324
rect 125928 92284 125934 92296
rect 183002 92284 183008 92296
rect 183060 92284 183066 92336
rect 116762 92216 116768 92268
rect 116820 92256 116826 92268
rect 170674 92256 170680 92268
rect 116820 92228 170680 92256
rect 116820 92216 116826 92228
rect 170674 92216 170680 92228
rect 170732 92216 170738 92268
rect 151538 92148 151544 92200
rect 151596 92188 151602 92200
rect 203610 92188 203616 92200
rect 151596 92160 203616 92188
rect 151596 92148 151602 92160
rect 203610 92148 203616 92160
rect 203668 92148 203674 92200
rect 119706 92080 119712 92132
rect 119764 92120 119770 92132
rect 166258 92120 166264 92132
rect 119764 92092 166264 92120
rect 119764 92080 119770 92092
rect 166258 92080 166264 92092
rect 166316 92080 166322 92132
rect 3142 91740 3148 91792
rect 3200 91780 3206 91792
rect 25498 91780 25504 91792
rect 3200 91752 25504 91780
rect 3200 91740 3206 91752
rect 25498 91740 25504 91752
rect 25556 91740 25562 91792
rect 228358 91740 228364 91792
rect 228416 91780 228422 91792
rect 278314 91780 278320 91792
rect 228416 91752 278320 91780
rect 228416 91740 228422 91752
rect 278314 91740 278320 91752
rect 278372 91740 278378 91792
rect 88058 91196 88064 91248
rect 88116 91236 88122 91248
rect 111058 91236 111064 91248
rect 88116 91208 111064 91236
rect 88116 91196 88122 91208
rect 111058 91196 111064 91208
rect 111116 91196 111122 91248
rect 74810 91128 74816 91180
rect 74868 91168 74874 91180
rect 100018 91168 100024 91180
rect 74868 91140 100024 91168
rect 74868 91128 74874 91140
rect 100018 91128 100024 91140
rect 100076 91128 100082 91180
rect 100570 91128 100576 91180
rect 100628 91168 100634 91180
rect 116578 91168 116584 91180
rect 100628 91140 116584 91168
rect 100628 91128 100634 91140
rect 116578 91128 116584 91140
rect 116636 91128 116642 91180
rect 85758 91060 85764 91112
rect 85816 91100 85822 91112
rect 128998 91100 129004 91112
rect 85816 91072 129004 91100
rect 85816 91060 85822 91072
rect 128998 91060 129004 91072
rect 129056 91060 129062 91112
rect 128170 90992 128176 91044
rect 128228 91032 128234 91044
rect 188338 91032 188344 91044
rect 128228 91004 188344 91032
rect 128228 90992 128234 91004
rect 188338 90992 188344 91004
rect 188396 90992 188402 91044
rect 112162 90924 112168 90976
rect 112220 90964 112226 90976
rect 169018 90964 169024 90976
rect 112220 90936 169024 90964
rect 112220 90924 112226 90936
rect 169018 90924 169024 90936
rect 169076 90924 169082 90976
rect 115474 90856 115480 90908
rect 115532 90896 115538 90908
rect 167822 90896 167828 90908
rect 115532 90868 167828 90896
rect 115532 90856 115538 90868
rect 167822 90856 167828 90868
rect 167880 90856 167886 90908
rect 126514 90788 126520 90840
rect 126572 90828 126578 90840
rect 166442 90828 166448 90840
rect 126572 90800 166448 90828
rect 126572 90788 126578 90800
rect 166442 90788 166448 90800
rect 166500 90788 166506 90840
rect 152918 90720 152924 90772
rect 152976 90760 152982 90772
rect 191098 90760 191104 90772
rect 152976 90732 191104 90760
rect 152976 90720 152982 90732
rect 191098 90720 191104 90732
rect 191156 90720 191162 90772
rect 151354 90652 151360 90704
rect 151412 90692 151418 90704
rect 184198 90692 184204 90704
rect 151412 90664 184204 90692
rect 151412 90652 151418 90664
rect 184198 90652 184204 90664
rect 184256 90652 184262 90704
rect 256050 90312 256056 90364
rect 256108 90352 256114 90364
rect 266354 90352 266360 90364
rect 256108 90324 266360 90352
rect 256108 90312 256114 90324
rect 266354 90312 266360 90324
rect 266412 90312 266418 90364
rect 67450 89632 67456 89684
rect 67508 89672 67514 89684
rect 214834 89672 214840 89684
rect 67508 89644 214840 89672
rect 67508 89632 67514 89644
rect 214834 89632 214840 89644
rect 214892 89632 214898 89684
rect 66070 89564 66076 89616
rect 66128 89604 66134 89616
rect 207842 89604 207848 89616
rect 66128 89576 207848 89604
rect 66128 89564 66134 89576
rect 207842 89564 207848 89576
rect 207900 89564 207906 89616
rect 109218 89496 109224 89548
rect 109276 89536 109282 89548
rect 189902 89536 189908 89548
rect 109276 89508 189908 89536
rect 109276 89496 109282 89508
rect 189902 89496 189908 89508
rect 189960 89496 189966 89548
rect 101858 89428 101864 89480
rect 101916 89468 101922 89480
rect 177390 89468 177396 89480
rect 101916 89440 177396 89468
rect 101916 89428 101922 89440
rect 177390 89428 177396 89440
rect 177448 89428 177454 89480
rect 122834 89360 122840 89412
rect 122892 89400 122898 89412
rect 166350 89400 166356 89412
rect 122892 89372 166356 89400
rect 122892 89360 122898 89372
rect 166350 89360 166356 89372
rect 166408 89360 166414 89412
rect 132218 89292 132224 89344
rect 132276 89332 132282 89344
rect 171962 89332 171968 89344
rect 132276 89304 171968 89332
rect 132276 89292 132282 89304
rect 171962 89292 171968 89304
rect 172020 89292 172026 89344
rect 224218 89156 224224 89208
rect 224276 89196 224282 89208
rect 260374 89196 260380 89208
rect 224276 89168 260380 89196
rect 224276 89156 224282 89168
rect 260374 89156 260380 89168
rect 260432 89156 260438 89208
rect 242894 89088 242900 89140
rect 242952 89128 242958 89140
rect 296714 89128 296720 89140
rect 242952 89100 296720 89128
rect 242952 89088 242958 89100
rect 296714 89088 296720 89100
rect 296772 89088 296778 89140
rect 176378 89020 176384 89072
rect 176436 89060 176442 89072
rect 245654 89060 245660 89072
rect 176436 89032 245660 89060
rect 176436 89020 176442 89032
rect 245654 89020 245660 89032
rect 245712 89020 245718 89072
rect 204898 88952 204904 89004
rect 204956 88992 204962 89004
rect 378778 88992 378784 89004
rect 204956 88964 378784 88992
rect 204956 88952 204962 88964
rect 378778 88952 378784 88964
rect 378836 88952 378842 89004
rect 39942 88272 39948 88324
rect 40000 88312 40006 88324
rect 323026 88312 323032 88324
rect 40000 88284 323032 88312
rect 40000 88272 40006 88284
rect 323026 88272 323032 88284
rect 323084 88272 323090 88324
rect 111426 88204 111432 88256
rect 111484 88244 111490 88256
rect 203702 88244 203708 88256
rect 111484 88216 203708 88244
rect 111484 88204 111490 88216
rect 203702 88204 203708 88216
rect 203760 88204 203766 88256
rect 100478 88136 100484 88188
rect 100536 88176 100542 88188
rect 192662 88176 192668 88188
rect 100536 88148 192668 88176
rect 100536 88136 100542 88148
rect 192662 88136 192668 88148
rect 192720 88136 192726 88188
rect 136450 88068 136456 88120
rect 136508 88108 136514 88120
rect 198090 88108 198096 88120
rect 136508 88080 198096 88108
rect 136508 88068 136514 88080
rect 198090 88068 198096 88080
rect 198148 88068 198154 88120
rect 124030 88000 124036 88052
rect 124088 88040 124094 88052
rect 180058 88040 180064 88052
rect 124088 88012 180064 88040
rect 124088 88000 124094 88012
rect 180058 88000 180064 88012
rect 180116 88000 180122 88052
rect 203610 87592 203616 87644
rect 203668 87632 203674 87644
rect 307110 87632 307116 87644
rect 203668 87604 307116 87632
rect 203668 87592 203674 87604
rect 307110 87592 307116 87604
rect 307168 87592 307174 87644
rect 67726 86912 67732 86964
rect 67784 86952 67790 86964
rect 214650 86952 214656 86964
rect 67784 86924 214656 86952
rect 67784 86912 67790 86924
rect 214650 86912 214656 86924
rect 214708 86912 214714 86964
rect 122098 86844 122104 86896
rect 122156 86884 122162 86896
rect 206370 86884 206376 86896
rect 122156 86856 206376 86884
rect 122156 86844 122162 86856
rect 206370 86844 206376 86856
rect 206428 86844 206434 86896
rect 107838 86776 107844 86828
rect 107896 86816 107902 86828
rect 187050 86816 187056 86828
rect 107896 86788 187056 86816
rect 107896 86776 107902 86788
rect 187050 86776 187056 86788
rect 187108 86776 187114 86828
rect 118234 86708 118240 86760
rect 118292 86748 118298 86760
rect 186958 86748 186964 86760
rect 118292 86720 186964 86748
rect 118292 86708 118298 86720
rect 186958 86708 186964 86720
rect 187016 86708 187022 86760
rect 238018 86300 238024 86352
rect 238076 86340 238082 86352
rect 251266 86340 251272 86352
rect 238076 86312 251272 86340
rect 238076 86300 238082 86312
rect 251266 86300 251272 86312
rect 251324 86300 251330 86352
rect 216582 86232 216588 86284
rect 216640 86272 216646 86284
rect 310514 86272 310520 86284
rect 216640 86244 310520 86272
rect 216640 86232 216646 86244
rect 310514 86232 310520 86244
rect 310572 86232 310578 86284
rect 104618 85484 104624 85536
rect 104676 85524 104682 85536
rect 202230 85524 202236 85536
rect 104676 85496 202236 85524
rect 104676 85484 104682 85496
rect 202230 85484 202236 85496
rect 202288 85484 202294 85536
rect 120442 85416 120448 85468
rect 120500 85456 120506 85468
rect 213178 85456 213184 85468
rect 120500 85428 213184 85456
rect 120500 85416 120506 85428
rect 213178 85416 213184 85428
rect 213236 85416 213242 85468
rect 105722 85348 105728 85400
rect 105780 85388 105786 85400
rect 185670 85388 185676 85400
rect 105780 85360 185676 85388
rect 105780 85348 105786 85360
rect 185670 85348 185676 85360
rect 185728 85348 185734 85400
rect 104342 85280 104348 85332
rect 104400 85320 104406 85332
rect 181438 85320 181444 85332
rect 104400 85292 181444 85320
rect 104400 85280 104406 85292
rect 181438 85280 181444 85292
rect 181496 85280 181502 85332
rect 97258 85212 97264 85264
rect 97316 85252 97322 85264
rect 170582 85252 170588 85264
rect 97316 85224 170588 85252
rect 97316 85212 97322 85224
rect 170582 85212 170588 85224
rect 170640 85212 170646 85264
rect 115842 85144 115848 85196
rect 115900 85184 115906 85196
rect 169110 85184 169116 85196
rect 115900 85156 169116 85184
rect 115900 85144 115906 85156
rect 169110 85144 169116 85156
rect 169168 85144 169174 85196
rect 308490 84804 308496 84856
rect 308548 84844 308554 84856
rect 317414 84844 317420 84856
rect 308548 84816 317420 84844
rect 308548 84804 308554 84816
rect 317414 84804 317420 84816
rect 317472 84804 317478 84856
rect 92382 84124 92388 84176
rect 92440 84164 92446 84176
rect 211798 84164 211804 84176
rect 92440 84136 211804 84164
rect 92440 84124 92446 84136
rect 211798 84124 211804 84136
rect 211856 84124 211862 84176
rect 99098 84056 99104 84108
rect 99156 84096 99162 84108
rect 169202 84096 169208 84108
rect 99156 84068 169208 84096
rect 99156 84056 99162 84068
rect 169202 84056 169208 84068
rect 169260 84056 169266 84108
rect 103422 83988 103428 84040
rect 103480 84028 103486 84040
rect 172054 84028 172060 84040
rect 103480 84000 172060 84028
rect 103480 83988 103486 84000
rect 172054 83988 172060 84000
rect 172112 83988 172118 84040
rect 126790 83920 126796 83972
rect 126848 83960 126854 83972
rect 195238 83960 195244 83972
rect 126848 83932 195244 83960
rect 126848 83920 126854 83932
rect 195238 83920 195244 83932
rect 195296 83920 195302 83972
rect 121362 83852 121368 83904
rect 121420 83892 121426 83904
rect 185578 83892 185584 83904
rect 121420 83864 185584 83892
rect 121420 83852 121426 83864
rect 185578 83852 185584 83864
rect 185636 83852 185642 83904
rect 258074 83512 258080 83564
rect 258132 83552 258138 83564
rect 284294 83552 284300 83564
rect 258132 83524 284300 83552
rect 258132 83512 258138 83524
rect 284294 83512 284300 83524
rect 284352 83512 284358 83564
rect 309870 83512 309876 83564
rect 309928 83552 309934 83564
rect 324314 83552 324320 83564
rect 309928 83524 324320 83552
rect 309928 83512 309934 83524
rect 324314 83512 324320 83524
rect 324372 83512 324378 83564
rect 207014 83444 207020 83496
rect 207072 83484 207078 83496
rect 319438 83484 319444 83496
rect 207072 83456 319444 83484
rect 207072 83444 207078 83456
rect 319438 83444 319444 83456
rect 319496 83444 319502 83496
rect 50982 82764 50988 82816
rect 51040 82804 51046 82816
rect 321554 82804 321560 82816
rect 51040 82776 321560 82804
rect 51040 82764 51046 82776
rect 321554 82764 321560 82776
rect 321612 82764 321618 82816
rect 124122 82696 124128 82748
rect 124180 82736 124186 82748
rect 210510 82736 210516 82748
rect 124180 82708 210516 82736
rect 124180 82696 124186 82708
rect 210510 82696 210516 82708
rect 210568 82696 210574 82748
rect 110322 82628 110328 82680
rect 110380 82668 110386 82680
rect 189810 82668 189816 82680
rect 110380 82640 189816 82668
rect 110380 82628 110386 82640
rect 189810 82628 189816 82640
rect 189868 82628 189874 82680
rect 113082 82560 113088 82612
rect 113140 82600 113146 82612
rect 192570 82600 192576 82612
rect 113140 82572 192576 82600
rect 113140 82560 113146 82572
rect 192570 82560 192576 82572
rect 192628 82560 192634 82612
rect 108942 82492 108948 82544
rect 109000 82532 109006 82544
rect 173250 82532 173256 82544
rect 109000 82504 173256 82532
rect 109000 82492 109006 82504
rect 173250 82492 173256 82504
rect 173308 82492 173314 82544
rect 251266 82084 251272 82136
rect 251324 82124 251330 82136
rect 293954 82124 293960 82136
rect 251324 82096 293960 82124
rect 251324 82084 251330 82096
rect 293954 82084 293960 82096
rect 294012 82084 294018 82136
rect 95050 81336 95056 81388
rect 95108 81376 95114 81388
rect 199378 81376 199384 81388
rect 95108 81348 199384 81376
rect 95108 81336 95114 81348
rect 199378 81336 199384 81348
rect 199436 81336 199442 81388
rect 86862 81268 86868 81320
rect 86920 81308 86926 81320
rect 166534 81308 166540 81320
rect 86920 81280 166540 81308
rect 86920 81268 86926 81280
rect 166534 81268 166540 81280
rect 166592 81268 166598 81320
rect 117222 81200 117228 81252
rect 117280 81240 117286 81252
rect 196710 81240 196716 81252
rect 117280 81212 196716 81240
rect 117280 81200 117286 81212
rect 196710 81200 196716 81212
rect 196768 81200 196774 81252
rect 114462 81132 114468 81184
rect 114520 81172 114526 81184
rect 193858 81172 193864 81184
rect 114520 81144 193864 81172
rect 114520 81132 114526 81144
rect 193858 81132 193864 81144
rect 193916 81132 193922 81184
rect 129642 81064 129648 81116
rect 129700 81104 129706 81116
rect 204990 81104 204996 81116
rect 129700 81076 204996 81104
rect 129700 81064 129706 81076
rect 204990 81064 204996 81076
rect 205048 81064 205054 81116
rect 177850 80724 177856 80776
rect 177908 80764 177914 80776
rect 247678 80764 247684 80776
rect 177908 80736 247684 80764
rect 177908 80724 177914 80736
rect 247678 80724 247684 80736
rect 247736 80724 247742 80776
rect 198734 80656 198740 80708
rect 198792 80696 198798 80708
rect 269942 80696 269948 80708
rect 198792 80668 269948 80696
rect 198792 80656 198798 80668
rect 269942 80656 269948 80668
rect 270000 80656 270006 80708
rect 298738 80656 298744 80708
rect 298796 80696 298802 80708
rect 322934 80696 322940 80708
rect 298796 80668 322940 80696
rect 298796 80656 298802 80668
rect 322934 80656 322940 80668
rect 322992 80656 322998 80708
rect 95142 79976 95148 80028
rect 95200 80016 95206 80028
rect 207658 80016 207664 80028
rect 95200 79988 207664 80016
rect 95200 79976 95206 79988
rect 207658 79976 207664 79988
rect 207716 79976 207722 80028
rect 116578 79908 116584 79960
rect 116636 79948 116642 79960
rect 214742 79948 214748 79960
rect 116636 79920 214748 79948
rect 116636 79908 116642 79920
rect 214742 79908 214748 79920
rect 214800 79908 214806 79960
rect 122742 79840 122748 79892
rect 122800 79880 122806 79892
rect 211982 79880 211988 79892
rect 122800 79852 211988 79880
rect 122800 79840 122806 79852
rect 211982 79840 211988 79852
rect 212040 79840 212046 79892
rect 102042 79772 102048 79824
rect 102100 79812 102106 79824
rect 174538 79812 174544 79824
rect 102100 79784 174544 79812
rect 102100 79772 102106 79784
rect 174538 79772 174544 79784
rect 174596 79772 174602 79824
rect 99190 79704 99196 79756
rect 99248 79744 99254 79756
rect 170398 79744 170404 79756
rect 99248 79716 170404 79744
rect 99248 79704 99254 79716
rect 170398 79704 170404 79716
rect 170456 79704 170462 79756
rect 211798 79296 211804 79348
rect 211856 79336 211862 79348
rect 307294 79336 307300 79348
rect 211856 79308 307300 79336
rect 211856 79296 211862 79308
rect 307294 79296 307300 79308
rect 307352 79296 307358 79348
rect 309686 79296 309692 79348
rect 309744 79336 309750 79348
rect 328454 79336 328460 79348
rect 309744 79308 328460 79336
rect 309744 79296 309750 79308
rect 328454 79296 328460 79308
rect 328512 79296 328518 79348
rect 97902 78616 97908 78668
rect 97960 78656 97966 78668
rect 188430 78656 188436 78668
rect 97960 78628 188436 78656
rect 97960 78616 97966 78628
rect 188430 78616 188436 78628
rect 188488 78616 188494 78668
rect 125502 78548 125508 78600
rect 125560 78588 125566 78600
rect 211890 78588 211896 78600
rect 125560 78560 211896 78588
rect 125560 78548 125566 78560
rect 211890 78548 211896 78560
rect 211948 78548 211954 78600
rect 125410 78480 125416 78532
rect 125468 78520 125474 78532
rect 206278 78520 206284 78532
rect 125468 78492 206284 78520
rect 125468 78480 125474 78492
rect 206278 78480 206284 78492
rect 206336 78480 206342 78532
rect 100018 77188 100024 77240
rect 100076 77228 100082 77240
rect 214558 77228 214564 77240
rect 100076 77200 214564 77228
rect 100076 77188 100082 77200
rect 214558 77188 214564 77200
rect 214616 77188 214622 77240
rect 93762 77120 93768 77172
rect 93820 77160 93826 77172
rect 167730 77160 167736 77172
rect 93820 77132 167736 77160
rect 93820 77120 93826 77132
rect 167730 77120 167736 77132
rect 167788 77120 167794 77172
rect 128998 77052 129004 77104
rect 129056 77092 129062 77104
rect 196802 77092 196808 77104
rect 129056 77064 196808 77092
rect 129056 77052 129062 77064
rect 196802 77052 196808 77064
rect 196860 77052 196866 77104
rect 184934 76576 184940 76628
rect 184992 76616 184998 76628
rect 315298 76616 315304 76628
rect 184992 76588 315304 76616
rect 184992 76576 184998 76588
rect 315298 76576 315304 76588
rect 315356 76576 315362 76628
rect 73154 76508 73160 76560
rect 73212 76548 73218 76560
rect 296162 76548 296168 76560
rect 73212 76520 296168 76548
rect 73212 76508 73218 76520
rect 296162 76508 296168 76520
rect 296220 76508 296226 76560
rect 63402 75828 63408 75880
rect 63460 75868 63466 75880
rect 191190 75868 191196 75880
rect 63460 75840 191196 75868
rect 63460 75828 63466 75840
rect 191190 75828 191196 75840
rect 191248 75828 191254 75880
rect 107562 75760 107568 75812
rect 107620 75800 107626 75812
rect 182910 75800 182916 75812
rect 107620 75772 182916 75800
rect 107620 75760 107626 75772
rect 182910 75760 182916 75772
rect 182968 75760 182974 75812
rect 77294 75216 77300 75268
rect 77352 75256 77358 75268
rect 270034 75256 270040 75268
rect 77352 75228 270040 75256
rect 77352 75216 77358 75228
rect 270034 75216 270040 75228
rect 270092 75216 270098 75268
rect 103514 75148 103520 75200
rect 103572 75188 103578 75200
rect 303154 75188 303160 75200
rect 103572 75160 303160 75188
rect 103572 75148 103578 75160
rect 303154 75148 303160 75160
rect 303212 75148 303218 75200
rect 91002 74468 91008 74520
rect 91060 74508 91066 74520
rect 194042 74508 194048 74520
rect 91060 74480 194048 74508
rect 91060 74468 91066 74480
rect 194042 74468 194048 74480
rect 194100 74468 194106 74520
rect 81434 73856 81440 73908
rect 81492 73896 81498 73908
rect 294690 73896 294696 73908
rect 81492 73868 294696 73896
rect 81492 73856 81498 73868
rect 294690 73856 294696 73868
rect 294748 73856 294754 73908
rect 46934 73788 46940 73840
rect 46992 73828 46998 73840
rect 274174 73828 274180 73840
rect 46992 73800 274180 73828
rect 46992 73788 46998 73800
rect 274174 73788 274180 73800
rect 274232 73788 274238 73840
rect 85482 73108 85488 73160
rect 85540 73148 85546 73160
rect 206462 73148 206468 73160
rect 85540 73120 206468 73148
rect 85540 73108 85546 73120
rect 206462 73108 206468 73120
rect 206520 73108 206526 73160
rect 418798 73108 418804 73160
rect 418856 73148 418862 73160
rect 580166 73148 580172 73160
rect 418856 73120 580172 73148
rect 418856 73108 418862 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 111058 73040 111064 73092
rect 111116 73080 111122 73092
rect 198182 73080 198188 73092
rect 111116 73052 198188 73080
rect 111116 73040 111122 73052
rect 198182 73040 198188 73052
rect 198240 73040 198246 73092
rect 85574 72428 85580 72480
rect 85632 72468 85638 72480
rect 289354 72468 289360 72480
rect 85632 72440 289360 72468
rect 85632 72428 85638 72440
rect 289354 72428 289360 72440
rect 289412 72428 289418 72480
rect 88334 71068 88340 71120
rect 88392 71108 88398 71120
rect 304258 71108 304264 71120
rect 88392 71080 304264 71108
rect 88392 71068 88398 71080
rect 304258 71068 304264 71080
rect 304316 71068 304322 71120
rect 64874 71000 64880 71052
rect 64932 71040 64938 71052
rect 293494 71040 293500 71052
rect 64932 71012 293500 71040
rect 64932 71000 64938 71012
rect 293494 71000 293500 71012
rect 293552 71000 293558 71052
rect 92474 69708 92480 69760
rect 92532 69748 92538 69760
rect 297450 69748 297456 69760
rect 92532 69720 297456 69748
rect 92532 69708 92538 69720
rect 297450 69708 297456 69720
rect 297508 69708 297514 69760
rect 53834 69640 53840 69692
rect 53892 69680 53898 69692
rect 304534 69680 304540 69692
rect 53892 69652 304540 69680
rect 53892 69640 53898 69652
rect 304534 69640 304540 69652
rect 304592 69640 304598 69692
rect 95234 68348 95240 68400
rect 95292 68388 95298 68400
rect 290550 68388 290556 68400
rect 95292 68360 290556 68388
rect 95292 68348 95298 68360
rect 290550 68348 290556 68360
rect 290608 68348 290614 68400
rect 57974 68280 57980 68332
rect 58032 68320 58038 68332
rect 296254 68320 296260 68332
rect 58032 68292 296260 68320
rect 58032 68280 58038 68292
rect 296254 68280 296260 68292
rect 296312 68280 296318 68332
rect 99374 66920 99380 66972
rect 99432 66960 99438 66972
rect 282362 66960 282368 66972
rect 99432 66932 282368 66960
rect 99432 66920 99438 66932
rect 282362 66920 282368 66932
rect 282420 66920 282426 66972
rect 69014 66852 69020 66904
rect 69072 66892 69078 66904
rect 305914 66892 305920 66904
rect 69072 66864 305920 66892
rect 69072 66852 69078 66864
rect 305914 66852 305920 66864
rect 305972 66852 305978 66904
rect 177942 65628 177948 65680
rect 178000 65668 178006 65680
rect 282362 65668 282368 65680
rect 178000 65640 282368 65668
rect 178000 65628 178006 65640
rect 282362 65628 282368 65640
rect 282420 65628 282426 65680
rect 106274 65560 106280 65612
rect 106332 65600 106338 65612
rect 258810 65600 258816 65612
rect 106332 65572 258816 65600
rect 106332 65560 106338 65572
rect 258810 65560 258816 65572
rect 258868 65560 258874 65612
rect 71774 65492 71780 65544
rect 71832 65532 71838 65544
rect 304442 65532 304448 65544
rect 71832 65504 304448 65532
rect 71832 65492 71838 65504
rect 304442 65492 304448 65504
rect 304500 65492 304506 65544
rect 110414 64200 110420 64252
rect 110472 64240 110478 64252
rect 280890 64240 280896 64252
rect 110472 64212 280896 64240
rect 110472 64200 110478 64212
rect 280890 64200 280896 64212
rect 280948 64200 280954 64252
rect 24854 64132 24860 64184
rect 24912 64172 24918 64184
rect 307202 64172 307208 64184
rect 24912 64144 307208 64172
rect 24912 64132 24918 64144
rect 307202 64132 307208 64144
rect 307260 64132 307266 64184
rect 82814 62772 82820 62824
rect 82872 62812 82878 62824
rect 300210 62812 300216 62824
rect 82872 62784 300216 62812
rect 82872 62772 82878 62784
rect 300210 62772 300216 62784
rect 300268 62772 300274 62824
rect 114554 61412 114560 61464
rect 114612 61452 114618 61464
rect 283742 61452 283748 61464
rect 114612 61424 283748 61452
rect 114612 61412 114618 61424
rect 283742 61412 283748 61424
rect 283800 61412 283806 61464
rect 13814 61344 13820 61396
rect 13872 61384 13878 61396
rect 271322 61384 271328 61396
rect 13872 61356 271328 61384
rect 13872 61344 13878 61356
rect 271322 61344 271328 61356
rect 271380 61344 271386 61396
rect 353938 60664 353944 60716
rect 353996 60704 354002 60716
rect 580166 60704 580172 60716
rect 353996 60676 580172 60704
rect 353996 60664 354002 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 74534 60052 74540 60104
rect 74592 60092 74598 60104
rect 282270 60092 282276 60104
rect 74592 60064 282276 60092
rect 74592 60052 74598 60064
rect 282270 60052 282276 60064
rect 282328 60052 282334 60104
rect 89714 59984 89720 60036
rect 89772 60024 89778 60036
rect 301774 60024 301780 60036
rect 89772 59996 301780 60024
rect 89772 59984 89778 59996
rect 301774 59984 301780 59996
rect 301832 59984 301838 60036
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 31018 59344 31024 59356
rect 3108 59316 31024 59344
rect 3108 59304 3114 59316
rect 31018 59304 31024 59316
rect 31076 59304 31082 59356
rect 93854 58692 93860 58744
rect 93912 58732 93918 58744
rect 305822 58732 305828 58744
rect 93912 58704 305828 58732
rect 93912 58692 93918 58704
rect 305822 58692 305828 58704
rect 305880 58692 305886 58744
rect 70394 58624 70400 58676
rect 70452 58664 70458 58676
rect 302970 58664 302976 58676
rect 70452 58636 302976 58664
rect 70452 58624 70458 58636
rect 302970 58624 302976 58636
rect 303028 58624 303034 58676
rect 113174 57332 113180 57384
rect 113232 57372 113238 57384
rect 287882 57372 287888 57384
rect 113232 57344 287888 57372
rect 113232 57332 113238 57344
rect 287882 57332 287888 57344
rect 287940 57332 287946 57384
rect 96614 57264 96620 57316
rect 96672 57304 96678 57316
rect 296070 57304 296076 57316
rect 96672 57276 296076 57304
rect 96672 57264 96678 57276
rect 296070 57264 296076 57276
rect 296128 57264 296134 57316
rect 63494 57196 63500 57248
rect 63552 57236 63558 57248
rect 266998 57236 267004 57248
rect 63552 57208 267004 57236
rect 63552 57196 63558 57208
rect 266998 57196 267004 57208
rect 267056 57196 267062 57248
rect 100754 55836 100760 55888
rect 100812 55876 100818 55888
rect 272518 55876 272524 55888
rect 100812 55848 272524 55876
rect 100812 55836 100818 55848
rect 272518 55836 272524 55848
rect 272576 55836 272582 55888
rect 110506 54544 110512 54596
rect 110564 54584 110570 54596
rect 300118 54584 300124 54596
rect 110564 54556 300124 54584
rect 110564 54544 110570 54556
rect 300118 54544 300124 54556
rect 300176 54544 300182 54596
rect 44174 54476 44180 54528
rect 44232 54516 44238 54528
rect 285030 54516 285036 54528
rect 44232 54488 285036 54516
rect 44232 54476 44238 54488
rect 285030 54476 285036 54488
rect 285088 54476 285094 54528
rect 37274 53116 37280 53168
rect 37332 53156 37338 53168
rect 253290 53156 253296 53168
rect 37332 53128 253296 53156
rect 37332 53116 37338 53128
rect 253290 53116 253296 53128
rect 253348 53116 253354 53168
rect 44266 53048 44272 53100
rect 44324 53088 44330 53100
rect 299014 53088 299020 53100
rect 44324 53060 299020 53088
rect 44324 53048 44330 53060
rect 299014 53048 299020 53060
rect 299072 53048 299078 53100
rect 117314 51824 117320 51876
rect 117372 51864 117378 51876
rect 261570 51864 261576 51876
rect 117372 51836 261576 51864
rect 117372 51824 117378 51836
rect 261570 51824 261576 51836
rect 261628 51824 261634 51876
rect 179230 51756 179236 51808
rect 179288 51796 179294 51808
rect 332594 51796 332600 51808
rect 179288 51768 332600 51796
rect 179288 51756 179294 51768
rect 332594 51756 332600 51768
rect 332652 51756 332658 51808
rect 16574 51688 16580 51740
rect 16632 51728 16638 51740
rect 294782 51728 294788 51740
rect 16632 51700 294788 51728
rect 16632 51688 16638 51700
rect 294782 51688 294788 51700
rect 294840 51688 294846 51740
rect 121454 50396 121460 50448
rect 121512 50436 121518 50448
rect 304350 50436 304356 50448
rect 121512 50408 304356 50436
rect 121512 50396 121518 50408
rect 304350 50396 304356 50408
rect 304408 50396 304414 50448
rect 27614 50328 27620 50380
rect 27672 50368 27678 50380
rect 264330 50368 264336 50380
rect 27672 50340 264336 50368
rect 27672 50328 27678 50340
rect 264330 50328 264336 50340
rect 264388 50328 264394 50380
rect 118694 49036 118700 49088
rect 118752 49076 118758 49088
rect 303062 49076 303068 49088
rect 118752 49048 303068 49076
rect 118752 49036 118758 49048
rect 303062 49036 303068 49048
rect 303120 49036 303126 49088
rect 30374 48968 30380 49020
rect 30432 49008 30438 49020
rect 287974 49008 287980 49020
rect 30432 48980 287980 49008
rect 30432 48968 30438 48980
rect 287974 48968 287980 48980
rect 288032 48968 288038 49020
rect 120074 47608 120080 47660
rect 120132 47648 120138 47660
rect 250438 47648 250444 47660
rect 120132 47620 250444 47648
rect 120132 47608 120138 47620
rect 250438 47608 250444 47620
rect 250496 47608 250502 47660
rect 20714 47540 20720 47592
rect 20772 47580 20778 47592
rect 291838 47580 291844 47592
rect 20772 47552 291844 47580
rect 20772 47540 20778 47552
rect 291838 47540 291844 47552
rect 291896 47540 291902 47592
rect 124214 46248 124220 46300
rect 124272 46288 124278 46300
rect 286318 46288 286324 46300
rect 124272 46260 286324 46288
rect 124272 46248 124278 46260
rect 286318 46248 286324 46260
rect 286376 46248 286382 46300
rect 26234 46180 26240 46232
rect 26292 46220 26298 46232
rect 260190 46220 260196 46232
rect 26292 46192 260196 46220
rect 26292 46180 26298 46192
rect 260190 46180 260196 46192
rect 260248 46180 260254 46232
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 18598 45540 18604 45552
rect 3476 45512 18604 45540
rect 3476 45500 3482 45512
rect 18598 45500 18604 45512
rect 18656 45500 18662 45552
rect 38654 44820 38660 44872
rect 38712 44860 38718 44872
rect 276658 44860 276664 44872
rect 38712 44832 276664 44860
rect 38712 44820 38718 44832
rect 276658 44820 276664 44832
rect 276716 44820 276722 44872
rect 31754 43460 31760 43512
rect 31812 43500 31818 43512
rect 275370 43500 275376 43512
rect 31812 43472 275376 43500
rect 31812 43460 31818 43472
rect 275370 43460 275376 43472
rect 275428 43460 275434 43512
rect 33134 43392 33140 43444
rect 33192 43432 33198 43444
rect 297542 43432 297548 43444
rect 33192 43404 297548 43432
rect 33192 43392 33198 43404
rect 297542 43392 297548 43404
rect 297600 43392 297606 43444
rect 107654 42100 107660 42152
rect 107712 42140 107718 42152
rect 295978 42140 295984 42152
rect 107712 42112 295984 42140
rect 107712 42100 107718 42112
rect 295978 42100 295984 42112
rect 296036 42100 296042 42152
rect 41414 42032 41420 42084
rect 41472 42072 41478 42084
rect 307018 42072 307024 42084
rect 41472 42044 307024 42072
rect 41472 42032 41478 42044
rect 307018 42032 307024 42044
rect 307076 42032 307082 42084
rect 35894 40740 35900 40792
rect 35952 40780 35958 40792
rect 297358 40780 297364 40792
rect 35952 40752 297364 40780
rect 35952 40740 35958 40752
rect 297358 40740 297364 40752
rect 297416 40740 297422 40792
rect 2774 40672 2780 40724
rect 2832 40712 2838 40724
rect 271138 40712 271144 40724
rect 2832 40684 271144 40712
rect 2832 40672 2838 40684
rect 271138 40672 271144 40684
rect 271196 40672 271202 40724
rect 42794 39380 42800 39432
rect 42852 39420 42858 39432
rect 283650 39420 283656 39432
rect 42852 39392 283656 39420
rect 42852 39380 42858 39392
rect 283650 39380 283656 39392
rect 283708 39380 283714 39432
rect 35986 39312 35992 39364
rect 36044 39352 36050 39364
rect 305730 39352 305736 39364
rect 36044 39324 305736 39352
rect 36044 39312 36050 39324
rect 305730 39312 305736 39324
rect 305788 39312 305794 39364
rect 78674 37952 78680 38004
rect 78732 37992 78738 38004
rect 298922 37992 298928 38004
rect 78732 37964 298928 37992
rect 78732 37952 78738 37964
rect 298922 37952 298928 37964
rect 298980 37952 298986 38004
rect 19334 37884 19340 37936
rect 19392 37924 19398 37936
rect 269850 37924 269856 37936
rect 19392 37896 269856 37924
rect 19392 37884 19398 37896
rect 269850 37884 269856 37896
rect 269908 37884 269914 37936
rect 60734 36592 60740 36644
rect 60792 36632 60798 36644
rect 305638 36632 305644 36644
rect 60792 36604 305644 36632
rect 60792 36592 60798 36604
rect 305638 36592 305644 36604
rect 305696 36592 305702 36644
rect 23474 36524 23480 36576
rect 23532 36564 23538 36576
rect 279510 36564 279516 36576
rect 23532 36536 279516 36564
rect 23532 36524 23538 36536
rect 279510 36524 279516 36536
rect 279568 36524 279574 36576
rect 35802 35844 35808 35896
rect 35860 35884 35866 35896
rect 249150 35884 249156 35896
rect 35860 35856 249156 35884
rect 35860 35844 35866 35856
rect 249150 35844 249156 35856
rect 249208 35844 249214 35896
rect 67634 35164 67640 35216
rect 67692 35204 67698 35216
rect 293218 35204 293224 35216
rect 67692 35176 293224 35204
rect 67692 35164 67698 35176
rect 293218 35164 293224 35176
rect 293276 35164 293282 35216
rect 35158 34484 35164 34536
rect 35216 34524 35222 34536
rect 35802 34524 35808 34536
rect 35216 34496 35808 34524
rect 35216 34484 35222 34496
rect 35802 34484 35808 34496
rect 35860 34484 35866 34536
rect 180794 33940 180800 33992
rect 180852 33980 180858 33992
rect 261570 33980 261576 33992
rect 180852 33952 261576 33980
rect 180852 33940 180858 33952
rect 261570 33940 261576 33952
rect 261628 33940 261634 33992
rect 201494 33872 201500 33924
rect 201552 33912 201558 33924
rect 343634 33912 343640 33924
rect 201552 33884 343640 33912
rect 201552 33872 201558 33884
rect 343634 33872 343640 33884
rect 343692 33872 343698 33924
rect 93946 33804 93952 33856
rect 94004 33844 94010 33856
rect 278222 33844 278228 33856
rect 94004 33816 278228 33844
rect 94004 33804 94010 33816
rect 278222 33804 278228 33816
rect 278280 33804 278286 33856
rect 4154 33736 4160 33788
rect 4212 33776 4218 33788
rect 251818 33776 251824 33788
rect 4212 33748 251824 33776
rect 4212 33736 4218 33748
rect 251818 33736 251824 33748
rect 251876 33736 251882 33788
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 46198 33096 46204 33108
rect 3568 33068 46204 33096
rect 3568 33056 3574 33068
rect 46198 33056 46204 33068
rect 46256 33056 46262 33108
rect 189718 32444 189724 32496
rect 189776 32484 189782 32496
rect 259546 32484 259552 32496
rect 189776 32456 259552 32484
rect 189776 32444 189782 32456
rect 259546 32444 259552 32456
rect 259604 32444 259610 32496
rect 111794 32376 111800 32428
rect 111852 32416 111858 32428
rect 301498 32416 301504 32428
rect 111852 32388 301504 32416
rect 111852 32376 111858 32388
rect 301498 32376 301504 32388
rect 301556 32376 301562 32428
rect 8294 31016 8300 31068
rect 8352 31056 8358 31068
rect 293310 31056 293316 31068
rect 8352 31028 293316 31056
rect 8352 31016 8358 31028
rect 293310 31016 293316 31028
rect 293368 31016 293374 31068
rect 200114 29724 200120 29776
rect 200172 29764 200178 29776
rect 311894 29764 311900 29776
rect 200172 29736 311900 29764
rect 200172 29724 200178 29736
rect 311894 29724 311900 29736
rect 311952 29724 311958 29776
rect 102134 29656 102140 29708
rect 102192 29696 102198 29708
rect 275278 29696 275284 29708
rect 102192 29668 275284 29696
rect 102192 29656 102198 29668
rect 275278 29656 275284 29668
rect 275336 29656 275342 29708
rect 15194 29588 15200 29640
rect 15252 29628 15258 29640
rect 253198 29628 253204 29640
rect 15252 29600 253204 29628
rect 15252 29588 15258 29600
rect 253198 29588 253204 29600
rect 253256 29588 253262 29640
rect 179506 28364 179512 28416
rect 179564 28404 179570 28416
rect 293954 28404 293960 28416
rect 179564 28376 293960 28404
rect 179564 28364 179570 28376
rect 293954 28364 293960 28376
rect 294012 28364 294018 28416
rect 84194 28296 84200 28348
rect 84252 28336 84258 28348
rect 302878 28336 302884 28348
rect 84252 28308 302884 28336
rect 84252 28296 84258 28308
rect 302878 28296 302884 28308
rect 302936 28296 302942 28348
rect 17954 28228 17960 28280
rect 18012 28268 18018 28280
rect 260098 28268 260104 28280
rect 18012 28240 260104 28268
rect 18012 28228 18018 28240
rect 260098 28228 260104 28240
rect 260156 28228 260162 28280
rect 176470 27004 176476 27056
rect 176528 27044 176534 27056
rect 296714 27044 296720 27056
rect 176528 27016 296720 27044
rect 176528 27004 176534 27016
rect 296714 27004 296720 27016
rect 296772 27004 296778 27056
rect 55214 26936 55220 26988
rect 55272 26976 55278 26988
rect 301682 26976 301688 26988
rect 55272 26948 301688 26976
rect 55272 26936 55278 26948
rect 301682 26936 301688 26948
rect 301740 26936 301746 26988
rect 2866 26868 2872 26920
rect 2924 26908 2930 26920
rect 250530 26908 250536 26920
rect 2924 26880 250536 26908
rect 2924 26868 2930 26880
rect 250530 26868 250536 26880
rect 250588 26868 250594 26920
rect 28994 25508 29000 25560
rect 29052 25548 29058 25560
rect 254578 25548 254584 25560
rect 29052 25520 254584 25548
rect 29052 25508 29058 25520
rect 254578 25508 254584 25520
rect 254636 25508 254642 25560
rect 187694 24284 187700 24336
rect 187752 24324 187758 24336
rect 254578 24324 254584 24336
rect 187752 24296 254584 24324
rect 187752 24284 187758 24296
rect 254578 24284 254584 24296
rect 254636 24284 254642 24336
rect 208394 24216 208400 24268
rect 208452 24256 208458 24268
rect 324406 24256 324412 24268
rect 208452 24228 324412 24256
rect 208452 24216 208458 24228
rect 324406 24216 324412 24228
rect 324464 24216 324470 24268
rect 86954 24148 86960 24200
rect 87012 24188 87018 24200
rect 284938 24188 284944 24200
rect 87012 24160 284944 24188
rect 87012 24148 87018 24160
rect 284938 24148 284944 24160
rect 284996 24148 285002 24200
rect 52454 24080 52460 24132
rect 52512 24120 52518 24132
rect 268470 24120 268476 24132
rect 52512 24092 268476 24120
rect 52512 24080 52518 24092
rect 268470 24080 268476 24092
rect 268528 24080 268534 24132
rect 69106 22788 69112 22840
rect 69164 22828 69170 22840
rect 294598 22828 294604 22840
rect 69164 22800 294604 22828
rect 69164 22788 69170 22800
rect 294598 22788 294604 22800
rect 294656 22788 294662 22840
rect 40034 22720 40040 22772
rect 40092 22760 40098 22772
rect 271230 22760 271236 22772
rect 40092 22732 271236 22760
rect 40092 22720 40098 22732
rect 271230 22720 271236 22732
rect 271288 22720 271294 22772
rect 183554 21496 183560 21548
rect 183612 21536 183618 21548
rect 349338 21536 349344 21548
rect 183612 21508 349344 21536
rect 183612 21496 183618 21508
rect 349338 21496 349344 21508
rect 349396 21496 349402 21548
rect 91094 21428 91100 21480
rect 91152 21468 91158 21480
rect 291930 21468 291936 21480
rect 91152 21440 291936 21468
rect 91152 21428 91158 21440
rect 291930 21428 291936 21440
rect 291988 21428 291994 21480
rect 19426 21360 19432 21412
rect 19484 21400 19490 21412
rect 261662 21400 261668 21412
rect 19484 21372 261668 21400
rect 19484 21360 19490 21372
rect 261662 21360 261668 21372
rect 261720 21360 261726 21412
rect 378778 20612 378784 20664
rect 378836 20652 378842 20664
rect 579982 20652 579988 20664
rect 378836 20624 579988 20652
rect 378836 20612 378842 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 102226 20000 102232 20052
rect 102284 20040 102290 20052
rect 249058 20040 249064 20052
rect 102284 20012 249064 20040
rect 102284 20000 102290 20012
rect 249058 20000 249064 20012
rect 249116 20000 249122 20052
rect 80054 19932 80060 19984
rect 80112 19972 80118 19984
rect 280798 19972 280804 19984
rect 80112 19944 280804 19972
rect 80112 19932 80118 19944
rect 280798 19932 280804 19944
rect 280856 19932 280862 19984
rect 3418 19456 3424 19508
rect 3476 19496 3482 19508
rect 7558 19496 7564 19508
rect 3476 19468 7564 19496
rect 3476 19456 3482 19468
rect 7558 19456 7564 19468
rect 7616 19456 7622 19508
rect 75914 18572 75920 18624
rect 75972 18612 75978 18624
rect 261478 18612 261484 18624
rect 75972 18584 261484 18612
rect 75972 18572 75978 18584
rect 261478 18572 261484 18584
rect 261536 18572 261542 18624
rect 193214 17280 193220 17332
rect 193272 17320 193278 17332
rect 247034 17320 247040 17332
rect 193272 17292 247040 17320
rect 193272 17280 193278 17292
rect 247034 17280 247040 17292
rect 247092 17280 247098 17332
rect 128354 17212 128360 17264
rect 128412 17252 128418 17264
rect 215938 17252 215944 17264
rect 128412 17224 215944 17252
rect 128412 17212 128418 17224
rect 215938 17212 215944 17224
rect 215996 17212 216002 17264
rect 217962 17212 217968 17264
rect 218020 17252 218026 17264
rect 248414 17252 248420 17264
rect 218020 17224 248420 17252
rect 218020 17212 218026 17224
rect 248414 17212 248420 17224
rect 248472 17212 248478 17264
rect 192478 15988 192484 16040
rect 192536 16028 192542 16040
rect 273254 16028 273260 16040
rect 192536 16000 273260 16028
rect 192536 15988 192542 16000
rect 273254 15988 273260 16000
rect 273312 15988 273318 16040
rect 105722 15920 105728 15972
rect 105780 15960 105786 15972
rect 289170 15960 289176 15972
rect 105780 15932 289176 15960
rect 105780 15920 105786 15932
rect 289170 15920 289176 15932
rect 289228 15920 289234 15972
rect 11882 15852 11888 15904
rect 11940 15892 11946 15904
rect 258718 15892 258724 15904
rect 11940 15864 258724 15892
rect 11940 15852 11946 15864
rect 258718 15852 258724 15864
rect 258776 15852 258782 15904
rect 212534 14560 212540 14612
rect 212592 14600 212598 14612
rect 327994 14600 328000 14612
rect 212592 14572 328000 14600
rect 212592 14560 212598 14572
rect 327994 14560 328000 14572
rect 328052 14560 328058 14612
rect 77386 14492 77392 14544
rect 77444 14532 77450 14544
rect 273990 14532 273996 14544
rect 77444 14504 273996 14532
rect 77444 14492 77450 14504
rect 273990 14492 273996 14504
rect 274048 14492 274054 14544
rect 34514 14424 34520 14476
rect 34572 14464 34578 14476
rect 298830 14464 298836 14476
rect 34572 14436 298836 14464
rect 34572 14424 34578 14436
rect 298830 14424 298836 14436
rect 298888 14424 298894 14476
rect 173802 13132 173808 13184
rect 173860 13172 173866 13184
rect 301498 13172 301504 13184
rect 173860 13144 301504 13172
rect 173860 13132 173866 13144
rect 301498 13132 301504 13144
rect 301556 13132 301562 13184
rect 109034 13064 109040 13116
rect 109092 13104 109098 13116
rect 265618 13104 265624 13116
rect 109092 13076 265624 13104
rect 109092 13064 109098 13076
rect 265618 13064 265624 13076
rect 265676 13064 265682 13116
rect 211062 11908 211068 11960
rect 211120 11948 211126 11960
rect 252370 11948 252376 11960
rect 211120 11920 252376 11948
rect 211120 11908 211126 11920
rect 252370 11908 252376 11920
rect 252428 11908 252434 11960
rect 176562 11840 176568 11892
rect 176620 11880 176626 11892
rect 262490 11880 262496 11892
rect 176620 11852 262496 11880
rect 176620 11840 176626 11852
rect 262490 11840 262496 11852
rect 262548 11840 262554 11892
rect 51074 11772 51080 11824
rect 51132 11812 51138 11824
rect 228358 11812 228364 11824
rect 51132 11784 228364 11812
rect 51132 11772 51138 11784
rect 228358 11772 228364 11784
rect 228416 11772 228422 11824
rect 98178 11704 98184 11756
rect 98236 11744 98242 11756
rect 283558 11744 283564 11756
rect 98236 11716 283564 11744
rect 98236 11704 98242 11716
rect 283558 11704 283564 11716
rect 283616 11704 283622 11756
rect 106 10956 112 11008
rect 164 10996 170 11008
rect 1302 10996 1308 11008
rect 164 10968 1308 10996
rect 164 10956 170 10968
rect 1302 10956 1308 10968
rect 1360 10996 1366 11008
rect 251174 10996 251180 11008
rect 1360 10968 251180 10996
rect 1360 10956 1366 10968
rect 251174 10956 251180 10968
rect 251232 10956 251238 11008
rect 179414 10344 179420 10396
rect 179472 10384 179478 10396
rect 299658 10384 299664 10396
rect 179472 10356 299664 10384
rect 179472 10344 179478 10356
rect 299658 10344 299664 10356
rect 299716 10344 299722 10396
rect 28442 10276 28448 10328
rect 28500 10316 28506 10328
rect 278130 10316 278136 10328
rect 28500 10288 278136 10316
rect 28500 10276 28506 10288
rect 278130 10276 278136 10288
rect 278188 10276 278194 10328
rect 197998 9052 198004 9104
rect 198056 9092 198062 9104
rect 287790 9092 287796 9104
rect 198056 9064 287796 9092
rect 198056 9052 198062 9064
rect 287790 9052 287796 9064
rect 287848 9052 287854 9104
rect 46658 8984 46664 9036
rect 46716 9024 46722 9036
rect 273898 9024 273904 9036
rect 46716 8996 273904 9024
rect 46716 8984 46722 8996
rect 273898 8984 273904 8996
rect 273956 8984 273962 9036
rect 6454 8916 6460 8968
rect 6512 8956 6518 8968
rect 289262 8956 289268 8968
rect 6512 8928 289268 8956
rect 6512 8916 6518 8928
rect 289262 8916 289268 8928
rect 289320 8916 289326 8968
rect 308398 8916 308404 8968
rect 308456 8956 308462 8968
rect 317322 8956 317328 8968
rect 308456 8928 317328 8956
rect 308456 8916 308462 8928
rect 317322 8916 317328 8928
rect 317380 8916 317386 8968
rect 331858 8236 331864 8288
rect 331916 8276 331922 8288
rect 333882 8276 333888 8288
rect 331916 8248 333888 8276
rect 331916 8236 331922 8248
rect 333882 8236 333888 8248
rect 333940 8236 333946 8288
rect 116394 7624 116400 7676
rect 116452 7664 116458 7676
rect 287698 7664 287704 7676
rect 116452 7636 287704 7664
rect 116452 7624 116458 7636
rect 287698 7624 287704 7636
rect 287756 7624 287762 7676
rect 7650 7556 7656 7608
rect 7708 7596 7714 7608
rect 269758 7596 269764 7608
rect 7708 7568 269764 7596
rect 7708 7556 7714 7568
rect 269758 7556 269764 7568
rect 269816 7556 269822 7608
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 48958 6848 48964 6860
rect 3476 6820 48964 6848
rect 3476 6808 3482 6820
rect 48958 6808 48964 6820
rect 49016 6808 49022 6860
rect 203518 6332 203524 6384
rect 203576 6372 203582 6384
rect 266538 6372 266544 6384
rect 203576 6344 266544 6372
rect 203576 6332 203582 6344
rect 266538 6332 266544 6344
rect 266596 6332 266602 6384
rect 175182 6264 175188 6316
rect 175240 6304 175246 6316
rect 311434 6304 311440 6316
rect 175240 6276 311440 6304
rect 175240 6264 175246 6276
rect 311434 6264 311440 6276
rect 311492 6264 311498 6316
rect 123478 6196 123484 6248
rect 123536 6236 123542 6248
rect 290458 6236 290464 6248
rect 123536 6208 290464 6236
rect 123536 6196 123542 6208
rect 290458 6196 290464 6208
rect 290516 6196 290522 6248
rect 86862 6128 86868 6180
rect 86920 6168 86926 6180
rect 255958 6168 255964 6180
rect 86920 6140 255964 6168
rect 86920 6128 86926 6140
rect 255958 6128 255964 6140
rect 256016 6128 256022 6180
rect 1670 4768 1676 4820
rect 1728 4808 1734 4820
rect 35158 4808 35164 4820
rect 1728 4780 35164 4808
rect 1728 4768 1734 4780
rect 35158 4768 35164 4780
rect 35216 4768 35222 4820
rect 48958 4768 48964 4820
rect 49016 4808 49022 4820
rect 262858 4808 262864 4820
rect 49016 4780 262864 4808
rect 49016 4768 49022 4780
rect 262858 4768 262864 4780
rect 262916 4768 262922 4820
rect 309778 4768 309784 4820
rect 309836 4808 309842 4820
rect 320910 4808 320916 4820
rect 309836 4780 320916 4808
rect 309836 4768 309842 4780
rect 320910 4768 320916 4780
rect 320968 4768 320974 4820
rect 345658 4156 345664 4208
rect 345716 4196 345722 4208
rect 350442 4196 350448 4208
rect 345716 4168 350448 4196
rect 345716 4156 345722 4168
rect 350442 4156 350448 4168
rect 350500 4156 350506 4208
rect 261570 4088 261576 4140
rect 261628 4128 261634 4140
rect 268838 4128 268844 4140
rect 261628 4100 268844 4128
rect 261628 4088 261634 4100
rect 268838 4088 268844 4100
rect 268896 4088 268902 4140
rect 315298 4088 315304 4140
rect 315356 4128 315362 4140
rect 316218 4128 316224 4140
rect 315356 4100 316224 4128
rect 315356 4088 315362 4100
rect 316218 4088 316224 4100
rect 316276 4088 316282 4140
rect 348050 3952 348056 4004
rect 348108 3992 348114 4004
rect 354674 3992 354680 4004
rect 348108 3964 354680 3992
rect 348108 3952 348114 3964
rect 354674 3952 354680 3964
rect 354732 3952 354738 4004
rect 202138 3680 202144 3732
rect 202196 3720 202202 3732
rect 267734 3720 267740 3732
rect 202196 3692 267740 3720
rect 202196 3680 202202 3692
rect 267734 3680 267740 3692
rect 267792 3680 267798 3732
rect 278038 3680 278044 3732
rect 278096 3720 278102 3732
rect 278096 3692 287054 3720
rect 278096 3680 278102 3692
rect 125870 3612 125876 3664
rect 125928 3652 125934 3664
rect 173894 3652 173900 3664
rect 125928 3624 173900 3652
rect 125928 3612 125934 3624
rect 173894 3612 173900 3624
rect 173952 3612 173958 3664
rect 196618 3612 196624 3664
rect 196676 3652 196682 3664
rect 281902 3652 281908 3664
rect 196676 3624 281908 3652
rect 196676 3612 196682 3624
rect 281902 3612 281908 3624
rect 281960 3612 281966 3664
rect 77294 3544 77300 3596
rect 77352 3584 77358 3596
rect 78214 3584 78220 3596
rect 77352 3556 78220 3584
rect 77352 3544 77358 3556
rect 78214 3544 78220 3556
rect 78272 3544 78278 3596
rect 119890 3544 119896 3596
rect 119948 3584 119954 3596
rect 224218 3584 224224 3596
rect 119948 3556 224224 3584
rect 119948 3544 119954 3556
rect 224218 3544 224224 3556
rect 224276 3544 224282 3596
rect 254578 3544 254584 3596
rect 254636 3584 254642 3596
rect 261754 3584 261760 3596
rect 254636 3556 261760 3584
rect 254636 3544 254642 3556
rect 261754 3544 261760 3556
rect 261812 3544 261818 3596
rect 282178 3544 282184 3596
rect 282236 3584 282242 3596
rect 287026 3584 287054 3692
rect 288986 3584 288992 3596
rect 282236 3556 284616 3584
rect 287026 3556 288992 3584
rect 282236 3544 282242 3556
rect 44174 3476 44180 3528
rect 44232 3516 44238 3528
rect 45094 3516 45100 3528
rect 44232 3488 45100 3516
rect 44232 3476 44238 3488
rect 45094 3476 45100 3488
rect 45152 3476 45158 3528
rect 60826 3476 60832 3528
rect 60884 3516 60890 3528
rect 203610 3516 203616 3528
rect 60884 3488 203616 3516
rect 60884 3476 60890 3488
rect 203610 3476 203616 3488
rect 203668 3476 203674 3528
rect 210418 3476 210424 3528
rect 210476 3516 210482 3528
rect 210476 3488 242848 3516
rect 210476 3476 210482 3488
rect 11146 3408 11152 3460
rect 11204 3448 11210 3460
rect 211798 3448 211804 3460
rect 11204 3420 211804 3448
rect 11204 3408 11210 3420
rect 211798 3408 211804 3420
rect 211856 3408 211862 3460
rect 216030 3408 216036 3460
rect 216088 3448 216094 3460
rect 240502 3448 240508 3460
rect 216088 3420 240508 3448
rect 216088 3408 216094 3420
rect 240502 3408 240508 3420
rect 240560 3408 240566 3460
rect 242820 3448 242848 3488
rect 242894 3476 242900 3528
rect 242952 3516 242958 3528
rect 244090 3516 244096 3528
rect 242952 3488 244096 3516
rect 242952 3476 242958 3488
rect 244090 3476 244096 3488
rect 244148 3476 244154 3528
rect 246942 3476 246948 3528
rect 247000 3516 247006 3528
rect 259454 3516 259460 3528
rect 247000 3488 259460 3516
rect 247000 3476 247006 3488
rect 259454 3476 259460 3488
rect 259512 3476 259518 3528
rect 268378 3476 268384 3528
rect 268436 3516 268442 3528
rect 278314 3516 278320 3528
rect 268436 3488 278320 3516
rect 268436 3476 268442 3488
rect 278314 3476 278320 3488
rect 278372 3476 278378 3528
rect 282362 3476 282368 3528
rect 282420 3516 282426 3528
rect 284294 3516 284300 3528
rect 282420 3488 284300 3516
rect 282420 3476 282426 3488
rect 284294 3476 284300 3488
rect 284352 3476 284358 3528
rect 284588 3516 284616 3556
rect 288986 3544 288992 3556
rect 289044 3544 289050 3596
rect 289078 3544 289084 3596
rect 289136 3584 289142 3596
rect 298462 3584 298468 3596
rect 289136 3556 298468 3584
rect 289136 3544 289142 3556
rect 298462 3544 298468 3556
rect 298520 3544 298526 3596
rect 319438 3544 319444 3596
rect 319496 3584 319502 3596
rect 319496 3556 319852 3584
rect 319496 3544 319502 3556
rect 292574 3516 292580 3528
rect 284588 3488 292580 3516
rect 292574 3476 292580 3488
rect 292632 3476 292638 3528
rect 299474 3476 299480 3528
rect 299532 3516 299538 3528
rect 300762 3516 300768 3528
rect 299532 3488 300768 3516
rect 299532 3476 299538 3488
rect 300762 3476 300768 3488
rect 300820 3476 300826 3528
rect 301590 3476 301596 3528
rect 301648 3516 301654 3528
rect 319714 3516 319720 3528
rect 301648 3488 319720 3516
rect 301648 3476 301654 3488
rect 319714 3476 319720 3488
rect 319772 3476 319778 3528
rect 319824 3516 319852 3556
rect 324406 3544 324412 3596
rect 324464 3584 324470 3596
rect 325602 3584 325608 3596
rect 324464 3556 325608 3584
rect 324464 3544 324470 3556
rect 325602 3544 325608 3556
rect 325660 3544 325666 3596
rect 338666 3544 338672 3596
rect 338724 3584 338730 3596
rect 349154 3584 349160 3596
rect 338724 3556 349160 3584
rect 338724 3544 338730 3556
rect 349154 3544 349160 3556
rect 349212 3544 349218 3596
rect 349338 3544 349344 3596
rect 349396 3544 349402 3596
rect 345750 3516 345756 3528
rect 319824 3488 345756 3516
rect 345750 3476 345756 3488
rect 345808 3476 345814 3528
rect 245194 3448 245200 3460
rect 242820 3420 245200 3448
rect 245194 3408 245200 3420
rect 245252 3408 245258 3460
rect 247678 3408 247684 3460
rect 247736 3448 247742 3460
rect 254670 3448 254676 3460
rect 247736 3420 254676 3448
rect 247736 3408 247742 3420
rect 254670 3408 254676 3420
rect 254728 3408 254734 3460
rect 256602 3408 256608 3460
rect 256660 3448 256666 3460
rect 271230 3448 271236 3460
rect 256660 3420 271236 3448
rect 256660 3408 256666 3420
rect 271230 3408 271236 3420
rect 271288 3408 271294 3460
rect 279418 3408 279424 3460
rect 279476 3448 279482 3460
rect 326798 3448 326804 3460
rect 279476 3420 326804 3448
rect 279476 3408 279482 3420
rect 326798 3408 326804 3420
rect 326856 3408 326862 3460
rect 330386 3408 330392 3460
rect 330444 3448 330450 3460
rect 349356 3448 349384 3544
rect 330444 3420 349384 3448
rect 330444 3408 330450 3420
rect 356698 3408 356704 3460
rect 356756 3448 356762 3460
rect 579798 3448 579804 3460
rect 356756 3420 579804 3448
rect 356756 3408 356762 3420
rect 579798 3408 579804 3420
rect 579856 3408 579862 3460
rect 308582 3340 308588 3392
rect 308640 3380 308646 3392
rect 315022 3380 315028 3392
rect 308640 3352 315028 3380
rect 308640 3340 308646 3352
rect 315022 3340 315028 3352
rect 315080 3340 315086 3392
rect 264238 3272 264244 3324
rect 264296 3312 264302 3324
rect 270034 3312 270040 3324
rect 264296 3284 270040 3312
rect 264296 3272 264302 3284
rect 270034 3272 270040 3284
rect 270092 3272 270098 3324
rect 249978 3204 249984 3256
rect 250036 3244 250042 3256
rect 256050 3244 256056 3256
rect 250036 3216 256056 3244
rect 250036 3204 250042 3216
rect 256050 3204 256056 3216
rect 256108 3204 256114 3256
rect 269942 3000 269948 3052
rect 270000 3040 270006 3052
rect 276014 3040 276020 3052
rect 270000 3012 276020 3040
rect 270000 3000 270006 3012
rect 276014 3000 276020 3012
rect 276072 3000 276078 3052
rect 235810 2932 235816 2984
rect 235868 2972 235874 2984
rect 238018 2972 238024 2984
rect 235868 2944 238024 2972
rect 235868 2932 235874 2944
rect 238018 2932 238024 2944
rect 238076 2932 238082 2984
rect 179322 2116 179328 2168
rect 179380 2156 179386 2168
rect 306742 2156 306748 2168
rect 179380 2128 306748 2156
rect 179380 2116 179386 2128
rect 306742 2116 306748 2128
rect 306800 2116 306806 2168
rect 59630 2048 59636 2100
rect 59688 2088 59694 2100
rect 287882 2088 287888 2100
rect 59688 2060 287888 2088
rect 59688 2048 59694 2060
rect 287882 2048 287888 2060
rect 287940 2048 287946 2100
<< via1 >>
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 301504 702652 301556 702704
rect 494796 702652 494848 702704
rect 209780 702584 209832 702636
rect 462320 702584 462372 702636
rect 177948 702516 178000 702568
rect 478512 702516 478564 702568
rect 206284 702448 206336 702500
rect 559656 702448 559708 702500
rect 72976 700340 73028 700392
rect 82084 700340 82136 700392
rect 105452 700340 105504 700392
rect 193220 700340 193272 700392
rect 235172 700340 235224 700392
rect 305000 700340 305052 700392
rect 24308 700272 24360 700324
rect 43444 700272 43496 700324
rect 62764 700272 62816 700324
rect 170312 700272 170364 700324
rect 218980 700272 219032 700324
rect 310520 700272 310572 700324
rect 319444 700272 319496 700324
rect 429844 700272 429896 700324
rect 300124 699660 300176 699712
rect 306472 699660 306524 699712
rect 525064 699660 525116 699712
rect 527180 699660 527232 699712
rect 324964 698912 325016 698964
rect 397460 698912 397512 698964
rect 266360 697620 266412 697672
rect 267648 697620 267700 697672
rect 211804 697552 211856 697604
rect 348792 697552 348844 697604
rect 3424 683136 3476 683188
rect 189724 683136 189776 683188
rect 297364 683136 297416 683188
rect 580172 683136 580224 683188
rect 3516 670692 3568 670744
rect 22744 670692 22796 670744
rect 2780 656956 2832 657008
rect 4804 656956 4856 657008
rect 3424 632068 3476 632120
rect 44824 632068 44876 632120
rect 179328 630640 179380 630692
rect 579988 630640 580040 630692
rect 3148 618264 3200 618316
rect 18604 618264 18656 618316
rect 337384 616836 337436 616888
rect 580172 616836 580224 616888
rect 3424 606024 3476 606076
rect 8944 606024 8996 606076
rect 309784 590656 309836 590708
rect 580172 590656 580224 590708
rect 3332 579640 3384 579692
rect 116584 579640 116636 579692
rect 3424 565836 3476 565888
rect 21364 565836 21416 565888
rect 158628 563048 158680 563100
rect 579896 563048 579948 563100
rect 3424 553392 3476 553444
rect 17224 553392 17276 553444
rect 3424 527144 3476 527196
rect 13084 527144 13136 527196
rect 347044 524424 347096 524476
rect 580172 524424 580224 524476
rect 400864 510620 400916 510672
rect 580172 510620 580224 510672
rect 3056 474716 3108 474768
rect 202880 474716 202932 474768
rect 278044 470568 278096 470620
rect 580172 470568 580224 470620
rect 3516 462340 3568 462392
rect 111064 462340 111116 462392
rect 166908 456764 166960 456816
rect 580172 456764 580224 456816
rect 3148 448536 3200 448588
rect 39304 448536 39356 448588
rect 3516 422288 3568 422340
rect 32404 422288 32456 422340
rect 2872 409844 2924 409896
rect 53104 409844 53156 409896
rect 160836 404336 160888 404388
rect 579988 404336 580040 404388
rect 3516 397468 3568 397520
rect 58624 397468 58676 397520
rect 220084 378156 220136 378208
rect 580172 378156 580224 378208
rect 179420 377408 179472 377460
rect 266360 377408 266412 377460
rect 195888 375980 195940 376032
rect 331220 375980 331272 376032
rect 179052 374620 179104 374672
rect 580264 374620 580316 374672
rect 122748 373260 122800 373312
rect 201500 373260 201552 373312
rect 189724 371832 189776 371884
rect 198740 371832 198792 371884
rect 3516 371220 3568 371272
rect 128360 371220 128412 371272
rect 206376 371220 206428 371272
rect 327724 371220 327776 371272
rect 179144 370472 179196 370524
rect 580356 370472 580408 370524
rect 209044 369112 209096 369164
rect 220084 369112 220136 369164
rect 39304 368908 39356 368960
rect 39948 368908 40000 368960
rect 194600 368908 194652 368960
rect 195888 368908 195940 368960
rect 64696 368568 64748 368620
rect 194600 368568 194652 368620
rect 39948 368500 40000 368552
rect 295616 368500 295668 368552
rect 109040 367072 109092 367124
rect 254584 367072 254636 367124
rect 142804 365780 142856 365832
rect 276020 365780 276072 365832
rect 124864 365712 124916 365764
rect 287060 365712 287112 365764
rect 190460 364488 190512 364540
rect 315304 364488 315356 364540
rect 69204 364420 69256 364472
rect 242900 364420 242952 364472
rect 179880 364352 179932 364404
rect 580172 364352 580224 364404
rect 117964 363060 118016 363112
rect 214472 363060 214524 363112
rect 130384 362992 130436 363044
rect 295340 362992 295392 363044
rect 179236 362924 179288 362976
rect 580264 362924 580316 362976
rect 282920 362176 282972 362228
rect 295432 362176 295484 362228
rect 174728 361700 174780 361752
rect 237472 361700 237524 361752
rect 273536 361700 273588 361752
rect 278044 361700 278096 361752
rect 134524 361632 134576 361684
rect 256792 361632 256844 361684
rect 79324 361564 79376 361616
rect 245844 361564 245896 361616
rect 162768 360476 162820 360528
rect 197728 360476 197780 360528
rect 126244 360408 126296 360460
rect 201592 360408 201644 360460
rect 225420 360408 225472 360460
rect 303620 360408 303672 360460
rect 167644 360340 167696 360392
rect 279332 360340 279384 360392
rect 170404 360272 170456 360324
rect 291844 360272 291896 360324
rect 69112 360204 69164 360256
rect 220268 360204 220320 360256
rect 254400 360204 254452 360256
rect 254584 360204 254636 360256
rect 373264 360204 373316 360256
rect 144184 359048 144236 359100
rect 283380 359048 283432 359100
rect 157248 358980 157300 359032
rect 184940 358980 184992 359032
rect 282092 358912 282144 358964
rect 311900 358912 311952 358964
rect 181628 358844 181680 358896
rect 349160 358844 349212 358896
rect 101404 358776 101456 358828
rect 294144 358776 294196 358828
rect 187424 358028 187476 358080
rect 206376 358028 206428 358080
rect 269028 357824 269080 357876
rect 349252 357824 349304 357876
rect 242808 357756 242860 357808
rect 270500 357756 270552 357808
rect 174636 357688 174688 357740
rect 241520 357688 241572 357740
rect 260748 357688 260800 357740
rect 296812 357688 296864 357740
rect 179788 357620 179840 357672
rect 211804 357620 211856 357672
rect 223488 357620 223540 357672
rect 291752 357620 291804 357672
rect 148324 357552 148376 357604
rect 193220 357552 193272 357604
rect 217048 357552 217100 357604
rect 317420 357552 317472 357604
rect 3056 357484 3108 357536
rect 90364 357484 90416 357536
rect 107660 357484 107712 357536
rect 289452 357484 289504 357536
rect 290464 357484 290516 357536
rect 308404 357484 308456 357536
rect 55036 357416 55088 357468
rect 265164 357416 265216 357468
rect 287152 357416 287204 357468
rect 293316 357416 293368 357468
rect 154028 357348 154080 357400
rect 242808 357348 242860 357400
rect 68652 356668 68704 356720
rect 153200 356668 153252 356720
rect 154028 356668 154080 356720
rect 174544 356328 174596 356380
rect 208768 356328 208820 356380
rect 258908 356328 258960 356380
rect 299572 356328 299624 356380
rect 171876 356260 171928 356312
rect 273536 356260 273588 356312
rect 285956 356260 286008 356312
rect 313280 356260 313332 356312
rect 140136 356192 140188 356244
rect 247960 356192 248012 356244
rect 252468 356192 252520 356244
rect 301596 356192 301648 356244
rect 111156 356124 111208 356176
rect 295524 356124 295576 356176
rect 80060 356056 80112 356108
rect 298192 356056 298244 356108
rect 289452 355988 289504 356040
rect 294236 355988 294288 356040
rect 111064 355308 111116 355360
rect 135260 355308 135312 355360
rect 202880 355240 202932 355292
rect 203846 355240 203898 355292
rect 171784 355036 171836 355088
rect 198740 355036 198792 355088
rect 199660 355036 199712 355088
rect 169024 354968 169076 355020
rect 202880 354968 202932 355020
rect 275652 354968 275704 355020
rect 299756 354968 299808 355020
rect 175924 354900 175976 354952
rect 235080 354900 235132 354952
rect 256792 354900 256844 354952
rect 297456 354900 297508 354952
rect 97264 354832 97316 354884
rect 293040 354832 293092 354884
rect 75920 354764 75972 354816
rect 294052 354764 294104 354816
rect 135260 354696 135312 354748
rect 266636 354696 266688 354748
rect 279516 354696 279568 354748
rect 449164 354696 449216 354748
rect 84292 354016 84344 354068
rect 179788 354016 179840 354068
rect 44824 353948 44876 354000
rect 45468 353948 45520 354000
rect 176660 353948 176712 354000
rect 293316 353948 293368 354000
rect 580356 353948 580408 354000
rect 177856 353268 177908 353320
rect 179880 353268 179932 353320
rect 113180 352520 113232 352572
rect 179604 352520 179656 352572
rect 50896 351160 50948 351212
rect 174728 351160 174780 351212
rect 293132 351160 293184 351212
rect 580264 351160 580316 351212
rect 127716 347760 127768 347812
rect 176660 347760 176712 347812
rect 6920 347012 6972 347064
rect 62856 347012 62908 347064
rect 3332 345040 3384 345092
rect 25504 345040 25556 345092
rect 296168 345040 296220 345092
rect 472624 345040 472676 345092
rect 72424 344292 72476 344344
rect 174636 344292 174688 344344
rect 295340 343544 295392 343596
rect 295616 343544 295668 343596
rect 295340 342864 295392 342916
rect 300860 342728 300912 342780
rect 301504 342728 301556 342780
rect 175188 342252 175240 342304
rect 176660 342252 176712 342304
rect 124128 340892 124180 340944
rect 176660 340892 176712 340944
rect 295340 339464 295392 339516
rect 308496 339464 308548 339516
rect 90364 335996 90416 336048
rect 98644 335996 98696 336048
rect 161572 334568 161624 334620
rect 177948 334568 178000 334620
rect 104164 332596 104216 332648
rect 176660 332596 176712 332648
rect 106280 330488 106332 330540
rect 161572 330488 161624 330540
rect 374644 330488 374696 330540
rect 412640 330488 412692 330540
rect 294420 327088 294472 327140
rect 311164 327088 311216 327140
rect 130568 325660 130620 325712
rect 179512 325660 179564 325712
rect 355324 324300 355376 324352
rect 580172 324300 580224 324352
rect 173808 321580 173860 321632
rect 176660 321580 176712 321632
rect 3424 320832 3476 320884
rect 120080 320832 120132 320884
rect 295524 320152 295576 320204
rect 305644 320152 305696 320204
rect 3424 318792 3476 318844
rect 100024 318792 100076 318844
rect 295524 318792 295576 318844
rect 350540 318792 350592 318844
rect 295616 316684 295668 316736
rect 468484 316684 468536 316736
rect 166264 314644 166316 314696
rect 176660 314644 176712 314696
rect 295524 314576 295576 314628
rect 299480 314576 299532 314628
rect 25504 313896 25556 313948
rect 119620 313896 119672 313948
rect 299480 313896 299532 313948
rect 418804 313896 418856 313948
rect 116584 312740 116636 312792
rect 121460 312740 121512 312792
rect 8944 312536 8996 312588
rect 94504 312536 94556 312588
rect 302240 312536 302292 312588
rect 309784 312536 309836 312588
rect 129188 311924 129240 311976
rect 166264 311924 166316 311976
rect 138112 311856 138164 311908
rect 178960 311856 179012 311908
rect 295524 311856 295576 311908
rect 302240 311856 302292 311908
rect 4804 311108 4856 311160
rect 121552 311108 121604 311160
rect 295524 309748 295576 309800
rect 298192 309748 298244 309800
rect 471244 309748 471296 309800
rect 173164 309136 173216 309188
rect 176660 309136 176712 309188
rect 158536 307844 158588 307896
rect 176660 307844 176712 307896
rect 82176 307776 82228 307828
rect 164976 307776 165028 307828
rect 295524 307776 295576 307828
rect 303712 307776 303764 307828
rect 91100 307028 91152 307080
rect 138112 307028 138164 307080
rect 85580 306348 85632 306400
rect 140228 306348 140280 306400
rect 314660 305600 314712 305652
rect 347044 305600 347096 305652
rect 75368 305056 75420 305108
rect 147036 305056 147088 305108
rect 3240 304988 3292 305040
rect 120172 304988 120224 305040
rect 176660 304988 176712 305040
rect 295432 304988 295484 305040
rect 314660 304988 314712 305040
rect 32404 304920 32456 304972
rect 72240 304920 72292 304972
rect 82084 304240 82136 304292
rect 115848 304240 115900 304292
rect 98736 303696 98788 303748
rect 149704 303696 149756 303748
rect 94596 303628 94648 303680
rect 146944 303628 146996 303680
rect 88340 303560 88392 303612
rect 104164 303560 104216 303612
rect 104440 303560 104492 303612
rect 294236 303560 294288 303612
rect 374644 303560 374696 303612
rect 43444 302880 43496 302932
rect 84384 302880 84436 302932
rect 89720 302268 89772 302320
rect 163596 302268 163648 302320
rect 74540 302200 74592 302252
rect 162216 302200 162268 302252
rect 114744 302132 114796 302184
rect 115848 302132 115900 302184
rect 173164 302132 173216 302184
rect 100024 301452 100076 301504
rect 116584 301452 116636 301504
rect 106924 301044 106976 301096
rect 133144 301044 133196 301096
rect 103704 300976 103756 301028
rect 143080 300976 143132 301028
rect 90272 300908 90324 300960
rect 142896 300908 142948 300960
rect 7564 300840 7616 300892
rect 117964 300840 118016 300892
rect 160008 300772 160060 300824
rect 160836 300772 160888 300824
rect 39948 300092 40000 300144
rect 70952 300092 71004 300144
rect 99380 299820 99432 299872
rect 124956 299820 125008 299872
rect 92848 299752 92900 299804
rect 130476 299752 130528 299804
rect 109132 299684 109184 299736
rect 153936 299684 153988 299736
rect 85672 299616 85724 299668
rect 137284 299616 137336 299668
rect 81440 299548 81492 299600
rect 157984 299548 158036 299600
rect 66168 299480 66220 299532
rect 160008 299480 160060 299532
rect 166448 299412 166500 299464
rect 166908 299412 166960 299464
rect 176660 299412 176712 299464
rect 297456 299412 297508 299464
rect 579620 299412 579672 299464
rect 102232 298392 102284 298444
rect 145656 298392 145708 298444
rect 106740 298324 106792 298376
rect 151084 298324 151136 298376
rect 88064 298256 88116 298308
rect 133236 298256 133288 298308
rect 88708 298188 88760 298240
rect 135904 298188 135956 298240
rect 67548 298120 67600 298172
rect 151268 298120 151320 298172
rect 157340 298052 157392 298104
rect 158628 298052 158680 298104
rect 176660 298052 176712 298104
rect 84200 297032 84252 297084
rect 153844 297032 153896 297084
rect 99012 296964 99064 297016
rect 123484 296964 123536 297016
rect 94504 296896 94556 296948
rect 144368 296896 144420 296948
rect 75184 296828 75236 296880
rect 134616 296828 134668 296880
rect 31024 296760 31076 296812
rect 97080 296760 97132 296812
rect 111248 296760 111300 296812
rect 159364 296760 159416 296812
rect 113824 296692 113876 296744
rect 120724 296692 120776 296744
rect 97724 295672 97776 295724
rect 129004 295672 129056 295724
rect 83556 295604 83608 295656
rect 126336 295604 126388 295656
rect 82268 295536 82320 295588
rect 138756 295536 138808 295588
rect 68560 295468 68612 295520
rect 129280 295468 129332 295520
rect 14464 295400 14516 295452
rect 92572 295400 92624 295452
rect 167736 295400 167788 295452
rect 67272 295332 67324 295384
rect 147128 295332 147180 295384
rect 295432 295332 295484 295384
rect 309876 295332 309928 295384
rect 73252 294720 73304 294772
rect 82176 294720 82228 294772
rect 79692 294652 79744 294704
rect 94596 294652 94648 294704
rect 71964 294584 72016 294636
rect 106924 294584 106976 294636
rect 111892 294312 111944 294364
rect 126428 294312 126480 294364
rect 91928 294244 91980 294296
rect 131764 294244 131816 294296
rect 80980 294176 81032 294228
rect 125048 294176 125100 294228
rect 78588 294108 78640 294160
rect 101404 294108 101456 294160
rect 105452 294108 105504 294160
rect 152464 294108 152516 294160
rect 65616 294040 65668 294092
rect 79324 294040 79376 294092
rect 93860 294040 93912 294092
rect 115848 294040 115900 294092
rect 116584 294040 116636 294092
rect 172060 294040 172112 294092
rect 75920 293972 75972 294024
rect 76748 293972 76800 294024
rect 82912 293972 82964 294024
rect 148416 293972 148468 294024
rect 158628 293972 158680 294024
rect 176660 293972 176712 294024
rect 295340 293972 295392 294024
rect 306380 293972 306432 294024
rect 84292 293904 84344 293956
rect 85212 293904 85264 293956
rect 85580 293904 85632 293956
rect 86500 293904 86552 293956
rect 109040 293904 109092 293956
rect 109684 293904 109736 293956
rect 114560 293904 114612 293956
rect 115388 293904 115440 293956
rect 3424 293224 3476 293276
rect 78588 293224 78640 293276
rect 87420 293224 87472 293276
rect 98736 293224 98788 293276
rect 115848 293224 115900 293276
rect 140044 293224 140096 293276
rect 3332 292816 3384 292868
rect 8944 292816 8996 292868
rect 112536 292816 112588 292868
rect 141424 292816 141476 292868
rect 102876 292748 102928 292800
rect 134708 292748 134760 292800
rect 117044 292680 117096 292732
rect 166264 292680 166316 292732
rect 68836 292612 68888 292664
rect 123668 292612 123720 292664
rect 67364 292544 67416 292596
rect 70676 292544 70728 292596
rect 98644 292544 98696 292596
rect 170496 292544 170548 292596
rect 71688 292476 71740 292528
rect 111156 292476 111208 292528
rect 121552 292476 121604 292528
rect 175924 292476 175976 292528
rect 101312 291864 101364 291916
rect 103612 291864 103664 291916
rect 67456 291184 67508 291236
rect 69756 291184 69808 291236
rect 110880 291864 110932 291916
rect 119344 291864 119396 291916
rect 119712 291864 119764 291916
rect 135996 291388 136048 291440
rect 127624 291320 127676 291372
rect 119804 291252 119856 291304
rect 152648 291252 152700 291304
rect 156604 291184 156656 291236
rect 168288 291184 168340 291236
rect 176660 291184 176712 291236
rect 26884 290436 26936 290488
rect 67732 290436 67784 290488
rect 302332 290436 302384 290488
rect 400864 290436 400916 290488
rect 121644 289960 121696 290012
rect 138664 289960 138716 290012
rect 121552 289892 121604 289944
rect 144276 289892 144328 289944
rect 53656 289824 53708 289876
rect 67640 289824 67692 289876
rect 120816 289824 120868 289876
rect 176660 289824 176712 289876
rect 295524 289824 295576 289876
rect 302332 289824 302384 289876
rect 121552 289756 121604 289808
rect 174544 289756 174596 289808
rect 67272 289280 67324 289332
rect 67548 289280 67600 289332
rect 64788 288396 64840 288448
rect 67640 288396 67692 288448
rect 121552 288396 121604 288448
rect 148508 288396 148560 288448
rect 121644 288328 121696 288380
rect 167644 288328 167696 288380
rect 3516 287648 3568 287700
rect 65616 287648 65668 287700
rect 52368 287036 52420 287088
rect 67640 287036 67692 287088
rect 121736 287036 121788 287088
rect 145564 287036 145616 287088
rect 22744 286968 22796 287020
rect 67548 286968 67600 287020
rect 121460 286424 121512 286476
rect 124128 286424 124180 286476
rect 136088 286424 136140 286476
rect 122748 286356 122800 286408
rect 171968 286356 172020 286408
rect 123576 286288 123628 286340
rect 177856 286288 177908 286340
rect 60648 285744 60700 285796
rect 67732 285744 67784 285796
rect 39948 285676 40000 285728
rect 67640 285676 67692 285728
rect 295524 285676 295576 285728
rect 309692 285676 309744 285728
rect 121552 285608 121604 285660
rect 171876 285608 171928 285660
rect 121460 284316 121512 284368
rect 167828 284316 167880 284368
rect 66168 284248 66220 284300
rect 67640 284248 67692 284300
rect 310980 283568 311032 283620
rect 355324 283568 355376 283620
rect 121460 282888 121512 282940
rect 174544 282888 174596 282940
rect 295524 282888 295576 282940
rect 310612 282888 310664 282940
rect 310980 282888 311032 282940
rect 64696 282820 64748 282872
rect 67640 282820 67692 282872
rect 167736 282820 167788 282872
rect 176660 282820 176712 282872
rect 121552 281596 121604 281648
rect 164884 281596 164936 281648
rect 121460 281528 121512 281580
rect 167644 281528 167696 281580
rect 295524 281528 295576 281580
rect 353944 281528 353996 281580
rect 54944 280236 54996 280288
rect 67640 280236 67692 280288
rect 121552 280236 121604 280288
rect 137376 280236 137428 280288
rect 55128 280168 55180 280220
rect 67732 280168 67784 280220
rect 121460 280168 121512 280220
rect 156696 280168 156748 280220
rect 129280 280100 129332 280152
rect 176752 280100 176804 280152
rect 48964 279420 49016 279472
rect 67916 279420 67968 279472
rect 121460 278740 121512 278792
rect 129096 278740 129148 278792
rect 295524 278740 295576 278792
rect 299480 278740 299532 278792
rect 152464 278060 152516 278112
rect 162676 278060 162728 278112
rect 121736 277992 121788 278044
rect 167736 277992 167788 278044
rect 56508 277448 56560 277500
rect 67640 277448 67692 277500
rect 46848 277380 46900 277432
rect 67732 277380 67784 277432
rect 121460 277380 121512 277432
rect 149888 277380 149940 277432
rect 162676 277380 162728 277432
rect 176660 277380 176712 277432
rect 305092 276632 305144 276684
rect 337384 276632 337436 276684
rect 64696 276088 64748 276140
rect 67640 276088 67692 276140
rect 121552 276088 121604 276140
rect 147220 276088 147272 276140
rect 53748 276020 53800 276072
rect 67732 276020 67784 276072
rect 121460 276020 121512 276072
rect 166540 276020 166592 276072
rect 295616 276020 295668 276072
rect 305092 276020 305144 276072
rect 172060 275952 172112 276004
rect 176660 275952 176712 276004
rect 121460 274728 121512 274780
rect 151176 274728 151228 274780
rect 63408 274660 63460 274712
rect 67640 274660 67692 274712
rect 121552 274660 121604 274712
rect 155500 274660 155552 274712
rect 121460 274388 121512 274440
rect 124864 274388 124916 274440
rect 18604 273912 18656 273964
rect 57244 273912 57296 273964
rect 64604 273300 64656 273352
rect 67640 273300 67692 273352
rect 57244 273232 57296 273284
rect 57612 273232 57664 273284
rect 67732 273232 67784 273284
rect 121460 273232 121512 273284
rect 143172 273232 143224 273284
rect 128360 273164 128412 273216
rect 176660 273164 176712 273216
rect 120908 272484 120960 272536
rect 128360 272484 128412 272536
rect 62028 271940 62080 271992
rect 67732 271940 67784 271992
rect 45376 271872 45428 271924
rect 67640 271872 67692 271924
rect 121460 271872 121512 271924
rect 155224 271872 155276 271924
rect 295616 271872 295668 271924
rect 300952 271872 301004 271924
rect 62304 271804 62356 271856
rect 62764 271804 62816 271856
rect 67732 271804 67784 271856
rect 50988 270512 51040 270564
rect 67640 270512 67692 270564
rect 121460 270512 121512 270564
rect 138848 270512 138900 270564
rect 66076 269152 66128 269204
rect 68192 269152 68244 269204
rect 121460 269152 121512 269204
rect 145748 269152 145800 269204
rect 44088 269084 44140 269136
rect 67640 269084 67692 269136
rect 121552 269084 121604 269136
rect 165068 269084 165120 269136
rect 295616 269084 295668 269136
rect 345664 269084 345716 269136
rect 66168 268200 66220 268252
rect 68192 268200 68244 268252
rect 121460 267792 121512 267844
rect 134800 267792 134852 267844
rect 161388 267792 161440 267844
rect 176660 267792 176712 267844
rect 46756 267724 46808 267776
rect 67640 267724 67692 267776
rect 120080 267724 120132 267776
rect 163688 267724 163740 267776
rect 63224 266976 63276 267028
rect 67640 266976 67692 267028
rect 121552 266432 121604 266484
rect 152464 266432 152516 266484
rect 121460 266364 121512 266416
rect 163504 266364 163556 266416
rect 45468 266296 45520 266348
rect 67732 266296 67784 266348
rect 123668 266296 123720 266348
rect 176660 266296 176712 266348
rect 121552 265004 121604 265056
rect 127808 265004 127860 265056
rect 53564 264936 53616 264988
rect 67640 264936 67692 264988
rect 121460 264936 121512 264988
rect 178684 264936 178736 264988
rect 295616 264936 295668 264988
rect 331864 264936 331916 264988
rect 48228 263644 48280 263696
rect 67640 263644 67692 263696
rect 21364 263576 21416 263628
rect 60464 263576 60516 263628
rect 67732 263576 67784 263628
rect 121552 263576 121604 263628
rect 148600 263576 148652 263628
rect 295616 263576 295668 263628
rect 305092 263576 305144 263628
rect 121460 263508 121512 263560
rect 169024 263508 169076 263560
rect 17224 262828 17276 262880
rect 53840 262828 53892 262880
rect 56416 262284 56468 262336
rect 67640 262284 67692 262336
rect 53840 262216 53892 262268
rect 54852 262216 54904 262268
rect 67732 262216 67784 262268
rect 121460 262216 121512 262268
rect 129280 262216 129332 262268
rect 121552 262148 121604 262200
rect 171784 262148 171836 262200
rect 160008 262080 160060 262132
rect 176660 262080 176712 262132
rect 3056 261468 3108 261520
rect 62764 261468 62816 261520
rect 121644 260856 121696 260908
rect 170588 260856 170640 260908
rect 295616 260856 295668 260908
rect 309784 260856 309836 260908
rect 13084 260788 13136 260840
rect 55036 260788 55088 260840
rect 67640 260788 67692 260840
rect 121460 260788 121512 260840
rect 170404 260788 170456 260840
rect 160008 259496 160060 259548
rect 176660 259496 176712 259548
rect 121460 259428 121512 259480
rect 169024 259428 169076 259480
rect 311164 259360 311216 259412
rect 579620 259360 579672 259412
rect 57704 258136 57756 258188
rect 67732 258136 67784 258188
rect 55036 258068 55088 258120
rect 67640 258068 67692 258120
rect 121460 258068 121512 258120
rect 171876 258068 171928 258120
rect 305644 257320 305696 257372
rect 340880 257320 340932 257372
rect 295708 257048 295760 257100
rect 298192 257048 298244 257100
rect 60372 256776 60424 256828
rect 67640 256776 67692 256828
rect 121552 256776 121604 256828
rect 140320 256776 140372 256828
rect 13084 256708 13136 256760
rect 69020 256708 69072 256760
rect 121460 256708 121512 256760
rect 159456 256708 159508 256760
rect 122104 255960 122156 256012
rect 169208 255960 169260 256012
rect 63316 255280 63368 255332
rect 67640 255280 67692 255332
rect 122472 254532 122524 254584
rect 169116 254532 169168 254584
rect 2780 254056 2832 254108
rect 4804 254056 4856 254108
rect 61936 253988 61988 254040
rect 67640 253988 67692 254040
rect 61844 253920 61896 253972
rect 67732 253920 67784 253972
rect 121460 253920 121512 253972
rect 170404 253920 170456 253972
rect 295708 253920 295760 253972
rect 335360 253920 335412 253972
rect 50528 253852 50580 253904
rect 50896 253852 50948 253904
rect 67640 253852 67692 253904
rect 295524 253444 295576 253496
rect 295708 253444 295760 253496
rect 25504 253172 25556 253224
rect 50528 253172 50580 253224
rect 121552 252628 121604 252680
rect 155316 252628 155368 252680
rect 50896 252560 50948 252612
rect 67640 252560 67692 252612
rect 121460 252560 121512 252612
rect 173256 252560 173308 252612
rect 64512 251880 64564 251932
rect 68100 251880 68152 251932
rect 59268 251812 59320 251864
rect 68376 251812 68428 251864
rect 302424 251812 302476 251864
rect 319444 251812 319496 251864
rect 56324 251268 56376 251320
rect 67640 251268 67692 251320
rect 121460 251200 121512 251252
rect 166448 251200 166500 251252
rect 296444 251200 296496 251252
rect 302424 251200 302476 251252
rect 120632 251132 120684 251184
rect 127716 251132 127768 251184
rect 295340 250860 295392 250912
rect 295524 250860 295576 250912
rect 60556 249772 60608 249824
rect 67640 249772 67692 249824
rect 121460 249772 121512 249824
rect 130660 249772 130712 249824
rect 172428 249772 172480 249824
rect 176660 249772 176712 249824
rect 295800 249772 295852 249824
rect 319444 249772 319496 249824
rect 68928 249704 68980 249756
rect 69664 249704 69716 249756
rect 65984 248616 66036 248668
rect 67824 248616 67876 248668
rect 121552 248480 121604 248532
rect 161020 248480 161072 248532
rect 121460 248412 121512 248464
rect 173348 248412 173400 248464
rect 121552 248344 121604 248396
rect 140136 248344 140188 248396
rect 296628 248344 296680 248396
rect 299664 248344 299716 248396
rect 324964 248344 325016 248396
rect 59176 247120 59228 247172
rect 67640 247120 67692 247172
rect 57796 247052 57848 247104
rect 67732 247052 67784 247104
rect 121460 247052 121512 247104
rect 144552 247052 144604 247104
rect 143080 246304 143132 246356
rect 174636 246304 174688 246356
rect 121460 245692 121512 245744
rect 142988 245692 143040 245744
rect 121552 245624 121604 245676
rect 149796 245624 149848 245676
rect 296904 245624 296956 245676
rect 467104 245624 467156 245676
rect 121460 245556 121512 245608
rect 162124 245556 162176 245608
rect 147036 245012 147088 245064
rect 171784 245012 171836 245064
rect 120724 244944 120776 244996
rect 158076 244944 158128 244996
rect 53104 244876 53156 244928
rect 59084 244876 59136 244928
rect 119804 244876 119856 244928
rect 162308 244876 162360 244928
rect 59084 244264 59136 244316
rect 67640 244264 67692 244316
rect 121552 244264 121604 244316
rect 170680 244264 170732 244316
rect 574744 244264 574796 244316
rect 579896 244264 579948 244316
rect 8944 244196 8996 244248
rect 69204 244196 69256 244248
rect 121552 242972 121604 243024
rect 147036 242972 147088 243024
rect 121460 242904 121512 242956
rect 179696 242904 179748 242956
rect 295340 242904 295392 242956
rect 299664 242904 299716 242956
rect 395344 242904 395396 242956
rect 121552 242836 121604 242888
rect 160744 242836 160796 242888
rect 121460 242768 121512 242820
rect 158628 242768 158680 242820
rect 160928 242768 160980 242820
rect 147128 242700 147180 242752
rect 176844 242700 176896 242752
rect 143172 242224 143224 242276
rect 152740 242224 152792 242276
rect 125048 242156 125100 242208
rect 154120 242156 154172 242208
rect 61752 241476 61804 241528
rect 67732 241476 67784 241528
rect 57888 241408 57940 241460
rect 67640 241408 67692 241460
rect 163688 241408 163740 241460
rect 295524 241408 295576 241460
rect 127808 240796 127860 240848
rect 156788 240796 156840 240848
rect 140228 240728 140280 240780
rect 182824 240592 182876 240644
rect 179696 240320 179748 240372
rect 69848 240184 69900 240236
rect 121460 240116 121512 240168
rect 144460 240116 144512 240168
rect 179880 240116 179932 240168
rect 152648 240048 152700 240100
rect 295708 240048 295760 240100
rect 75276 239912 75328 239964
rect 118976 239912 119028 239964
rect 119804 239912 119856 239964
rect 64512 239436 64564 239488
rect 116584 239436 116636 239488
rect 3332 239368 3384 239420
rect 70308 239368 70360 239420
rect 118608 239368 118660 239420
rect 135260 239368 135312 239420
rect 287704 239368 287756 239420
rect 296812 239368 296864 239420
rect 121552 238960 121604 239012
rect 323584 238960 323636 239012
rect 60464 238892 60516 238944
rect 252560 238892 252612 238944
rect 61936 238824 61988 238876
rect 262220 238824 262272 238876
rect 262772 238824 262824 238876
rect 278872 238824 278924 238876
rect 279976 238824 280028 238876
rect 310520 238824 310572 238876
rect 58624 238756 58676 238808
rect 81532 238756 81584 238808
rect 82268 238756 82320 238808
rect 109040 238756 109092 238808
rect 109960 238756 110012 238808
rect 120816 238756 120868 238808
rect 174544 238756 174596 238808
rect 215300 238756 215352 238808
rect 525064 238756 525116 238808
rect 62764 238688 62816 238740
rect 86776 238688 86828 238740
rect 114468 238688 114520 238740
rect 118608 238688 118660 238740
rect 190000 238688 190052 238740
rect 582564 238688 582616 238740
rect 70308 238620 70360 238672
rect 103520 238620 103572 238672
rect 104716 238620 104768 238672
rect 107384 238620 107436 238672
rect 130568 238620 130620 238672
rect 176016 238620 176068 238672
rect 223856 238620 223908 238672
rect 236000 238620 236052 238672
rect 582472 238620 582524 238672
rect 117688 238552 117740 238604
rect 250812 238552 250864 238604
rect 99012 238484 99064 238536
rect 120908 238484 120960 238536
rect 170496 238484 170548 238536
rect 195980 238484 196032 238536
rect 110604 238416 110656 238468
rect 126244 238416 126296 238468
rect 89352 238348 89404 238400
rect 148324 238348 148376 238400
rect 86132 238212 86184 238264
rect 95700 238212 95752 238264
rect 75828 238144 75880 238196
rect 86224 238144 86276 238196
rect 70676 238076 70728 238128
rect 147128 238076 147180 238128
rect 4804 238008 4856 238060
rect 112536 238008 112588 238060
rect 155408 238008 155460 238060
rect 189724 238008 189776 238060
rect 110604 237804 110656 237856
rect 111064 237804 111116 237856
rect 104164 237396 104216 237448
rect 106924 237396 106976 237448
rect 215944 237396 215996 237448
rect 217048 237396 217100 237448
rect 224132 237396 224184 237448
rect 240048 237396 240100 237448
rect 291844 237396 291896 237448
rect 292580 237396 292632 237448
rect 91928 237328 91980 237380
rect 134524 237328 134576 237380
rect 166356 237328 166408 237380
rect 580356 237328 580408 237380
rect 112536 237260 112588 237312
rect 144184 237260 144236 237312
rect 161020 237260 161072 237312
rect 314660 237260 314712 237312
rect 63224 237192 63276 237244
rect 191932 237192 191984 237244
rect 233884 237192 233936 237244
rect 364340 237192 364392 237244
rect 188344 237124 188396 237176
rect 254400 237124 254452 237176
rect 173348 236716 173400 236768
rect 192484 236716 192536 236768
rect 40040 236648 40092 236700
rect 95056 236648 95108 236700
rect 95792 236648 95844 236700
rect 141516 236648 141568 236700
rect 242256 236648 242308 236700
rect 113824 235900 113876 235952
rect 300860 235900 300912 235952
rect 72608 235832 72660 235884
rect 123576 235832 123628 235884
rect 159456 235832 159508 235884
rect 310612 235832 310664 235884
rect 95056 235764 95108 235816
rect 142804 235764 142856 235816
rect 169208 235764 169260 235816
rect 295616 235764 295668 235816
rect 276296 235696 276348 235748
rect 276664 235696 276716 235748
rect 305000 235696 305052 235748
rect 170588 235356 170640 235408
rect 198004 235356 198056 235408
rect 60372 235288 60424 235340
rect 159548 235288 159600 235340
rect 171876 235288 171928 235340
rect 222844 235288 222896 235340
rect 152556 235220 152608 235272
rect 260104 235220 260156 235272
rect 46756 234540 46808 234592
rect 303712 234540 303764 234592
rect 91284 234472 91336 234524
rect 129188 234472 129240 234524
rect 151268 234472 151320 234524
rect 298192 234472 298244 234524
rect 264980 234404 265032 234456
rect 265624 234404 265676 234456
rect 306472 234404 306524 234456
rect 46204 234132 46256 234184
rect 46756 234132 46808 234184
rect 149888 233996 149940 234048
rect 186964 233996 187016 234048
rect 69020 233928 69072 233980
rect 69756 233928 69808 233980
rect 75920 233928 75972 233980
rect 77116 233928 77168 233980
rect 77300 233928 77352 233980
rect 78404 233928 78456 233980
rect 78680 233928 78732 233980
rect 79692 233928 79744 233980
rect 84292 233928 84344 233980
rect 85488 233928 85540 233980
rect 93860 233928 93912 233980
rect 94504 233928 94556 233980
rect 96620 233928 96672 233980
rect 97724 233928 97776 233980
rect 100760 233928 100812 233980
rect 101588 233928 101640 233980
rect 102140 233928 102192 233980
rect 102876 233928 102928 233980
rect 104900 233928 104952 233980
rect 106096 233928 106148 233980
rect 114560 233928 114612 233980
rect 115756 233928 115808 233980
rect 174636 233928 174688 233980
rect 255964 233928 256016 233980
rect 62028 233860 62080 233912
rect 196716 233860 196768 233912
rect 289820 233656 289872 233708
rect 294144 233656 294196 233708
rect 92480 233384 92532 233436
rect 93216 233384 93268 233436
rect 59084 233180 59136 233232
rect 218980 233180 219032 233232
rect 223856 233180 223908 233232
rect 582656 233180 582708 233232
rect 86776 233112 86828 233164
rect 210608 233112 210660 233164
rect 240048 233112 240100 233164
rect 582380 233112 582432 233164
rect 115112 233044 115164 233096
rect 236000 233044 236052 233096
rect 395344 233044 395396 233096
rect 579620 233044 579672 233096
rect 171968 232976 172020 233028
rect 271144 232976 271196 233028
rect 278780 232636 278832 232688
rect 294236 232636 294288 232688
rect 274640 232568 274692 232620
rect 293224 232568 293276 232620
rect 68652 232500 68704 232552
rect 328552 232500 328604 232552
rect 84108 231820 84160 231872
rect 84844 231820 84896 231872
rect 61844 231752 61896 231804
rect 302424 231752 302476 231804
rect 83556 231684 83608 231736
rect 130384 231684 130436 231736
rect 179880 231684 179932 231736
rect 295432 231684 295484 231736
rect 118332 231616 118384 231668
rect 224132 231616 224184 231668
rect 167828 231072 167880 231124
rect 224224 231072 224276 231124
rect 319444 231072 319496 231124
rect 333980 231072 334032 231124
rect 54852 230392 54904 230444
rect 289912 230392 289964 230444
rect 104716 230324 104768 230376
rect 293132 230324 293184 230376
rect 98368 230256 98420 230308
rect 233884 230256 233936 230308
rect 170680 229712 170732 229764
rect 264336 229712 264388 229764
rect 73160 229304 73212 229356
rect 73896 229304 73948 229356
rect 81532 229032 81584 229084
rect 277400 229032 277452 229084
rect 57612 228964 57664 229016
rect 241520 228964 241572 229016
rect 100300 228488 100352 228540
rect 163688 228488 163740 228540
rect 165068 228488 165120 228540
rect 206284 228488 206336 228540
rect 108672 228420 108724 228472
rect 328460 228420 328512 228472
rect 67364 228352 67416 228404
rect 98644 228352 98696 228404
rect 162676 228352 162728 228404
rect 582380 228352 582432 228404
rect 86224 227672 86276 227724
rect 302240 227672 302292 227724
rect 92572 227128 92624 227180
rect 220084 227128 220136 227180
rect 280160 227128 280212 227180
rect 311900 227128 311952 227180
rect 113180 227060 113232 227112
rect 283564 227060 283616 227112
rect 66076 226992 66128 227044
rect 324596 226992 324648 227044
rect 155500 226244 155552 226296
rect 296904 226244 296956 226296
rect 182824 225700 182876 225752
rect 319444 225700 319496 225752
rect 156788 225632 156840 225684
rect 336740 225632 336792 225684
rect 67272 225564 67324 225616
rect 253204 225564 253256 225616
rect 81440 224884 81492 224936
rect 278872 224884 278924 224936
rect 147220 224816 147272 224868
rect 299664 224816 299716 224868
rect 129280 224340 129332 224392
rect 257344 224340 257396 224392
rect 97080 224272 97132 224324
rect 129188 224272 129240 224324
rect 164976 224272 165028 224324
rect 311164 224272 311216 224324
rect 3608 224204 3660 224256
rect 120172 224204 120224 224256
rect 136088 224204 136140 224256
rect 580356 224204 580408 224256
rect 160928 223524 160980 223576
rect 574744 223524 574796 223576
rect 69112 222980 69164 223032
rect 249800 222980 249852 223032
rect 56416 222912 56468 222964
rect 240784 222912 240836 222964
rect 256700 222912 256752 222964
rect 278044 222912 278096 222964
rect 131856 222844 131908 222896
rect 345020 222844 345072 222896
rect 162216 221620 162268 221672
rect 214564 221620 214616 221672
rect 88064 221552 88116 221604
rect 247684 221552 247736 221604
rect 64696 221484 64748 221536
rect 324412 221484 324464 221536
rect 77760 221416 77812 221468
rect 351920 221416 351972 221468
rect 111892 220328 111944 220380
rect 267740 220328 267792 220380
rect 79048 220260 79100 220312
rect 242164 220260 242216 220312
rect 159364 220192 159416 220244
rect 346492 220192 346544 220244
rect 56324 220124 56376 220176
rect 313924 220124 313976 220176
rect 179052 220056 179104 220108
rect 580448 220056 580500 220108
rect 76012 219376 76064 219428
rect 150348 219376 150400 219428
rect 471244 219376 471296 219428
rect 580172 219376 580224 219428
rect 170404 218968 170456 219020
rect 273352 218968 273404 219020
rect 153936 218900 153988 218952
rect 318064 218900 318116 218952
rect 65984 218832 66036 218884
rect 278872 218832 278924 218884
rect 48228 218764 48280 218816
rect 343640 218764 343692 218816
rect 150348 218696 150400 218748
rect 582472 218696 582524 218748
rect 145656 217540 145708 217592
rect 266452 217540 266504 217592
rect 148600 217472 148652 217524
rect 270500 217472 270552 217524
rect 138756 217404 138808 217456
rect 274732 217404 274784 217456
rect 106924 217336 106976 217388
rect 160744 217336 160796 217388
rect 160836 217336 160888 217388
rect 356060 217336 356112 217388
rect 102232 217268 102284 217320
rect 319536 217268 319588 217320
rect 100852 216112 100904 216164
rect 255320 216112 255372 216164
rect 159548 216044 159600 216096
rect 345112 216044 345164 216096
rect 116584 215976 116636 216028
rect 315396 215976 315448 216028
rect 134800 215908 134852 215960
rect 338120 215908 338172 215960
rect 3332 215228 3384 215280
rect 21364 215228 21416 215280
rect 258080 215024 258132 215076
rect 264244 215024 264296 215076
rect 144276 214752 144328 214804
rect 210424 214752 210476 214804
rect 163688 214684 163740 214736
rect 276020 214684 276072 214736
rect 114560 214616 114612 214668
rect 325700 214616 325752 214668
rect 46848 214548 46900 214600
rect 311256 214548 311308 214600
rect 255964 213868 256016 213920
rect 258724 213868 258776 213920
rect 152740 213392 152792 213444
rect 236644 213392 236696 213444
rect 149704 213324 149756 213376
rect 277400 213324 277452 213376
rect 99380 213256 99432 213308
rect 325884 213256 325936 213308
rect 86960 213188 87012 213240
rect 322940 213188 322992 213240
rect 124956 211896 125008 211948
rect 273260 211896 273312 211948
rect 89812 211828 89864 211880
rect 274824 211828 274876 211880
rect 61752 211760 61804 211812
rect 259460 211760 259512 211812
rect 260104 211760 260156 211812
rect 332600 211760 332652 211812
rect 231860 210604 231912 210656
rect 282920 210604 282972 210656
rect 133236 210536 133288 210588
rect 232504 210536 232556 210588
rect 4804 210468 4856 210520
rect 83464 210468 83516 210520
rect 144552 210468 144604 210520
rect 246396 210468 246448 210520
rect 74632 210400 74684 210452
rect 246304 210400 246356 210452
rect 271880 210400 271932 210452
rect 294052 210400 294104 210452
rect 138848 209176 138900 209228
rect 258172 209176 258224 209228
rect 67456 209108 67508 209160
rect 247776 209108 247828 209160
rect 103704 209040 103756 209092
rect 327080 209040 327132 209092
rect 237380 207952 237432 208004
rect 279424 207952 279476 208004
rect 198004 207884 198056 207936
rect 305644 207884 305696 207936
rect 151176 207816 151228 207868
rect 281632 207816 281684 207868
rect 55036 207748 55088 207800
rect 239404 207748 239456 207800
rect 126428 207680 126480 207732
rect 339684 207680 339736 207732
rect 53656 207612 53708 207664
rect 271972 207612 272024 207664
rect 281540 207612 281592 207664
rect 342260 207612 342312 207664
rect 45376 206388 45428 206440
rect 228364 206388 228416 206440
rect 260840 206388 260892 206440
rect 289084 206388 289136 206440
rect 160744 206320 160796 206372
rect 347780 206320 347832 206372
rect 75920 206252 75972 206304
rect 327172 206252 327224 206304
rect 94044 205164 94096 205216
rect 189908 205164 189960 205216
rect 189724 205096 189776 205148
rect 339500 205096 339552 205148
rect 70400 205028 70452 205080
rect 252836 205028 252888 205080
rect 59176 204960 59228 205012
rect 259552 204960 259604 205012
rect 118700 204892 118752 204944
rect 328644 204892 328696 204944
rect 153844 203804 153896 203856
rect 243544 203804 243596 203856
rect 248420 203804 248472 203856
rect 291200 203804 291252 203856
rect 166540 203736 166592 203788
rect 342444 203736 342496 203788
rect 122104 203668 122156 203720
rect 325792 203668 325844 203720
rect 57704 203600 57756 203652
rect 273444 203600 273496 203652
rect 71780 203532 71832 203584
rect 327264 203532 327316 203584
rect 245660 202444 245712 202496
rect 308588 202444 308640 202496
rect 146944 202376 146996 202428
rect 281540 202376 281592 202428
rect 102140 202308 102192 202360
rect 252652 202308 252704 202360
rect 160008 202240 160060 202292
rect 354680 202240 354732 202292
rect 145564 202172 145616 202224
rect 343732 202172 343784 202224
rect 60556 202104 60608 202156
rect 276112 202104 276164 202156
rect 131764 200812 131816 200864
rect 258264 200812 258316 200864
rect 56508 200744 56560 200796
rect 231124 200744 231176 200796
rect 142896 199520 142948 199572
rect 269120 199520 269172 199572
rect 162308 199452 162360 199504
rect 342352 199452 342404 199504
rect 96528 199384 96580 199436
rect 582380 199384 582432 199436
rect 126336 198160 126388 198212
rect 239496 198160 239548 198212
rect 140320 198092 140372 198144
rect 264980 198092 265032 198144
rect 115940 198024 115992 198076
rect 260932 198024 260984 198076
rect 151084 197956 151136 198008
rect 319628 197956 319680 198008
rect 130660 196936 130712 196988
rect 250076 196936 250128 196988
rect 192484 196868 192536 196920
rect 312544 196868 312596 196920
rect 66168 196800 66220 196852
rect 251180 196800 251232 196852
rect 123484 196732 123536 196784
rect 349344 196732 349396 196784
rect 69664 196664 69716 196716
rect 320824 196664 320876 196716
rect 50896 196596 50948 196648
rect 334164 196596 334216 196648
rect 134616 195508 134668 195560
rect 267832 195508 267884 195560
rect 89720 195440 89772 195492
rect 263600 195440 263652 195492
rect 158076 195372 158128 195424
rect 347872 195372 347924 195424
rect 104900 195304 104952 195356
rect 336832 195304 336884 195356
rect 92480 195236 92532 195288
rect 328736 195236 328788 195288
rect 196716 194148 196768 194200
rect 244924 194148 244976 194200
rect 253204 194148 253256 194200
rect 329932 194148 329984 194200
rect 129188 194080 129240 194132
rect 262404 194080 262456 194132
rect 167736 194012 167788 194064
rect 318156 194012 318208 194064
rect 147128 193944 147180 193996
rect 331312 193944 331364 193996
rect 44088 193876 44140 193928
rect 270592 193876 270644 193928
rect 96620 193808 96672 193860
rect 331220 193808 331272 193860
rect 127624 192584 127676 192636
rect 272064 192584 272116 192636
rect 93952 192516 94004 192568
rect 254124 192516 254176 192568
rect 133144 192448 133196 192500
rect 341064 192448 341116 192500
rect 142988 191360 143040 191412
rect 242256 191360 242308 191412
rect 149796 191292 149848 191344
rect 260840 191292 260892 191344
rect 137284 191224 137336 191276
rect 255504 191224 255556 191276
rect 264336 191224 264388 191276
rect 338212 191224 338264 191276
rect 227720 191156 227772 191208
rect 346400 191156 346452 191208
rect 135904 191088 135956 191140
rect 343824 191088 343876 191140
rect 102048 190476 102100 190528
rect 203616 190476 203668 190528
rect 211068 190068 211120 190120
rect 244280 190068 244332 190120
rect 229100 190000 229152 190052
rect 268384 190000 268436 190052
rect 144460 189932 144512 189984
rect 261024 189932 261076 189984
rect 141424 189864 141476 189916
rect 269212 189864 269264 189916
rect 21364 189796 21416 189848
rect 111064 189796 111116 189848
rect 173256 189796 173308 189848
rect 324504 189796 324556 189848
rect 84292 189728 84344 189780
rect 254032 189728 254084 189780
rect 257344 189728 257396 189780
rect 340972 189728 341024 189780
rect 107568 189184 107620 189236
rect 171876 189184 171928 189236
rect 118608 189116 118660 189168
rect 189816 189116 189868 189168
rect 133788 189048 133840 189100
rect 214656 189048 214708 189100
rect 3148 188980 3200 189032
rect 14464 188980 14516 189032
rect 206284 188572 206336 188624
rect 263692 188572 263744 188624
rect 138664 188504 138716 188556
rect 258080 188504 258132 188556
rect 258724 188504 258776 188556
rect 339776 188504 339828 188556
rect 135996 188436 136048 188488
rect 266544 188436 266596 188488
rect 18604 188368 18656 188420
rect 109040 188368 109092 188420
rect 152464 188368 152516 188420
rect 349436 188368 349488 188420
rect 80152 188300 80204 188352
rect 327356 188300 327408 188352
rect 106188 187756 106240 187808
rect 167736 187756 167788 187808
rect 100668 187688 100720 187740
rect 170404 187688 170456 187740
rect 157248 187280 157300 187332
rect 189724 187280 189776 187332
rect 148416 187212 148468 187264
rect 252744 187212 252796 187264
rect 129096 187144 129148 187196
rect 256700 187144 256752 187196
rect 63408 187076 63460 187128
rect 249064 187076 249116 187128
rect 95332 187008 95384 187060
rect 321284 187008 321336 187060
rect 73252 186940 73304 186992
rect 320180 186940 320232 186992
rect 155316 185852 155368 185904
rect 255596 185852 255648 185904
rect 107660 185784 107712 185836
rect 346584 185784 346636 185836
rect 68928 185716 68980 185768
rect 321744 185716 321796 185768
rect 69020 185648 69072 185700
rect 323124 185648 323176 185700
rect 59268 185580 59320 185632
rect 337016 185580 337068 185632
rect 134524 184900 134576 184952
rect 210608 184900 210660 184952
rect 222844 184424 222896 184476
rect 350632 184424 350684 184476
rect 163504 184356 163556 184408
rect 334256 184356 334308 184408
rect 63316 184288 63368 184340
rect 256792 184288 256844 184340
rect 84200 184220 84252 184272
rect 325976 184220 326028 184272
rect 88340 184152 88392 184204
rect 346676 184152 346728 184204
rect 114468 183608 114520 183660
rect 169300 183608 169352 183660
rect 128268 183540 128320 183592
rect 214748 183540 214800 183592
rect 220084 183132 220136 183184
rect 258356 183132 258408 183184
rect 156696 183064 156748 183116
rect 245660 183064 245712 183116
rect 172428 182996 172480 183048
rect 282184 182996 282236 183048
rect 189908 182928 189960 182980
rect 334072 182928 334124 182980
rect 148508 182860 148560 182912
rect 338304 182860 338356 182912
rect 93860 182792 93912 182844
rect 330116 182792 330168 182844
rect 127808 182180 127860 182232
rect 206468 182180 206520 182232
rect 228364 181704 228416 181756
rect 265072 181704 265124 181756
rect 140044 181636 140096 181688
rect 249340 181636 249392 181688
rect 224224 181568 224276 181620
rect 332784 181568 332836 181620
rect 156604 181500 156656 181552
rect 341156 181500 341208 181552
rect 147036 181432 147088 181484
rect 342536 181432 342588 181484
rect 116952 180956 117004 181008
rect 166540 180956 166592 181008
rect 112996 180888 113048 180940
rect 167828 180888 167880 180940
rect 129464 180820 129516 180872
rect 206560 180820 206612 180872
rect 162768 180276 162820 180328
rect 203524 180276 203576 180328
rect 231124 180276 231176 180328
rect 262496 180276 262548 180328
rect 169116 180208 169168 180260
rect 318340 180208 318392 180260
rect 64788 180140 64840 180192
rect 251272 180140 251324 180192
rect 283564 180140 283616 180192
rect 335452 180140 335504 180192
rect 157984 180072 158036 180124
rect 345204 180072 345256 180124
rect 113916 179528 113968 179580
rect 166356 179528 166408 179580
rect 110696 179460 110748 179512
rect 166264 179460 166316 179512
rect 97816 179392 97868 179444
rect 169208 179392 169260 179444
rect 373264 179324 373316 179376
rect 580172 179324 580224 179376
rect 246396 178984 246448 179036
rect 252560 178984 252612 179036
rect 240784 178916 240836 178968
rect 256884 178916 256936 178968
rect 210424 178848 210476 178900
rect 249984 178848 250036 178900
rect 312544 178848 312596 178900
rect 339592 178848 339644 178900
rect 167644 178780 167696 178832
rect 251456 178780 251508 178832
rect 305644 178780 305696 178832
rect 335544 178780 335596 178832
rect 129004 178712 129056 178764
rect 318708 178712 318760 178764
rect 78680 178644 78732 178696
rect 343916 178644 343968 178696
rect 109868 178236 109920 178288
rect 162768 178236 162820 178288
rect 148232 178168 148284 178220
rect 206284 178168 206336 178220
rect 122012 178100 122064 178152
rect 196716 178100 196768 178152
rect 124956 178032 125008 178084
rect 214932 178032 214984 178084
rect 119712 177964 119764 178016
rect 134524 177964 134576 178016
rect 217968 177964 218020 178016
rect 220820 177964 220872 178016
rect 236644 177624 236696 177676
rect 249248 177624 249300 177676
rect 242256 177556 242308 177608
rect 256976 177556 257028 177608
rect 168288 177488 168340 177540
rect 202144 177488 202196 177540
rect 216588 177488 216640 177540
rect 224960 177488 225012 177540
rect 242164 177488 242216 177540
rect 262312 177488 262364 177540
rect 318064 177488 318116 177540
rect 169024 177420 169076 177472
rect 251364 177420 251416 177472
rect 318340 177420 318392 177472
rect 321836 177420 321888 177472
rect 332876 177420 332928 177472
rect 164884 177352 164936 177404
rect 249156 177352 249208 177404
rect 315396 177352 315448 177404
rect 331404 177352 331456 177404
rect 1308 177284 1360 177336
rect 120080 177284 120132 177336
rect 166448 177284 166500 177336
rect 330024 177284 330076 177336
rect 108120 177012 108172 177064
rect 165252 177012 165304 177064
rect 132040 176944 132092 176996
rect 165436 176944 165488 176996
rect 123024 176876 123076 176928
rect 165528 176876 165580 176928
rect 125876 176808 125928 176860
rect 167920 176808 167972 176860
rect 158996 176740 159048 176792
rect 187056 176740 187108 176792
rect 134432 176672 134484 176724
rect 195980 176672 196032 176724
rect 318156 176672 318208 176724
rect 321560 176672 321612 176724
rect 135720 176604 135772 176656
rect 213920 176604 213972 176656
rect 245660 176604 245712 176656
rect 249892 176604 249944 176656
rect 311256 176604 311308 176656
rect 321468 176604 321520 176656
rect 162768 176196 162820 176248
rect 206376 176196 206428 176248
rect 120816 176128 120868 176180
rect 167644 176128 167696 176180
rect 115756 176060 115808 176112
rect 166448 176060 166500 176112
rect 249064 176060 249116 176112
rect 253940 176060 253992 176112
rect 104624 175992 104676 176044
rect 169024 175992 169076 176044
rect 246304 175992 246356 176044
rect 255412 175992 255464 176044
rect 305644 175992 305696 176044
rect 306380 175992 306432 176044
rect 307576 175992 307628 176044
rect 319628 175992 319680 176044
rect 326068 175992 326120 176044
rect 130752 175924 130804 175976
rect 214012 175924 214064 175976
rect 247684 175924 247736 175976
rect 259644 175924 259696 175976
rect 319536 175924 319588 175976
rect 335636 175924 335688 175976
rect 318708 175856 318760 175908
rect 321928 175856 321980 175908
rect 243544 175788 243596 175840
rect 248052 175788 248104 175840
rect 195980 175176 196032 175228
rect 213920 175176 213972 175228
rect 3516 150356 3568 150408
rect 26884 150356 26936 150408
rect 3516 137912 3568 137964
rect 13084 137912 13136 137964
rect 59268 125604 59320 125656
rect 66168 125604 66220 125656
rect 63316 124176 63368 124228
rect 65524 124176 65576 124228
rect 62028 122816 62080 122868
rect 66076 122816 66128 122868
rect 63408 121456 63460 121508
rect 66076 121456 66128 121508
rect 3148 111732 3200 111784
rect 21364 111732 21416 111784
rect 2780 97724 2832 97776
rect 4804 97724 4856 97776
rect 165436 174496 165488 174548
rect 213920 174496 213972 174548
rect 288072 174020 288124 174072
rect 307668 174020 307720 174072
rect 282276 173952 282328 174004
rect 306748 173952 306800 174004
rect 264428 173884 264480 173936
rect 307576 173884 307628 173936
rect 324320 173816 324372 173868
rect 326068 173816 326120 173868
rect 252100 173680 252152 173732
rect 256700 173680 256752 173732
rect 165252 173136 165304 173188
rect 214288 173136 214340 173188
rect 271236 172592 271288 172644
rect 307300 172592 307352 172644
rect 269856 172524 269908 172576
rect 306932 172524 306984 172576
rect 206560 172456 206612 172508
rect 213920 172456 213972 172508
rect 252468 171504 252520 171556
rect 258172 171504 258224 171556
rect 280804 171232 280856 171284
rect 306932 171232 306984 171284
rect 265624 171164 265676 171216
rect 307668 171164 307720 171216
rect 168012 171096 168064 171148
rect 210516 171096 210568 171148
rect 261668 171096 261720 171148
rect 307576 171096 307628 171148
rect 167920 171028 167972 171080
rect 214012 171028 214064 171080
rect 206468 170960 206520 171012
rect 213920 170960 213972 171012
rect 251364 170892 251416 170944
rect 251548 170892 251600 170944
rect 251732 170892 251784 170944
rect 255504 170892 255556 170944
rect 294604 170348 294656 170400
rect 306564 170348 306616 170400
rect 251364 170280 251416 170332
rect 253940 170280 253992 170332
rect 251824 169804 251876 169856
rect 259552 169804 259604 169856
rect 267096 169804 267148 169856
rect 307668 169804 307720 169856
rect 260380 169736 260432 169788
rect 306748 169736 306800 169788
rect 252284 169668 252336 169720
rect 262404 169668 262456 169720
rect 324320 169668 324372 169720
rect 337016 169668 337068 169720
rect 169116 168988 169168 169040
rect 214656 168988 214708 169040
rect 283564 168512 283616 168564
rect 307668 168512 307720 168564
rect 273904 168444 273956 168496
rect 307484 168444 307536 168496
rect 262864 168376 262916 168428
rect 307576 168376 307628 168428
rect 167644 168308 167696 168360
rect 214012 168308 214064 168360
rect 251916 168308 251968 168360
rect 255596 168308 255648 168360
rect 324320 168308 324372 168360
rect 334164 168308 334216 168360
rect 196716 168240 196768 168292
rect 213920 168240 213972 168292
rect 252468 167220 252520 167272
rect 258264 167220 258316 167272
rect 291936 167152 291988 167204
rect 307300 167152 307352 167204
rect 278228 167084 278280 167136
rect 307668 167084 307720 167136
rect 275284 167016 275336 167068
rect 307484 167016 307536 167068
rect 166540 166948 166592 167000
rect 214012 166948 214064 167000
rect 252100 166948 252152 167000
rect 261024 166948 261076 167000
rect 189816 166880 189868 166932
rect 213920 166880 213972 166932
rect 210608 166812 210660 166864
rect 214104 166812 214156 166864
rect 252376 166744 252428 166796
rect 256884 166744 256936 166796
rect 252468 166472 252520 166524
rect 258356 166472 258408 166524
rect 269948 165656 270000 165708
rect 307576 165656 307628 165708
rect 259092 165588 259144 165640
rect 307668 165588 307720 165640
rect 166448 165520 166500 165572
rect 213920 165520 213972 165572
rect 252468 165520 252520 165572
rect 266544 165520 266596 165572
rect 324320 165520 324372 165572
rect 335636 165520 335688 165572
rect 169300 165452 169352 165504
rect 214012 165452 214064 165504
rect 252100 165452 252152 165504
rect 263600 165452 263652 165504
rect 251732 165384 251784 165436
rect 262496 165384 262548 165436
rect 271328 164908 271380 164960
rect 306932 164908 306984 164960
rect 257436 164840 257488 164892
rect 307484 164840 307536 164892
rect 300124 164296 300176 164348
rect 307668 164296 307720 164348
rect 287796 164228 287848 164280
rect 307300 164228 307352 164280
rect 166356 164160 166408 164212
rect 213920 164160 213972 164212
rect 252192 164160 252244 164212
rect 270500 164160 270552 164212
rect 324412 164160 324464 164212
rect 331404 164160 331456 164212
rect 167828 164092 167880 164144
rect 214012 164092 214064 164144
rect 324320 164092 324372 164144
rect 329932 164092 329984 164144
rect 290464 163004 290516 163056
rect 307300 163004 307352 163056
rect 272524 162936 272576 162988
rect 306748 162936 306800 162988
rect 265716 162868 265768 162920
rect 307668 162868 307720 162920
rect 166264 162800 166316 162852
rect 213920 162800 213972 162852
rect 252468 162800 252520 162852
rect 263692 162800 263744 162852
rect 324412 162800 324464 162852
rect 342536 162800 342588 162852
rect 206376 162732 206428 162784
rect 214012 162732 214064 162784
rect 324320 162732 324372 162784
rect 332876 162732 332928 162784
rect 262956 162120 263008 162172
rect 307116 162120 307168 162172
rect 289268 161508 289320 161560
rect 307484 161508 307536 161560
rect 279608 161440 279660 161492
rect 307668 161440 307720 161492
rect 171876 161372 171928 161424
rect 213920 161372 213972 161424
rect 252468 161372 252520 161424
rect 260932 161372 260984 161424
rect 324320 161372 324372 161424
rect 346492 161372 346544 161424
rect 324412 161304 324464 161356
rect 332784 161304 332836 161356
rect 260104 160760 260156 160812
rect 306472 160760 306524 160812
rect 254860 160692 254912 160744
rect 307208 160692 307260 160744
rect 303068 160148 303120 160200
rect 307668 160148 307720 160200
rect 276848 160080 276900 160132
rect 307576 160080 307628 160132
rect 167736 160012 167788 160064
rect 213920 160012 213972 160064
rect 324320 160012 324372 160064
rect 331312 160012 331364 160064
rect 169024 159944 169076 159996
rect 214012 159944 214064 159996
rect 251088 159332 251140 159384
rect 259644 159332 259696 159384
rect 278320 159332 278372 159384
rect 307392 159332 307444 159384
rect 264336 158788 264388 158840
rect 306932 158788 306984 158840
rect 261760 158720 261812 158772
rect 307668 158720 307720 158772
rect 203616 158652 203668 158704
rect 213920 158652 213972 158704
rect 251916 158652 251968 158704
rect 256792 158652 256844 158704
rect 324412 158652 324464 158704
rect 341156 158652 341208 158704
rect 324320 158584 324372 158636
rect 334256 158584 334308 158636
rect 287980 157496 288032 157548
rect 307668 157496 307720 157548
rect 260196 157428 260248 157480
rect 307484 157428 307536 157480
rect 257344 157360 257396 157412
rect 306932 157360 306984 157412
rect 170404 157292 170456 157344
rect 213920 157292 213972 157344
rect 252468 157292 252520 157344
rect 272064 157292 272116 157344
rect 252376 157224 252428 157276
rect 265072 157224 265124 157276
rect 324320 157224 324372 157276
rect 339776 157224 339828 157276
rect 285128 156068 285180 156120
rect 307484 156068 307536 156120
rect 258724 156000 258776 156052
rect 307576 156000 307628 156052
rect 254676 155932 254728 155984
rect 307668 155932 307720 155984
rect 169208 155864 169260 155916
rect 214012 155864 214064 155916
rect 251916 155864 251968 155916
rect 255320 155864 255372 155916
rect 324320 155864 324372 155916
rect 338396 155864 338448 155916
rect 170496 155796 170548 155848
rect 213920 155796 213972 155848
rect 251180 155796 251232 155848
rect 254032 155796 254084 155848
rect 324412 155796 324464 155848
rect 328552 155796 328604 155848
rect 252468 155728 252520 155780
rect 269120 155728 269172 155780
rect 295984 154640 296036 154692
rect 307668 154640 307720 154692
rect 261484 154572 261536 154624
rect 307484 154572 307536 154624
rect 251640 154504 251692 154556
rect 270592 154504 270644 154556
rect 324320 154504 324372 154556
rect 346676 154504 346728 154556
rect 283748 153348 283800 153400
rect 307576 153348 307628 153400
rect 184204 153280 184256 153332
rect 214012 153280 214064 153332
rect 263048 153280 263100 153332
rect 307668 153280 307720 153332
rect 324320 153280 324372 153332
rect 327356 153280 327408 153332
rect 171876 153212 171928 153264
rect 213920 153212 213972 153264
rect 255964 153212 256016 153264
rect 307484 153212 307536 153264
rect 251916 153144 251968 153196
rect 281632 153144 281684 153196
rect 252376 153076 252428 153128
rect 271972 153076 272024 153128
rect 252468 153008 252520 153060
rect 269212 153008 269264 153060
rect 258908 152464 258960 152516
rect 306564 152464 306616 152516
rect 203616 151852 203668 151904
rect 213920 151852 213972 151904
rect 300768 151852 300820 151904
rect 307576 151852 307628 151904
rect 191104 151784 191156 151836
rect 214012 151784 214064 151836
rect 253480 151784 253532 151836
rect 307668 151784 307720 151836
rect 251916 151716 251968 151768
rect 276020 151716 276072 151768
rect 324320 151716 324372 151768
rect 346584 151716 346636 151768
rect 252376 151648 252428 151700
rect 274824 151648 274876 151700
rect 252468 151580 252520 151632
rect 267740 151580 267792 151632
rect 177672 151036 177724 151088
rect 210424 151036 210476 151088
rect 298928 150560 298980 150612
rect 307668 150560 307720 150612
rect 211804 150492 211856 150544
rect 214012 150492 214064 150544
rect 268568 150492 268620 150544
rect 307484 150492 307536 150544
rect 207664 150424 207716 150476
rect 213920 150424 213972 150476
rect 254584 150424 254636 150476
rect 306748 150424 306800 150476
rect 206284 150356 206336 150408
rect 214012 150356 214064 150408
rect 251180 150356 251232 150408
rect 254124 150356 254176 150408
rect 324320 150356 324372 150408
rect 330024 150356 330076 150408
rect 210516 150288 210568 150340
rect 213920 150288 213972 150340
rect 252008 150288 252060 150340
rect 273352 150288 273404 150340
rect 252468 150220 252520 150272
rect 274732 150220 274784 150272
rect 296076 149676 296128 149728
rect 307116 149676 307168 149728
rect 300308 149200 300360 149252
rect 306748 149200 306800 149252
rect 301780 149132 301832 149184
rect 307668 149132 307720 149184
rect 253204 149064 253256 149116
rect 307576 149064 307628 149116
rect 187056 148996 187108 149048
rect 213920 148996 213972 149048
rect 252468 148996 252520 149048
rect 266452 148996 266504 149048
rect 324320 148928 324372 148980
rect 349436 148928 349488 148980
rect 251916 148860 251968 148912
rect 255412 148860 255464 148912
rect 324412 148792 324464 148844
rect 325976 148792 326028 148844
rect 252284 148588 252336 148640
rect 259460 148588 259512 148640
rect 269764 147704 269816 147756
rect 307576 147704 307628 147756
rect 198096 147636 198148 147688
rect 213920 147636 213972 147688
rect 254768 147636 254820 147688
rect 307668 147636 307720 147688
rect 252468 147568 252520 147620
rect 277400 147568 277452 147620
rect 324320 147568 324372 147620
rect 343824 147568 343876 147620
rect 252376 147500 252428 147552
rect 276112 147500 276164 147552
rect 251916 146888 251968 146940
rect 273904 146888 273956 146940
rect 276756 146888 276808 146940
rect 307392 146888 307444 146940
rect 304356 146412 304408 146464
rect 307668 146412 307720 146464
rect 182824 146344 182876 146396
rect 213920 146344 213972 146396
rect 274180 146344 274232 146396
rect 307576 146344 307628 146396
rect 167644 146276 167696 146328
rect 214012 146276 214064 146328
rect 256148 146276 256200 146328
rect 307484 146276 307536 146328
rect 252468 146208 252520 146260
rect 273444 146208 273496 146260
rect 252100 146140 252152 146192
rect 262312 146140 262364 146192
rect 251824 146072 251876 146124
rect 258080 146072 258132 146124
rect 282460 145732 282512 145784
rect 303620 145732 303672 145784
rect 265072 145664 265124 145716
rect 293040 145664 293092 145716
rect 256240 145596 256292 145648
rect 306656 145596 306708 145648
rect 196808 145528 196860 145580
rect 214380 145528 214432 145580
rect 253388 145528 253440 145580
rect 307300 145528 307352 145580
rect 252284 145460 252336 145512
rect 256976 145460 257028 145512
rect 193956 144984 194008 145036
rect 213920 144984 213972 145036
rect 304448 144984 304500 145036
rect 307668 144984 307720 145036
rect 171968 144916 172020 144968
rect 214012 144916 214064 144968
rect 293408 144916 293460 144968
rect 307484 144916 307536 144968
rect 252100 144848 252152 144900
rect 264980 144848 265032 144900
rect 324320 144848 324372 144900
rect 342444 144848 342496 144900
rect 252468 144780 252520 144832
rect 260840 144780 260892 144832
rect 204996 143624 205048 143676
rect 214012 143624 214064 143676
rect 188344 143556 188396 143608
rect 213920 143556 213972 143608
rect 274088 143556 274140 143608
rect 307668 143556 307720 143608
rect 323584 143488 323636 143540
rect 324504 143488 324556 143540
rect 324596 143488 324648 143540
rect 343732 143488 343784 143540
rect 324320 143420 324372 143472
rect 336924 143420 336976 143472
rect 250628 142808 250680 142860
rect 305092 142808 305144 142860
rect 256056 142264 256108 142316
rect 307668 142264 307720 142316
rect 272616 142196 272668 142248
rect 307576 142196 307628 142248
rect 195244 142128 195296 142180
rect 213920 142128 213972 142180
rect 324596 142060 324648 142112
rect 345204 142060 345256 142112
rect 324320 141992 324372 142044
rect 336740 141992 336792 142044
rect 171784 141380 171836 141432
rect 209044 141380 209096 141432
rect 253296 141380 253348 141432
rect 307024 141380 307076 141432
rect 210516 140836 210568 140888
rect 214012 140836 214064 140888
rect 280988 140836 281040 140888
rect 306932 140836 306984 140888
rect 206284 140768 206336 140820
rect 213920 140768 213972 140820
rect 252100 140700 252152 140752
rect 281540 140700 281592 140752
rect 324320 140700 324372 140752
rect 338304 140700 338356 140752
rect 177764 140020 177816 140072
rect 216036 140020 216088 140072
rect 252284 139816 252336 139868
rect 260380 139816 260432 139868
rect 286324 139544 286376 139596
rect 307668 139544 307720 139596
rect 271144 139476 271196 139528
rect 307576 139476 307628 139528
rect 206376 139408 206428 139460
rect 213920 139408 213972 139460
rect 260288 139408 260340 139460
rect 307484 139408 307536 139460
rect 324320 139340 324372 139392
rect 339684 139340 339736 139392
rect 472624 139340 472676 139392
rect 580172 139340 580224 139392
rect 287888 138116 287940 138168
rect 307668 138116 307720 138168
rect 170496 138048 170548 138100
rect 213920 138048 213972 138100
rect 261576 138048 261628 138100
rect 307576 138048 307628 138100
rect 166264 137980 166316 138032
rect 214012 137980 214064 138032
rect 250444 137980 250496 138032
rect 307484 137980 307536 138032
rect 252376 137912 252428 137964
rect 278872 137912 278924 137964
rect 324412 137912 324464 137964
rect 343916 137912 343968 137964
rect 252100 137844 252152 137896
rect 273260 137844 273312 137896
rect 324320 137844 324372 137896
rect 335544 137844 335596 137896
rect 252468 137776 252520 137828
rect 267832 137776 267884 137828
rect 167736 137232 167788 137284
rect 211804 137232 211856 137284
rect 252192 137096 252244 137148
rect 259092 137096 259144 137148
rect 280896 136756 280948 136808
rect 307576 136756 307628 136808
rect 258816 136688 258868 136740
rect 306564 136688 306616 136740
rect 177304 136620 177356 136672
rect 213920 136620 213972 136672
rect 249064 136620 249116 136672
rect 307668 136620 307720 136672
rect 252376 136552 252428 136604
rect 288072 136552 288124 136604
rect 324412 136552 324464 136604
rect 341064 136552 341116 136604
rect 252100 136484 252152 136536
rect 282276 136484 282328 136536
rect 252468 136416 252520 136468
rect 264428 136416 264480 136468
rect 324320 136348 324372 136400
rect 327264 136348 327316 136400
rect 251916 135872 251968 135924
rect 290464 135872 290516 135924
rect 282368 135464 282420 135516
rect 307484 135464 307536 135516
rect 297456 135396 297508 135448
rect 307668 135396 307720 135448
rect 193864 135328 193916 135380
rect 214012 135328 214064 135380
rect 290556 135328 290608 135380
rect 307576 135328 307628 135380
rect 169024 135260 169076 135312
rect 213920 135260 213972 135312
rect 304264 135260 304316 135312
rect 307668 135260 307720 135312
rect 251640 135192 251692 135244
rect 294604 135192 294656 135244
rect 252468 135124 252520 135176
rect 269856 135124 269908 135176
rect 294696 134036 294748 134088
rect 307668 134036 307720 134088
rect 289360 133968 289412 134020
rect 307484 133968 307536 134020
rect 189816 133900 189868 133952
rect 213920 133900 213972 133952
rect 270040 133900 270092 133952
rect 307576 133900 307628 133952
rect 251456 133832 251508 133884
rect 280804 133832 280856 133884
rect 252468 133764 252520 133816
rect 271236 133764 271288 133816
rect 252008 133696 252060 133748
rect 261668 133696 261720 133748
rect 271420 133152 271472 133204
rect 307116 133152 307168 133204
rect 302976 132608 303028 132660
rect 307576 132608 307628 132660
rect 293224 132540 293276 132592
rect 307668 132540 307720 132592
rect 173256 132472 173308 132524
rect 213920 132472 213972 132524
rect 282276 132472 282328 132524
rect 307392 132472 307444 132524
rect 252468 132404 252520 132456
rect 265624 132404 265676 132456
rect 324320 132404 324372 132456
rect 347872 132404 347924 132456
rect 251548 132132 251600 132184
rect 254860 132132 254912 132184
rect 202236 131112 202288 131164
rect 213920 131112 213972 131164
rect 267004 131112 267056 131164
rect 307668 131112 307720 131164
rect 252468 131044 252520 131096
rect 271328 131044 271380 131096
rect 324320 131044 324372 131096
rect 350632 131044 350684 131096
rect 251548 130976 251600 131028
rect 267096 130976 267148 131028
rect 324412 130976 324464 131028
rect 328736 130976 328788 131028
rect 183008 130364 183060 130416
rect 214748 130364 214800 130416
rect 283656 129888 283708 129940
rect 307668 129888 307720 129940
rect 273904 129820 273956 129872
rect 307576 129820 307628 129872
rect 171784 129752 171836 129804
rect 213920 129752 213972 129804
rect 268476 129752 268528 129804
rect 306748 129752 306800 129804
rect 251732 129684 251784 129736
rect 283564 129684 283616 129736
rect 324320 129684 324372 129736
rect 351920 129684 351972 129736
rect 252008 129616 252060 129668
rect 275284 129616 275336 129668
rect 324412 129616 324464 129668
rect 328644 129616 328696 129668
rect 252468 129548 252520 129600
rect 262864 129548 262916 129600
rect 297364 128460 297416 128512
rect 307668 128460 307720 128512
rect 276664 128392 276716 128444
rect 307392 128392 307444 128444
rect 174544 128324 174596 128376
rect 213920 128324 213972 128376
rect 275376 128324 275428 128376
rect 307576 128324 307628 128376
rect 252376 128256 252428 128308
rect 291936 128256 291988 128308
rect 324320 128256 324372 128308
rect 328460 128256 328512 128308
rect 252468 128188 252520 128240
rect 278228 128188 278280 128240
rect 252008 128120 252060 128172
rect 269948 128120 270000 128172
rect 324412 127916 324464 127968
rect 327172 127916 327224 127968
rect 251824 127576 251876 127628
rect 261760 127576 261812 127628
rect 279516 127100 279568 127152
rect 307116 127100 307168 127152
rect 188436 127032 188488 127084
rect 213920 127032 213972 127084
rect 278136 127032 278188 127084
rect 307668 127032 307720 127084
rect 170404 126964 170456 127016
rect 214012 126964 214064 127016
rect 269856 126964 269908 127016
rect 306748 126964 306800 127016
rect 252192 126896 252244 126948
rect 278320 126896 278372 126948
rect 449164 126896 449216 126948
rect 580172 126896 580224 126948
rect 252468 126692 252520 126744
rect 257436 126692 257488 126744
rect 251272 126216 251324 126268
rect 300124 126216 300176 126268
rect 211896 125672 211948 125724
rect 214472 125672 214524 125724
rect 290464 125672 290516 125724
rect 307668 125672 307720 125724
rect 166448 125604 166500 125656
rect 213920 125604 213972 125656
rect 271328 125604 271380 125656
rect 306748 125604 306800 125656
rect 252192 125536 252244 125588
rect 287796 125536 287848 125588
rect 324320 125536 324372 125588
rect 342352 125536 342404 125588
rect 251180 125332 251232 125384
rect 253296 125332 253348 125384
rect 252100 124856 252152 124908
rect 265716 124856 265768 124908
rect 301504 124380 301556 124432
rect 307668 124380 307720 124432
rect 287704 124312 287756 124364
rect 306748 124312 306800 124364
rect 180064 124244 180116 124296
rect 214012 124244 214064 124296
rect 265624 124244 265676 124296
rect 307116 124244 307168 124296
rect 166356 124176 166408 124228
rect 213920 124176 213972 124228
rect 260380 124176 260432 124228
rect 307576 124176 307628 124228
rect 252468 124108 252520 124160
rect 272524 124108 272576 124160
rect 324320 124108 324372 124160
rect 340972 124108 341024 124160
rect 252008 123428 252060 123480
rect 283748 123428 283800 123480
rect 211988 123360 212040 123412
rect 214012 123360 214064 123412
rect 289176 122952 289228 123004
rect 306564 122952 306616 123004
rect 283564 122884 283616 122936
rect 307668 122884 307720 122936
rect 185584 122816 185636 122868
rect 213920 122816 213972 122868
rect 252284 122816 252336 122868
rect 258724 122816 258776 122868
rect 275284 122816 275336 122868
rect 307576 122816 307628 122868
rect 252468 122748 252520 122800
rect 289268 122748 289320 122800
rect 324320 122748 324372 122800
rect 349344 122748 349396 122800
rect 252376 122680 252428 122732
rect 279608 122680 279660 122732
rect 291936 121592 291988 121644
rect 307576 121592 307628 121644
rect 186964 121524 187016 121576
rect 213920 121524 213972 121576
rect 252468 121524 252520 121576
rect 260104 121524 260156 121576
rect 284944 121524 284996 121576
rect 307668 121524 307720 121576
rect 178776 121456 178828 121508
rect 214012 121456 214064 121508
rect 278228 121456 278280 121508
rect 306748 121456 306800 121508
rect 251916 121388 251968 121440
rect 303068 121388 303120 121440
rect 324412 121388 324464 121440
rect 345020 121388 345072 121440
rect 252468 121320 252520 121372
rect 276848 121320 276900 121372
rect 324320 121320 324372 121372
rect 330116 121320 330168 121372
rect 252100 121252 252152 121304
rect 258908 121252 258960 121304
rect 302884 120232 302936 120284
rect 306748 120232 306800 120284
rect 196716 120164 196768 120216
rect 214012 120164 214064 120216
rect 280804 120164 280856 120216
rect 307576 120164 307628 120216
rect 169116 120096 169168 120148
rect 213920 120096 213972 120148
rect 273996 120096 274048 120148
rect 307668 120096 307720 120148
rect 252376 120028 252428 120080
rect 296076 120028 296128 120080
rect 324320 120028 324372 120080
rect 338212 120028 338264 120080
rect 252468 119960 252520 120012
rect 264336 119960 264388 120012
rect 261760 119348 261812 119400
rect 307484 119348 307536 119400
rect 192576 118804 192628 118856
rect 213920 118804 213972 118856
rect 173348 118736 173400 118788
rect 214012 118736 214064 118788
rect 296168 118736 296220 118788
rect 307668 118736 307720 118788
rect 167828 118668 167880 118720
rect 214104 118668 214156 118720
rect 252468 118668 252520 118720
rect 260196 118668 260248 118720
rect 294604 118668 294656 118720
rect 306748 118668 306800 118720
rect 252100 118600 252152 118652
rect 287980 118600 288032 118652
rect 324320 118600 324372 118652
rect 336832 118600 336884 118652
rect 324412 118532 324464 118584
rect 334072 118532 334124 118584
rect 251548 118396 251600 118448
rect 257344 118396 257396 118448
rect 251824 117920 251876 117972
rect 304356 117920 304408 117972
rect 203708 117376 203760 117428
rect 214012 117376 214064 117428
rect 301688 117376 301740 117428
rect 307668 117376 307720 117428
rect 167920 117308 167972 117360
rect 213920 117308 213972 117360
rect 287796 117308 287848 117360
rect 307484 117308 307536 117360
rect 252376 117240 252428 117292
rect 285128 117240 285180 117292
rect 324320 117240 324372 117292
rect 343640 117240 343692 117292
rect 324412 117172 324464 117224
rect 335452 117172 335504 117224
rect 251548 116900 251600 116952
rect 257528 116900 257580 116952
rect 251916 116560 251968 116612
rect 263048 116560 263100 116612
rect 296076 116560 296128 116612
rect 307208 116560 307260 116612
rect 189908 116016 189960 116068
rect 214012 116016 214064 116068
rect 285036 116016 285088 116068
rect 307484 116016 307536 116068
rect 187056 115948 187108 116000
rect 213920 115948 213972 116000
rect 262864 115948 262916 116000
rect 307668 115948 307720 116000
rect 252376 115880 252428 115932
rect 295984 115880 296036 115932
rect 324320 115880 324372 115932
rect 345112 115880 345164 115932
rect 251640 115812 251692 115864
rect 254676 115812 254728 115864
rect 298836 114656 298888 114708
rect 307576 114656 307628 114708
rect 185676 114588 185728 114640
rect 213920 114588 213972 114640
rect 287980 114588 288032 114640
rect 307668 114588 307720 114640
rect 182916 114520 182968 114572
rect 214012 114520 214064 114572
rect 253296 114520 253348 114572
rect 307484 114520 307536 114572
rect 252468 114452 252520 114504
rect 261484 114452 261536 114504
rect 324412 114452 324464 114504
rect 332692 114452 332744 114504
rect 324320 114384 324372 114436
rect 331220 114384 331272 114436
rect 252468 113704 252520 113756
rect 259000 113704 259052 113756
rect 251732 113364 251784 113416
rect 253480 113364 253532 113416
rect 181444 113228 181496 113280
rect 214012 113228 214064 113280
rect 264336 113228 264388 113280
rect 307576 113228 307628 113280
rect 172060 113160 172112 113212
rect 213920 113160 213972 113212
rect 260104 113160 260156 113212
rect 307668 113160 307720 113212
rect 252100 113092 252152 113144
rect 296076 113092 296128 113144
rect 324320 113092 324372 113144
rect 338120 113092 338172 113144
rect 468484 113092 468536 113144
rect 579804 113092 579856 113144
rect 252192 113024 252244 113076
rect 255964 113024 256016 113076
rect 174636 112412 174688 112464
rect 214932 112412 214984 112464
rect 252008 112412 252060 112464
rect 304448 112412 304500 112464
rect 303068 111936 303120 111988
rect 307300 111936 307352 111988
rect 167552 111868 167604 111920
rect 167736 111868 167788 111920
rect 304356 111868 304408 111920
rect 307668 111868 307720 111920
rect 177396 111800 177448 111852
rect 213920 111800 213972 111852
rect 293316 111800 293368 111852
rect 306564 111800 306616 111852
rect 167736 111732 167788 111784
rect 207664 111732 207716 111784
rect 252376 111732 252428 111784
rect 256240 111732 256292 111784
rect 324320 111732 324372 111784
rect 339500 111732 339552 111784
rect 252284 111188 252336 111240
rect 274180 111188 274232 111240
rect 256608 111120 256660 111172
rect 282460 111120 282512 111172
rect 251916 111052 251968 111104
rect 301780 111052 301832 111104
rect 300124 110576 300176 110628
rect 306564 110576 306616 110628
rect 192668 110508 192720 110560
rect 214012 110508 214064 110560
rect 295984 110508 296036 110560
rect 307300 110508 307352 110560
rect 169208 110440 169260 110492
rect 213920 110440 213972 110492
rect 283748 110440 283800 110492
rect 306748 110440 306800 110492
rect 251456 110372 251508 110424
rect 254584 110372 254636 110424
rect 324320 110372 324372 110424
rect 332600 110372 332652 110424
rect 251548 110304 251600 110356
rect 268568 110304 268620 110356
rect 252468 110236 252520 110288
rect 298928 110236 298980 110288
rect 303160 109148 303212 109200
rect 306748 109148 306800 109200
rect 296076 109080 296128 109132
rect 307668 109080 307720 109132
rect 170588 109012 170640 109064
rect 213920 109012 213972 109064
rect 272524 109012 272576 109064
rect 307576 109012 307628 109064
rect 167736 108944 167788 108996
rect 196808 108944 196860 108996
rect 251824 108944 251876 108996
rect 300308 108944 300360 108996
rect 251180 108876 251232 108928
rect 253204 108876 253256 108928
rect 324320 108876 324372 108928
rect 339592 108876 339644 108928
rect 252560 108264 252612 108316
rect 291844 108264 291896 108316
rect 255964 107856 256016 107908
rect 307668 107856 307720 107908
rect 207664 107720 207716 107772
rect 214012 107720 214064 107772
rect 300216 107720 300268 107772
rect 307300 107720 307352 107772
rect 199384 107652 199436 107704
rect 213920 107652 213972 107704
rect 301780 107652 301832 107704
rect 307484 107652 307536 107704
rect 252376 107584 252428 107636
rect 276756 107584 276808 107636
rect 252468 107516 252520 107568
rect 269764 107516 269816 107568
rect 251548 107380 251600 107432
rect 254768 107380 254820 107432
rect 292028 106972 292080 107024
rect 307208 106972 307260 107024
rect 276112 106904 276164 106956
rect 295340 106904 295392 106956
rect 304448 106428 304500 106480
rect 307668 106428 307720 106480
rect 211804 106360 211856 106412
rect 214472 106360 214524 106412
rect 298928 106360 298980 106412
rect 307484 106360 307536 106412
rect 167736 106292 167788 106344
rect 213920 106292 213972 106344
rect 261484 106292 261536 106344
rect 307300 106292 307352 106344
rect 324320 106224 324372 106276
rect 347780 106224 347832 106276
rect 251180 106156 251232 106208
rect 253388 106156 253440 106208
rect 252376 105680 252428 105732
rect 256148 105680 256200 105732
rect 252192 105612 252244 105664
rect 306012 105612 306064 105664
rect 251640 105544 251692 105596
rect 306104 105544 306156 105596
rect 293500 105000 293552 105052
rect 307668 105000 307720 105052
rect 196900 104932 196952 104984
rect 213920 104932 213972 104984
rect 194048 104864 194100 104916
rect 214012 104864 214064 104916
rect 252468 104796 252520 104848
rect 293408 104796 293460 104848
rect 324320 104796 324372 104848
rect 356060 104796 356112 104848
rect 324320 104660 324372 104712
rect 327080 104660 327132 104712
rect 252284 104116 252336 104168
rect 305736 104116 305788 104168
rect 304540 103640 304592 103692
rect 307668 103640 307720 103692
rect 202328 103572 202380 103624
rect 213920 103572 213972 103624
rect 296260 103572 296312 103624
rect 307484 103572 307536 103624
rect 199476 103504 199528 103556
rect 214012 103504 214064 103556
rect 278320 103504 278372 103556
rect 307576 103504 307628 103556
rect 252376 103436 252428 103488
rect 274088 103436 274140 103488
rect 252468 103368 252520 103420
rect 271420 103368 271472 103420
rect 299020 102280 299072 102332
rect 306564 102280 306616 102332
rect 207756 102212 207808 102264
rect 214012 102212 214064 102264
rect 274180 102212 274232 102264
rect 307576 102212 307628 102264
rect 191196 102144 191248 102196
rect 213920 102144 213972 102196
rect 271236 102144 271288 102196
rect 307668 102144 307720 102196
rect 252468 102076 252520 102128
rect 272616 102076 272668 102128
rect 252008 101192 252060 101244
rect 256056 101192 256108 101244
rect 254584 100920 254636 100972
rect 307668 100920 307720 100972
rect 297548 100852 297600 100904
rect 306564 100852 306616 100904
rect 260196 100784 260248 100836
rect 307668 100784 307720 100836
rect 206468 100716 206520 100768
rect 213920 100716 213972 100768
rect 252100 100648 252152 100700
rect 292028 100648 292080 100700
rect 467104 100648 467156 100700
rect 580172 100648 580224 100700
rect 252468 100580 252520 100632
rect 280988 100580 281040 100632
rect 170680 99968 170732 100020
rect 214656 99968 214708 100020
rect 294788 99492 294840 99544
rect 306564 99492 306616 99544
rect 291844 99424 291896 99476
rect 306748 99424 306800 99476
rect 198188 99356 198240 99408
rect 213920 99356 213972 99408
rect 258724 99356 258776 99408
rect 307668 99356 307720 99408
rect 252468 99288 252520 99340
rect 262956 99288 263008 99340
rect 252376 99220 252428 99272
rect 261760 99220 261812 99272
rect 252468 98132 252520 98184
rect 260288 98132 260340 98184
rect 196808 98064 196860 98116
rect 213920 98064 213972 98116
rect 269764 98064 269816 98116
rect 306748 98064 306800 98116
rect 166540 97996 166592 98048
rect 214012 97996 214064 98048
rect 261668 97996 261720 98048
rect 307668 97996 307720 98048
rect 169300 97248 169352 97300
rect 214564 97248 214616 97300
rect 289268 96772 289320 96824
rect 307668 96772 307720 96824
rect 253204 96704 253256 96756
rect 307576 96704 307628 96756
rect 207848 96636 207900 96688
rect 213920 96636 213972 96688
rect 250536 96636 250588 96688
rect 307668 96636 307720 96688
rect 165528 95888 165580 95940
rect 214104 95888 214156 95940
rect 251824 95208 251876 95260
rect 306932 95208 306984 95260
rect 178684 95140 178736 95192
rect 321468 95140 321520 95192
rect 59268 95004 59320 95056
rect 199476 95004 199528 95056
rect 246948 94460 247000 94512
rect 299572 94460 299624 94512
rect 133144 94052 133196 94104
rect 182824 94052 182876 94104
rect 113732 93984 113784 94036
rect 173348 93984 173400 94036
rect 115480 93916 115532 93968
rect 177304 93916 177356 93968
rect 102048 93848 102100 93900
rect 171784 93848 171836 93900
rect 62028 93780 62080 93832
rect 207756 93780 207808 93832
rect 209044 93780 209096 93832
rect 321652 93780 321704 93832
rect 151728 93372 151780 93424
rect 171876 93372 171928 93424
rect 134432 93304 134484 93356
rect 167644 93304 167696 93356
rect 118056 93236 118108 93288
rect 170496 93236 170548 93288
rect 110144 93168 110196 93220
rect 167920 93168 167972 93220
rect 119528 93100 119580 93152
rect 178776 93100 178828 93152
rect 238760 93100 238812 93152
rect 250628 93100 250680 93152
rect 88984 92420 89036 92472
rect 165528 92420 165580 92472
rect 173164 92420 173216 92472
rect 324596 92420 324648 92472
rect 130752 92352 130804 92404
rect 193956 92352 194008 92404
rect 125876 92284 125928 92336
rect 183008 92284 183060 92336
rect 116768 92216 116820 92268
rect 170680 92216 170732 92268
rect 151544 92148 151596 92200
rect 203616 92148 203668 92200
rect 119712 92080 119764 92132
rect 166264 92080 166316 92132
rect 3148 91740 3200 91792
rect 25504 91740 25556 91792
rect 228364 91740 228416 91792
rect 278320 91740 278372 91792
rect 88064 91196 88116 91248
rect 111064 91196 111116 91248
rect 74816 91128 74868 91180
rect 100024 91128 100076 91180
rect 100576 91128 100628 91180
rect 116584 91128 116636 91180
rect 85764 91060 85816 91112
rect 129004 91060 129056 91112
rect 128176 90992 128228 91044
rect 188344 90992 188396 91044
rect 112168 90924 112220 90976
rect 169024 90924 169076 90976
rect 115480 90856 115532 90908
rect 167828 90856 167880 90908
rect 126520 90788 126572 90840
rect 166448 90788 166500 90840
rect 152924 90720 152976 90772
rect 191104 90720 191156 90772
rect 151360 90652 151412 90704
rect 184204 90652 184256 90704
rect 256056 90312 256108 90364
rect 266360 90312 266412 90364
rect 67456 89632 67508 89684
rect 214840 89632 214892 89684
rect 66076 89564 66128 89616
rect 207848 89564 207900 89616
rect 109224 89496 109276 89548
rect 189908 89496 189960 89548
rect 101864 89428 101916 89480
rect 177396 89428 177448 89480
rect 122840 89360 122892 89412
rect 166356 89360 166408 89412
rect 132224 89292 132276 89344
rect 171968 89292 172020 89344
rect 224224 89156 224276 89208
rect 260380 89156 260432 89208
rect 242900 89088 242952 89140
rect 296720 89088 296772 89140
rect 176384 89020 176436 89072
rect 245660 89020 245712 89072
rect 204904 88952 204956 89004
rect 378784 88952 378836 89004
rect 39948 88272 40000 88324
rect 323032 88272 323084 88324
rect 111432 88204 111484 88256
rect 203708 88204 203760 88256
rect 100484 88136 100536 88188
rect 192668 88136 192720 88188
rect 136456 88068 136508 88120
rect 198096 88068 198148 88120
rect 124036 88000 124088 88052
rect 180064 88000 180116 88052
rect 203616 87592 203668 87644
rect 307116 87592 307168 87644
rect 67732 86912 67784 86964
rect 214656 86912 214708 86964
rect 122104 86844 122156 86896
rect 206376 86844 206428 86896
rect 107844 86776 107896 86828
rect 187056 86776 187108 86828
rect 118240 86708 118292 86760
rect 186964 86708 187016 86760
rect 238024 86300 238076 86352
rect 251272 86300 251324 86352
rect 216588 86232 216640 86284
rect 310520 86232 310572 86284
rect 104624 85484 104676 85536
rect 202236 85484 202288 85536
rect 120448 85416 120500 85468
rect 213184 85416 213236 85468
rect 105728 85348 105780 85400
rect 185676 85348 185728 85400
rect 104348 85280 104400 85332
rect 181444 85280 181496 85332
rect 97264 85212 97316 85264
rect 170588 85212 170640 85264
rect 115848 85144 115900 85196
rect 169116 85144 169168 85196
rect 308496 84804 308548 84856
rect 317420 84804 317472 84856
rect 92388 84124 92440 84176
rect 211804 84124 211856 84176
rect 99104 84056 99156 84108
rect 169208 84056 169260 84108
rect 103428 83988 103480 84040
rect 172060 83988 172112 84040
rect 126796 83920 126848 83972
rect 195244 83920 195296 83972
rect 121368 83852 121420 83904
rect 185584 83852 185636 83904
rect 258080 83512 258132 83564
rect 284300 83512 284352 83564
rect 309876 83512 309928 83564
rect 324320 83512 324372 83564
rect 207020 83444 207072 83496
rect 319444 83444 319496 83496
rect 50988 82764 51040 82816
rect 321560 82764 321612 82816
rect 124128 82696 124180 82748
rect 210516 82696 210568 82748
rect 110328 82628 110380 82680
rect 189816 82628 189868 82680
rect 113088 82560 113140 82612
rect 192576 82560 192628 82612
rect 108948 82492 109000 82544
rect 173256 82492 173308 82544
rect 251272 82084 251324 82136
rect 293960 82084 294012 82136
rect 95056 81336 95108 81388
rect 199384 81336 199436 81388
rect 86868 81268 86920 81320
rect 166540 81268 166592 81320
rect 117228 81200 117280 81252
rect 196716 81200 196768 81252
rect 114468 81132 114520 81184
rect 193864 81132 193916 81184
rect 129648 81064 129700 81116
rect 204996 81064 205048 81116
rect 177856 80724 177908 80776
rect 247684 80724 247736 80776
rect 198740 80656 198792 80708
rect 269948 80656 270000 80708
rect 298744 80656 298796 80708
rect 322940 80656 322992 80708
rect 95148 79976 95200 80028
rect 207664 79976 207716 80028
rect 116584 79908 116636 79960
rect 214748 79908 214800 79960
rect 122748 79840 122800 79892
rect 211988 79840 212040 79892
rect 102048 79772 102100 79824
rect 174544 79772 174596 79824
rect 99196 79704 99248 79756
rect 170404 79704 170456 79756
rect 211804 79296 211856 79348
rect 307300 79296 307352 79348
rect 309692 79296 309744 79348
rect 328460 79296 328512 79348
rect 97908 78616 97960 78668
rect 188436 78616 188488 78668
rect 125508 78548 125560 78600
rect 211896 78548 211948 78600
rect 125416 78480 125468 78532
rect 206284 78480 206336 78532
rect 100024 77188 100076 77240
rect 214564 77188 214616 77240
rect 93768 77120 93820 77172
rect 167736 77120 167788 77172
rect 129004 77052 129056 77104
rect 196808 77052 196860 77104
rect 184940 76576 184992 76628
rect 315304 76576 315356 76628
rect 73160 76508 73212 76560
rect 296168 76508 296220 76560
rect 63408 75828 63460 75880
rect 191196 75828 191248 75880
rect 107568 75760 107620 75812
rect 182916 75760 182968 75812
rect 77300 75216 77352 75268
rect 270040 75216 270092 75268
rect 103520 75148 103572 75200
rect 303160 75148 303212 75200
rect 91008 74468 91060 74520
rect 194048 74468 194100 74520
rect 81440 73856 81492 73908
rect 294696 73856 294748 73908
rect 46940 73788 46992 73840
rect 274180 73788 274232 73840
rect 85488 73108 85540 73160
rect 206468 73108 206520 73160
rect 418804 73108 418856 73160
rect 580172 73108 580224 73160
rect 111064 73040 111116 73092
rect 198188 73040 198240 73092
rect 85580 72428 85632 72480
rect 289360 72428 289412 72480
rect 88340 71068 88392 71120
rect 304264 71068 304316 71120
rect 64880 71000 64932 71052
rect 293500 71000 293552 71052
rect 92480 69708 92532 69760
rect 297456 69708 297508 69760
rect 53840 69640 53892 69692
rect 304540 69640 304592 69692
rect 95240 68348 95292 68400
rect 290556 68348 290608 68400
rect 57980 68280 58032 68332
rect 296260 68280 296312 68332
rect 99380 66920 99432 66972
rect 282368 66920 282420 66972
rect 69020 66852 69072 66904
rect 305920 66852 305972 66904
rect 177948 65628 178000 65680
rect 282368 65628 282420 65680
rect 106280 65560 106332 65612
rect 258816 65560 258868 65612
rect 71780 65492 71832 65544
rect 304448 65492 304500 65544
rect 110420 64200 110472 64252
rect 280896 64200 280948 64252
rect 24860 64132 24912 64184
rect 307208 64132 307260 64184
rect 82820 62772 82872 62824
rect 300216 62772 300268 62824
rect 114560 61412 114612 61464
rect 283748 61412 283800 61464
rect 13820 61344 13872 61396
rect 271328 61344 271380 61396
rect 353944 60664 353996 60716
rect 580172 60664 580224 60716
rect 74540 60052 74592 60104
rect 282276 60052 282328 60104
rect 89720 59984 89772 60036
rect 301780 59984 301832 60036
rect 3056 59304 3108 59356
rect 31024 59304 31076 59356
rect 93860 58692 93912 58744
rect 305828 58692 305880 58744
rect 70400 58624 70452 58676
rect 302976 58624 303028 58676
rect 113180 57332 113232 57384
rect 287888 57332 287940 57384
rect 96620 57264 96672 57316
rect 296076 57264 296128 57316
rect 63500 57196 63552 57248
rect 267004 57196 267056 57248
rect 100760 55836 100812 55888
rect 272524 55836 272576 55888
rect 110512 54544 110564 54596
rect 300124 54544 300176 54596
rect 44180 54476 44232 54528
rect 285036 54476 285088 54528
rect 37280 53116 37332 53168
rect 253296 53116 253348 53168
rect 44272 53048 44324 53100
rect 299020 53048 299072 53100
rect 117320 51824 117372 51876
rect 261576 51824 261628 51876
rect 179236 51756 179288 51808
rect 332600 51756 332652 51808
rect 16580 51688 16632 51740
rect 294788 51688 294840 51740
rect 121460 50396 121512 50448
rect 304356 50396 304408 50448
rect 27620 50328 27672 50380
rect 264336 50328 264388 50380
rect 118700 49036 118752 49088
rect 303068 49036 303120 49088
rect 30380 48968 30432 49020
rect 287980 48968 288032 49020
rect 120080 47608 120132 47660
rect 250444 47608 250496 47660
rect 20720 47540 20772 47592
rect 291844 47540 291896 47592
rect 124220 46248 124272 46300
rect 286324 46248 286376 46300
rect 26240 46180 26292 46232
rect 260196 46180 260248 46232
rect 3424 45500 3476 45552
rect 18604 45500 18656 45552
rect 38660 44820 38712 44872
rect 276664 44820 276716 44872
rect 31760 43460 31812 43512
rect 275376 43460 275428 43512
rect 33140 43392 33192 43444
rect 297548 43392 297600 43444
rect 107660 42100 107712 42152
rect 295984 42100 296036 42152
rect 41420 42032 41472 42084
rect 307024 42032 307076 42084
rect 35900 40740 35952 40792
rect 297364 40740 297416 40792
rect 2780 40672 2832 40724
rect 271144 40672 271196 40724
rect 42800 39380 42852 39432
rect 283656 39380 283708 39432
rect 35992 39312 36044 39364
rect 305736 39312 305788 39364
rect 78680 37952 78732 38004
rect 298928 37952 298980 38004
rect 19340 37884 19392 37936
rect 269856 37884 269908 37936
rect 60740 36592 60792 36644
rect 305644 36592 305696 36644
rect 23480 36524 23532 36576
rect 279516 36524 279568 36576
rect 35808 35844 35860 35896
rect 249156 35844 249208 35896
rect 67640 35164 67692 35216
rect 293224 35164 293276 35216
rect 35164 34484 35216 34536
rect 35808 34484 35860 34536
rect 180800 33940 180852 33992
rect 261576 33940 261628 33992
rect 201500 33872 201552 33924
rect 343640 33872 343692 33924
rect 93952 33804 94004 33856
rect 278228 33804 278280 33856
rect 4160 33736 4212 33788
rect 251824 33736 251876 33788
rect 3516 33056 3568 33108
rect 46204 33056 46256 33108
rect 189724 32444 189776 32496
rect 259552 32444 259604 32496
rect 111800 32376 111852 32428
rect 301504 32376 301556 32428
rect 8300 31016 8352 31068
rect 293316 31016 293368 31068
rect 200120 29724 200172 29776
rect 311900 29724 311952 29776
rect 102140 29656 102192 29708
rect 275284 29656 275336 29708
rect 15200 29588 15252 29640
rect 253204 29588 253256 29640
rect 179512 28364 179564 28416
rect 293960 28364 294012 28416
rect 84200 28296 84252 28348
rect 302884 28296 302936 28348
rect 17960 28228 18012 28280
rect 260104 28228 260156 28280
rect 176476 27004 176528 27056
rect 296720 27004 296772 27056
rect 55220 26936 55272 26988
rect 301688 26936 301740 26988
rect 2872 26868 2924 26920
rect 250536 26868 250588 26920
rect 29000 25508 29052 25560
rect 254584 25508 254636 25560
rect 187700 24284 187752 24336
rect 254584 24284 254636 24336
rect 208400 24216 208452 24268
rect 324412 24216 324464 24268
rect 86960 24148 87012 24200
rect 284944 24148 284996 24200
rect 52460 24080 52512 24132
rect 268476 24080 268528 24132
rect 69112 22788 69164 22840
rect 294604 22788 294656 22840
rect 40040 22720 40092 22772
rect 271236 22720 271288 22772
rect 183560 21496 183612 21548
rect 349344 21496 349396 21548
rect 91100 21428 91152 21480
rect 291936 21428 291988 21480
rect 19432 21360 19484 21412
rect 261668 21360 261720 21412
rect 378784 20612 378836 20664
rect 579988 20612 580040 20664
rect 102232 20000 102284 20052
rect 249064 20000 249116 20052
rect 80060 19932 80112 19984
rect 280804 19932 280856 19984
rect 3424 19456 3476 19508
rect 7564 19456 7616 19508
rect 75920 18572 75972 18624
rect 261484 18572 261536 18624
rect 193220 17280 193272 17332
rect 247040 17280 247092 17332
rect 128360 17212 128412 17264
rect 215944 17212 215996 17264
rect 217968 17212 218020 17264
rect 248420 17212 248472 17264
rect 192484 15988 192536 16040
rect 273260 15988 273312 16040
rect 105728 15920 105780 15972
rect 289176 15920 289228 15972
rect 11888 15852 11940 15904
rect 258724 15852 258776 15904
rect 212540 14560 212592 14612
rect 328000 14560 328052 14612
rect 77392 14492 77444 14544
rect 273996 14492 274048 14544
rect 34520 14424 34572 14476
rect 298836 14424 298888 14476
rect 173808 13132 173860 13184
rect 301504 13132 301556 13184
rect 109040 13064 109092 13116
rect 265624 13064 265676 13116
rect 211068 11908 211120 11960
rect 252376 11908 252428 11960
rect 176568 11840 176620 11892
rect 262496 11840 262548 11892
rect 51080 11772 51132 11824
rect 228364 11772 228416 11824
rect 98184 11704 98236 11756
rect 283564 11704 283616 11756
rect 112 10956 164 11008
rect 1308 10956 1360 11008
rect 251180 10956 251232 11008
rect 179420 10344 179472 10396
rect 299664 10344 299716 10396
rect 28448 10276 28500 10328
rect 278136 10276 278188 10328
rect 198004 9052 198056 9104
rect 287796 9052 287848 9104
rect 46664 8984 46716 9036
rect 273904 8984 273956 9036
rect 6460 8916 6512 8968
rect 289268 8916 289320 8968
rect 308404 8916 308456 8968
rect 317328 8916 317380 8968
rect 331864 8236 331916 8288
rect 333888 8236 333940 8288
rect 116400 7624 116452 7676
rect 287704 7624 287756 7676
rect 7656 7556 7708 7608
rect 269764 7556 269816 7608
rect 3424 6808 3476 6860
rect 48964 6808 49016 6860
rect 203524 6332 203576 6384
rect 266544 6332 266596 6384
rect 175188 6264 175240 6316
rect 311440 6264 311492 6316
rect 123484 6196 123536 6248
rect 290464 6196 290516 6248
rect 86868 6128 86920 6180
rect 255964 6128 256016 6180
rect 1676 4768 1728 4820
rect 35164 4768 35216 4820
rect 48964 4768 49016 4820
rect 262864 4768 262916 4820
rect 309784 4768 309836 4820
rect 320916 4768 320968 4820
rect 345664 4156 345716 4208
rect 350448 4156 350500 4208
rect 261576 4088 261628 4140
rect 268844 4088 268896 4140
rect 315304 4088 315356 4140
rect 316224 4088 316276 4140
rect 348056 3952 348108 4004
rect 354680 3952 354732 4004
rect 202144 3680 202196 3732
rect 267740 3680 267792 3732
rect 278044 3680 278096 3732
rect 125876 3612 125928 3664
rect 173900 3612 173952 3664
rect 196624 3612 196676 3664
rect 281908 3612 281960 3664
rect 77300 3544 77352 3596
rect 78220 3544 78272 3596
rect 119896 3544 119948 3596
rect 224224 3544 224276 3596
rect 254584 3544 254636 3596
rect 261760 3544 261812 3596
rect 282184 3544 282236 3596
rect 44180 3476 44232 3528
rect 45100 3476 45152 3528
rect 60832 3476 60884 3528
rect 203616 3476 203668 3528
rect 210424 3476 210476 3528
rect 11152 3408 11204 3460
rect 211804 3408 211856 3460
rect 216036 3408 216088 3460
rect 240508 3408 240560 3460
rect 242900 3476 242952 3528
rect 244096 3476 244148 3528
rect 246948 3476 247000 3528
rect 259460 3476 259512 3528
rect 268384 3476 268436 3528
rect 278320 3476 278372 3528
rect 282368 3476 282420 3528
rect 284300 3476 284352 3528
rect 288992 3544 289044 3596
rect 289084 3544 289136 3596
rect 298468 3544 298520 3596
rect 319444 3544 319496 3596
rect 292580 3476 292632 3528
rect 299480 3476 299532 3528
rect 300768 3476 300820 3528
rect 301596 3476 301648 3528
rect 319720 3476 319772 3528
rect 324412 3544 324464 3596
rect 325608 3544 325660 3596
rect 338672 3544 338724 3596
rect 349160 3544 349212 3596
rect 349344 3544 349396 3596
rect 345756 3476 345808 3528
rect 245200 3408 245252 3460
rect 247684 3408 247736 3460
rect 254676 3408 254728 3460
rect 256608 3408 256660 3460
rect 271236 3408 271288 3460
rect 279424 3408 279476 3460
rect 326804 3408 326856 3460
rect 330392 3408 330444 3460
rect 356704 3408 356756 3460
rect 579804 3408 579856 3460
rect 308588 3340 308640 3392
rect 315028 3340 315080 3392
rect 264244 3272 264296 3324
rect 270040 3272 270092 3324
rect 249984 3204 250036 3256
rect 256056 3204 256108 3256
rect 269948 3000 270000 3052
rect 276020 3000 276072 3052
rect 235816 2932 235868 2984
rect 238024 2932 238076 2984
rect 179328 2116 179380 2168
rect 306748 2116 306800 2168
rect 59636 2048 59688 2100
rect 287888 2048 287940 2100
<< obsm1 >>
rect 68800 95100 164756 174600
<< metal2 >>
rect 6932 703582 7972 703610
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 2778 658200 2834 658209
rect 2778 658135 2834 658144
rect 2792 657014 2820 658135
rect 2780 657008 2832 657014
rect 2780 656950 2832 656956
rect 4804 657008 4856 657014
rect 4804 656950 4856 656956
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3422 606112 3478 606121
rect 3422 606047 3424 606056
rect 3476 606047 3478 606056
rect 3424 606018 3476 606024
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 553450 3464 553823
rect 3424 553444 3476 553450
rect 3424 553386 3476 553392
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 527202 3464 527847
rect 3424 527196 3476 527202
rect 3424 527138 3476 527144
rect 3422 501800 3478 501809
rect 3422 501735 3478 501744
rect 3054 475688 3110 475697
rect 3054 475623 3110 475632
rect 3068 474774 3096 475623
rect 3056 474768 3108 474774
rect 3056 474710 3108 474716
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 2870 410544 2926 410553
rect 2870 410479 2926 410488
rect 2884 409902 2912 410479
rect 2872 409896 2924 409902
rect 2872 409838 2924 409844
rect 3054 358456 3110 358465
rect 3054 358391 3110 358400
rect 3068 357542 3096 358391
rect 3056 357536 3108 357542
rect 3056 357478 3108 357484
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 3436 320890 3464 501735
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3528 462398 3556 462567
rect 3516 462392 3568 462398
rect 3516 462334 3568 462340
rect 3514 423600 3570 423609
rect 3514 423535 3570 423544
rect 3528 422346 3556 423535
rect 3516 422340 3568 422346
rect 3516 422282 3568 422288
rect 3516 397520 3568 397526
rect 3514 397488 3516 397497
rect 3568 397488 3570 397497
rect 3514 397423 3570 397432
rect 3514 371376 3570 371385
rect 3514 371311 3570 371320
rect 3528 371278 3556 371311
rect 3516 371272 3568 371278
rect 3516 371214 3568 371220
rect 3424 320884 3476 320890
rect 3424 320826 3476 320832
rect 3422 319288 3478 319297
rect 3422 319223 3478 319232
rect 3436 318850 3464 319223
rect 3424 318844 3476 318850
rect 3424 318786 3476 318792
rect 4816 311166 4844 656950
rect 6932 347070 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 24320 700330 24348 703520
rect 24308 700324 24360 700330
rect 24308 700266 24360 700272
rect 22744 670744 22796 670750
rect 22744 670686 22796 670692
rect 18604 618316 18656 618322
rect 18604 618258 18656 618264
rect 8944 606076 8996 606082
rect 8944 606018 8996 606024
rect 6920 347064 6972 347070
rect 6920 347006 6972 347012
rect 8956 312594 8984 606018
rect 17224 553444 17276 553450
rect 17224 553386 17276 553392
rect 13084 527196 13136 527202
rect 13084 527138 13136 527144
rect 8944 312588 8996 312594
rect 8944 312530 8996 312536
rect 4804 311160 4856 311166
rect 4804 311102 4856 311108
rect 3238 306232 3294 306241
rect 3238 306167 3294 306176
rect 3252 305046 3280 306167
rect 3240 305040 3292 305046
rect 3240 304982 3292 304988
rect 7564 300892 7616 300898
rect 7564 300834 7616 300840
rect 3424 293276 3476 293282
rect 3424 293218 3476 293224
rect 3330 293176 3386 293185
rect 3330 293111 3386 293120
rect 3344 292874 3372 293111
rect 3332 292868 3384 292874
rect 3332 292810 3384 292816
rect 3054 267200 3110 267209
rect 3054 267135 3110 267144
rect 3068 261526 3096 267135
rect 3056 261520 3108 261526
rect 3056 261462 3108 261468
rect 2778 254144 2834 254153
rect 2778 254079 2780 254088
rect 2832 254079 2834 254088
rect 2780 254050 2832 254056
rect 3330 241088 3386 241097
rect 3330 241023 3386 241032
rect 3344 239426 3372 241023
rect 3332 239420 3384 239426
rect 3332 239362 3384 239368
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3148 189032 3200 189038
rect 3148 188974 3200 188980
rect 3160 188873 3188 188974
rect 3146 188864 3202 188873
rect 3146 188799 3202 188808
rect 1308 177336 1360 177342
rect 1308 177278 1360 177284
rect 1320 11014 1348 177278
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 2780 97776 2832 97782
rect 2780 97718 2832 97724
rect 2792 97617 2820 97718
rect 2778 97608 2834 97617
rect 2778 97543 2834 97552
rect 3148 91792 3200 91798
rect 3148 91734 3200 91740
rect 3160 84697 3188 91734
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 3436 71641 3464 293218
rect 3516 287700 3568 287706
rect 3516 287642 3568 287648
rect 3528 162897 3556 287642
rect 4804 254108 4856 254114
rect 4804 254050 4856 254056
rect 4816 238066 4844 254050
rect 4804 238060 4856 238066
rect 4804 238002 4856 238008
rect 3608 224256 3660 224262
rect 3608 224198 3660 224204
rect 3620 201929 3648 224198
rect 4804 210520 4856 210526
rect 4804 210462 4856 210468
rect 3606 201920 3662 201929
rect 3606 201855 3662 201864
rect 3514 162888 3570 162897
rect 3514 162823 3570 162832
rect 3516 150408 3568 150414
rect 3516 150350 3568 150356
rect 3528 149841 3556 150350
rect 3514 149832 3570 149841
rect 3514 149767 3570 149776
rect 3516 137964 3568 137970
rect 3516 137906 3568 137912
rect 3528 136785 3556 137906
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 4816 97782 4844 210462
rect 4804 97776 4856 97782
rect 4804 97718 4856 97724
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 2780 40724 2832 40730
rect 2780 40666 2832 40672
rect 112 11008 164 11014
rect 112 10950 164 10956
rect 1308 11008 1360 11014
rect 1308 10950 1360 10956
rect 124 354 152 10950
rect 2792 6914 2820 40666
rect 4160 33788 4212 33794
rect 4160 33730 4212 33736
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 2872 26920 2924 26926
rect 2872 26862 2924 26868
rect 2884 16574 2912 26862
rect 3424 19508 3476 19514
rect 3424 19450 3476 19456
rect 3436 19417 3464 19450
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 4172 16574 4200 33730
rect 7576 19514 7604 300834
rect 8944 292868 8996 292874
rect 8944 292810 8996 292816
rect 8956 244254 8984 292810
rect 13096 260846 13124 527138
rect 14464 295452 14516 295458
rect 14464 295394 14516 295400
rect 13084 260840 13136 260846
rect 13084 260782 13136 260788
rect 13084 256760 13136 256766
rect 13084 256702 13136 256708
rect 8944 244248 8996 244254
rect 8944 244190 8996 244196
rect 13096 137970 13124 256702
rect 14476 189038 14504 295394
rect 17236 262886 17264 553386
rect 18616 273970 18644 618258
rect 21364 565888 21416 565894
rect 21364 565830 21416 565836
rect 18604 273964 18656 273970
rect 18604 273906 18656 273912
rect 21376 266393 21404 565830
rect 22756 287026 22784 670686
rect 39304 448588 39356 448594
rect 39304 448530 39356 448536
rect 32404 422340 32456 422346
rect 32404 422282 32456 422288
rect 25504 345092 25556 345098
rect 25504 345034 25556 345040
rect 25516 313954 25544 345034
rect 25504 313948 25556 313954
rect 25504 313890 25556 313896
rect 32416 304978 32444 422282
rect 39316 368966 39344 448530
rect 39304 368960 39356 368966
rect 39304 368902 39356 368908
rect 39948 368960 40000 368966
rect 39948 368902 40000 368908
rect 39960 368558 39988 368902
rect 39948 368552 40000 368558
rect 39948 368494 40000 368500
rect 32404 304972 32456 304978
rect 32404 304914 32456 304920
rect 39960 300150 39988 368494
rect 39948 300144 40000 300150
rect 39948 300086 40000 300092
rect 31024 296812 31076 296818
rect 31024 296754 31076 296760
rect 26884 290488 26936 290494
rect 26884 290430 26936 290436
rect 22744 287020 22796 287026
rect 22744 286962 22796 286968
rect 21362 266384 21418 266393
rect 21362 266319 21418 266328
rect 21364 263628 21416 263634
rect 21364 263570 21416 263576
rect 17224 262880 17276 262886
rect 17224 262822 17276 262828
rect 21376 215286 21404 263570
rect 25504 253224 25556 253230
rect 25504 253166 25556 253172
rect 21364 215280 21416 215286
rect 21364 215222 21416 215228
rect 21364 189848 21416 189854
rect 21364 189790 21416 189796
rect 14464 189032 14516 189038
rect 14464 188974 14516 188980
rect 18604 188420 18656 188426
rect 18604 188362 18656 188368
rect 13084 137964 13136 137970
rect 13084 137906 13136 137912
rect 13820 61396 13872 61402
rect 13820 61338 13872 61344
rect 9678 46200 9734 46209
rect 9678 46135 9734 46144
rect 8300 31068 8352 31074
rect 8300 31010 8352 31016
rect 7564 19508 7616 19514
rect 7564 19450 7616 19456
rect 8312 16574 8340 31010
rect 2884 16546 3648 16574
rect 4172 16546 5304 16574
rect 8312 16546 8800 16574
rect 2792 6886 2912 6914
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1688 480 1716 4762
rect 2884 480 2912 6886
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 542 354 654 480
rect 124 326 654 354
rect 542 -960 654 326
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3620 354 3648 16546
rect 5276 480 5304 16546
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 6472 480 6500 8910
rect 7656 7608 7708 7614
rect 7656 7550 7708 7556
rect 7668 480 7696 7550
rect 8772 480 8800 16546
rect 4038 354 4150 480
rect 3620 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 46135
rect 12438 18592 12494 18601
rect 12438 18527 12494 18536
rect 12452 16574 12480 18527
rect 13832 16574 13860 61338
rect 16580 51740 16632 51746
rect 16580 51682 16632 51688
rect 15200 29640 15252 29646
rect 15200 29582 15252 29588
rect 15212 16574 15240 29582
rect 16592 16574 16620 51682
rect 18616 45558 18644 188362
rect 21376 111790 21404 189790
rect 21364 111784 21416 111790
rect 21364 111726 21416 111732
rect 25516 91798 25544 253166
rect 26896 150414 26924 290430
rect 26884 150408 26936 150414
rect 26884 150350 26936 150356
rect 25504 91792 25556 91798
rect 25504 91734 25556 91740
rect 24860 64184 24912 64190
rect 24860 64126 24912 64132
rect 20720 47592 20772 47598
rect 20720 47534 20772 47540
rect 18604 45552 18656 45558
rect 18604 45494 18656 45500
rect 19340 37936 19392 37942
rect 19340 37878 19392 37884
rect 17960 28280 18012 28286
rect 17960 28222 18012 28228
rect 12452 16546 13584 16574
rect 13832 16546 14320 16574
rect 15212 16546 15976 16574
rect 16592 16546 17080 16574
rect 11888 15904 11940 15910
rect 11888 15846 11940 15852
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11164 480 11192 3402
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 11900 354 11928 15846
rect 13556 480 13584 16546
rect 12318 354 12430 480
rect 11900 326 12430 354
rect 12318 -960 12430 326
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 15948 480 15976 16546
rect 17052 480 17080 16546
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 28222
rect 19352 6914 19380 37878
rect 19432 21412 19484 21418
rect 19432 21354 19484 21360
rect 19444 16574 19472 21354
rect 20732 16574 20760 47534
rect 23480 36576 23532 36582
rect 23480 36518 23532 36524
rect 22098 17232 22154 17241
rect 22098 17167 22154 17176
rect 22112 16574 22140 17167
rect 23492 16574 23520 36518
rect 24872 16574 24900 64126
rect 31036 59362 31064 296754
rect 35806 293992 35862 294001
rect 35806 293927 35862 293936
rect 31024 59356 31076 59362
rect 31024 59298 31076 59304
rect 27620 50380 27672 50386
rect 27620 50322 27672 50328
rect 26240 46232 26292 46238
rect 26240 46174 26292 46180
rect 19444 16546 20208 16574
rect 20732 16546 21864 16574
rect 22112 16546 22600 16574
rect 23492 16546 24256 16574
rect 24872 16546 25360 16574
rect 19352 6886 19472 6914
rect 19444 480 19472 6886
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20180 354 20208 16546
rect 21836 480 21864 16546
rect 20598 354 20710 480
rect 20180 326 20710 354
rect 20598 -960 20710 326
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 24228 480 24256 16546
rect 25332 480 25360 16546
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 46174
rect 27632 16574 27660 50322
rect 30380 49020 30432 49026
rect 30380 48962 30432 48968
rect 29000 25560 29052 25566
rect 29000 25502 29052 25508
rect 29012 16574 29040 25502
rect 30392 16574 30420 48962
rect 31760 43512 31812 43518
rect 31760 43454 31812 43460
rect 31772 16574 31800 43454
rect 33140 43444 33192 43450
rect 33140 43386 33192 43392
rect 33152 16574 33180 43386
rect 35820 35902 35848 293927
rect 39948 285728 40000 285734
rect 39948 285670 40000 285676
rect 39960 88330 39988 285670
rect 40052 236706 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 700398 73016 703520
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 72976 700392 73028 700398
rect 72976 700334 73028 700340
rect 82084 700392 82136 700398
rect 82084 700334 82136 700340
rect 43444 700324 43496 700330
rect 43444 700266 43496 700272
rect 62764 700324 62816 700330
rect 62764 700266 62816 700272
rect 43456 302938 43484 700266
rect 44824 632120 44876 632126
rect 44824 632062 44876 632068
rect 44836 354006 44864 632062
rect 53104 409896 53156 409902
rect 53104 409838 53156 409844
rect 44824 354000 44876 354006
rect 44824 353942 44876 353948
rect 45468 354000 45520 354006
rect 45468 353942 45520 353948
rect 43444 302932 43496 302938
rect 43444 302874 43496 302880
rect 45376 271924 45428 271930
rect 45376 271866 45428 271872
rect 44088 269136 44140 269142
rect 44088 269078 44140 269084
rect 40040 236700 40092 236706
rect 40040 236642 40092 236648
rect 44100 193934 44128 269078
rect 45388 206446 45416 271866
rect 45480 266354 45508 353942
rect 50896 351212 50948 351218
rect 50896 351154 50948 351160
rect 48964 279472 49016 279478
rect 48964 279414 49016 279420
rect 46848 277432 46900 277438
rect 46848 277374 46900 277380
rect 46756 267776 46808 267782
rect 46756 267718 46808 267724
rect 45468 266348 45520 266354
rect 45468 266290 45520 266296
rect 46768 234598 46796 267718
rect 46756 234592 46808 234598
rect 46756 234534 46808 234540
rect 46768 234190 46796 234534
rect 46204 234184 46256 234190
rect 46204 234126 46256 234132
rect 46756 234184 46808 234190
rect 46756 234126 46808 234132
rect 45376 206440 45428 206446
rect 45376 206382 45428 206388
rect 44088 193928 44140 193934
rect 44088 193870 44140 193876
rect 39948 88324 40000 88330
rect 39948 88266 40000 88272
rect 44180 54528 44232 54534
rect 44180 54470 44232 54476
rect 37280 53168 37332 53174
rect 37280 53110 37332 53116
rect 35900 40792 35952 40798
rect 35900 40734 35952 40740
rect 35808 35896 35860 35902
rect 35808 35838 35860 35844
rect 35820 34542 35848 35838
rect 35164 34536 35216 34542
rect 35164 34478 35216 34484
rect 35808 34536 35860 34542
rect 35808 34478 35860 34484
rect 27632 16546 27752 16574
rect 29012 16546 30144 16574
rect 30392 16546 30880 16574
rect 31772 16546 31984 16574
rect 33152 16546 33640 16574
rect 27724 480 27752 16546
rect 28448 10328 28500 10334
rect 28448 10270 28500 10276
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28460 354 28488 10270
rect 30116 480 30144 16546
rect 28878 354 28990 480
rect 28460 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 33612 480 33640 16546
rect 34520 14476 34572 14482
rect 34520 14418 34572 14424
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 14418
rect 35176 4826 35204 34478
rect 35912 6914 35940 40734
rect 35992 39364 36044 39370
rect 35992 39306 36044 39312
rect 36004 16574 36032 39306
rect 37292 16574 37320 53110
rect 38660 44872 38712 44878
rect 38660 44814 38712 44820
rect 38672 16574 38700 44814
rect 41420 42084 41472 42090
rect 41420 42026 41472 42032
rect 40040 22772 40092 22778
rect 40040 22714 40092 22720
rect 40052 16574 40080 22714
rect 41432 16574 41460 42026
rect 42800 39432 42852 39438
rect 42800 39374 42852 39380
rect 36004 16546 36768 16574
rect 37292 16546 38424 16574
rect 38672 16546 39160 16574
rect 40052 16546 40264 16574
rect 41432 16546 41920 16574
rect 35912 6886 36032 6914
rect 35164 4820 35216 4826
rect 35164 4762 35216 4768
rect 36004 480 36032 6886
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 16546
rect 38396 480 38424 16546
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 41892 480 41920 16546
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 42812 354 42840 39374
rect 44192 3534 44220 54470
rect 44272 53100 44324 53106
rect 44272 53042 44324 53048
rect 44180 3528 44232 3534
rect 44180 3470 44232 3476
rect 44284 480 44312 53042
rect 46216 33114 46244 234126
rect 46860 214606 46888 277374
rect 48228 263696 48280 263702
rect 48228 263638 48280 263644
rect 48240 218822 48268 263638
rect 48228 218816 48280 218822
rect 48228 218758 48280 218764
rect 46848 214600 46900 214606
rect 46848 214542 46900 214548
rect 46940 73840 46992 73846
rect 46940 73782 46992 73788
rect 46204 33108 46256 33114
rect 46204 33050 46256 33056
rect 46952 16574 46980 73782
rect 46952 16546 47440 16574
rect 46664 9036 46716 9042
rect 46664 8978 46716 8984
rect 45100 3528 45152 3534
rect 45100 3470 45152 3476
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45112 354 45140 3470
rect 46676 480 46704 8978
rect 45438 354 45550 480
rect 45112 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 48976 6866 49004 279414
rect 50908 253910 50936 351154
rect 52368 287088 52420 287094
rect 52368 287030 52420 287036
rect 50988 270564 51040 270570
rect 50988 270506 51040 270512
rect 50528 253904 50580 253910
rect 50528 253846 50580 253852
rect 50896 253904 50948 253910
rect 50896 253846 50948 253852
rect 50540 253230 50568 253846
rect 50528 253224 50580 253230
rect 50528 253166 50580 253172
rect 50896 252612 50948 252618
rect 50896 252554 50948 252560
rect 50908 196654 50936 252554
rect 50896 196648 50948 196654
rect 50896 196590 50948 196596
rect 51000 82822 51028 270506
rect 52380 210497 52408 287030
rect 53116 244934 53144 409838
rect 58624 397520 58676 397526
rect 58624 397462 58676 397468
rect 55036 357468 55088 357474
rect 55036 357410 55088 357416
rect 53656 289876 53708 289882
rect 53656 289818 53708 289824
rect 53564 264988 53616 264994
rect 53564 264930 53616 264936
rect 53104 244928 53156 244934
rect 53104 244870 53156 244876
rect 53576 211857 53604 264930
rect 53562 211848 53618 211857
rect 53562 211783 53618 211792
rect 52366 210488 52422 210497
rect 52366 210423 52422 210432
rect 53668 207670 53696 289818
rect 54944 280288 54996 280294
rect 54944 280230 54996 280236
rect 53748 276072 53800 276078
rect 53748 276014 53800 276020
rect 53656 207664 53708 207670
rect 53656 207606 53708 207612
rect 53760 180033 53788 276014
rect 53840 262880 53892 262886
rect 53840 262822 53892 262828
rect 53852 262274 53880 262822
rect 53840 262268 53892 262274
rect 53840 262210 53892 262216
rect 54852 262268 54904 262274
rect 54852 262210 54904 262216
rect 54864 230450 54892 262210
rect 54852 230444 54904 230450
rect 54852 230386 54904 230392
rect 54956 213217 54984 280230
rect 55048 260846 55076 357410
rect 57886 298752 57942 298761
rect 57886 298687 57942 298696
rect 55128 280220 55180 280226
rect 55128 280162 55180 280168
rect 55036 260840 55088 260846
rect 55036 260782 55088 260788
rect 55036 258120 55088 258126
rect 55036 258062 55088 258068
rect 54942 213208 54998 213217
rect 54942 213143 54998 213152
rect 55048 207806 55076 258062
rect 55036 207800 55088 207806
rect 55036 207742 55088 207748
rect 53746 180024 53802 180033
rect 53746 179959 53802 179968
rect 55140 178673 55168 280162
rect 56508 277500 56560 277506
rect 56508 277442 56560 277448
rect 56416 262336 56468 262342
rect 56416 262278 56468 262284
rect 56324 251320 56376 251326
rect 56324 251262 56376 251268
rect 56336 220182 56364 251262
rect 56428 222970 56456 262278
rect 56416 222964 56468 222970
rect 56416 222906 56468 222912
rect 56324 220176 56376 220182
rect 56324 220118 56376 220124
rect 56520 200802 56548 277442
rect 57244 273964 57296 273970
rect 57244 273906 57296 273912
rect 57256 273290 57284 273906
rect 57244 273284 57296 273290
rect 57244 273226 57296 273232
rect 57612 273284 57664 273290
rect 57612 273226 57664 273232
rect 57624 229022 57652 273226
rect 57704 258188 57756 258194
rect 57704 258130 57756 258136
rect 57612 229016 57664 229022
rect 57612 228958 57664 228964
rect 57716 203658 57744 258130
rect 57796 247104 57848 247110
rect 57796 247046 57848 247052
rect 57704 203652 57756 203658
rect 57704 203594 57756 203600
rect 56508 200796 56560 200802
rect 56508 200738 56560 200744
rect 57808 191049 57836 247046
rect 57900 241466 57928 298687
rect 57888 241460 57940 241466
rect 57888 241402 57940 241408
rect 58636 238814 58664 397462
rect 60648 285796 60700 285802
rect 60648 285738 60700 285744
rect 60464 263628 60516 263634
rect 60464 263570 60516 263576
rect 60372 256828 60424 256834
rect 60372 256770 60424 256776
rect 59268 251864 59320 251870
rect 59268 251806 59320 251812
rect 59176 247172 59228 247178
rect 59176 247114 59228 247120
rect 59084 244928 59136 244934
rect 59084 244870 59136 244876
rect 59096 244322 59124 244870
rect 59084 244316 59136 244322
rect 59084 244258 59136 244264
rect 58624 238808 58676 238814
rect 58624 238750 58676 238756
rect 59096 233238 59124 244258
rect 59084 233232 59136 233238
rect 59084 233174 59136 233180
rect 59188 205018 59216 247114
rect 59176 205012 59228 205018
rect 59176 204954 59228 204960
rect 57794 191040 57850 191049
rect 57794 190975 57850 190984
rect 59280 185638 59308 251806
rect 60384 235346 60412 256770
rect 60476 238950 60504 263570
rect 60556 249824 60608 249830
rect 60556 249766 60608 249772
rect 60464 238944 60516 238950
rect 60464 238886 60516 238892
rect 60372 235340 60424 235346
rect 60372 235282 60424 235288
rect 60568 202162 60596 249766
rect 60556 202156 60608 202162
rect 60556 202098 60608 202104
rect 60660 189689 60688 285738
rect 62028 271992 62080 271998
rect 62028 271934 62080 271940
rect 62302 271960 62358 271969
rect 61936 254040 61988 254046
rect 61936 253982 61988 253988
rect 61844 253972 61896 253978
rect 61844 253914 61896 253920
rect 61752 241528 61804 241534
rect 61752 241470 61804 241476
rect 61764 211818 61792 241470
rect 61856 231810 61884 253914
rect 61948 238882 61976 253982
rect 61936 238876 61988 238882
rect 61936 238818 61988 238824
rect 62040 233918 62068 271934
rect 62302 271895 62358 271904
rect 62316 271862 62344 271895
rect 62776 271862 62804 700266
rect 64696 368620 64748 368626
rect 64696 368562 64748 368568
rect 62856 347064 62908 347070
rect 62856 347006 62908 347012
rect 62868 287054 62896 347006
rect 62868 287026 63264 287054
rect 62304 271856 62356 271862
rect 62304 271798 62356 271804
rect 62764 271856 62816 271862
rect 62764 271798 62816 271804
rect 63236 267034 63264 287026
rect 64708 282878 64736 368562
rect 69204 364472 69256 364478
rect 69204 364414 69256 364420
rect 69112 360256 69164 360262
rect 69112 360198 69164 360204
rect 68652 356720 68704 356726
rect 68652 356662 68704 356668
rect 66168 299532 66220 299538
rect 66168 299474 66220 299480
rect 65616 294092 65668 294098
rect 65616 294034 65668 294040
rect 64788 288448 64840 288454
rect 64788 288390 64840 288396
rect 64696 282872 64748 282878
rect 64696 282814 64748 282820
rect 64696 276140 64748 276146
rect 64696 276082 64748 276088
rect 63408 274712 63460 274718
rect 63408 274654 63460 274660
rect 63224 267028 63276 267034
rect 63224 266970 63276 266976
rect 62764 261520 62816 261526
rect 62764 261462 62816 261468
rect 62776 238746 62804 261462
rect 62764 238740 62816 238746
rect 62764 238682 62816 238688
rect 63236 237250 63264 266970
rect 63316 255332 63368 255338
rect 63316 255274 63368 255280
rect 63224 237244 63276 237250
rect 63224 237186 63276 237192
rect 62028 233912 62080 233918
rect 62028 233854 62080 233860
rect 61844 231804 61896 231810
rect 61844 231746 61896 231752
rect 61752 211812 61804 211818
rect 61752 211754 61804 211760
rect 60646 189680 60702 189689
rect 60646 189615 60702 189624
rect 59268 185632 59320 185638
rect 59268 185574 59320 185580
rect 63328 184346 63356 255274
rect 63420 187134 63448 274654
rect 64604 273352 64656 273358
rect 64604 273294 64656 273300
rect 64512 251932 64564 251938
rect 64512 251874 64564 251880
rect 64524 239494 64552 251874
rect 64512 239488 64564 239494
rect 64512 239430 64564 239436
rect 64616 225593 64644 273294
rect 64602 225584 64658 225593
rect 64602 225519 64658 225528
rect 64708 221542 64736 276082
rect 64696 221536 64748 221542
rect 64696 221478 64748 221484
rect 63408 187128 63460 187134
rect 63408 187070 63460 187076
rect 63316 184340 63368 184346
rect 63316 184282 63368 184288
rect 64800 180198 64828 288390
rect 65628 287706 65656 294034
rect 65616 287700 65668 287706
rect 65616 287642 65668 287648
rect 66180 284306 66208 299474
rect 67548 298172 67600 298178
rect 67548 298114 67600 298120
rect 67272 295384 67324 295390
rect 67272 295326 67324 295332
rect 67284 289338 67312 295326
rect 67364 292596 67416 292602
rect 67364 292538 67416 292544
rect 67272 289332 67324 289338
rect 67272 289274 67324 289280
rect 66168 284300 66220 284306
rect 66168 284242 66220 284248
rect 66076 269204 66128 269210
rect 66076 269146 66128 269152
rect 65984 248668 66036 248674
rect 65984 248610 66036 248616
rect 65996 218890 66024 248610
rect 66088 227050 66116 269146
rect 66168 268252 66220 268258
rect 66168 268194 66220 268200
rect 66076 227044 66128 227050
rect 66076 226986 66128 226992
rect 65984 218884 66036 218890
rect 65984 218826 66036 218832
rect 66180 196858 66208 268194
rect 67270 261896 67326 261905
rect 67270 261831 67326 261840
rect 67284 225622 67312 261831
rect 67376 228410 67404 292538
rect 67456 291236 67508 291242
rect 67456 291178 67508 291184
rect 67364 228404 67416 228410
rect 67364 228346 67416 228352
rect 67272 225616 67324 225622
rect 67272 225558 67324 225564
rect 67468 209166 67496 291178
rect 67560 291122 67588 298114
rect 68664 295746 68692 356662
rect 68742 296848 68798 296857
rect 68742 296783 68798 296792
rect 68388 295718 68692 295746
rect 67730 291136 67786 291145
rect 67560 291094 67730 291122
rect 67730 291071 67786 291080
rect 67744 290494 67772 291071
rect 67732 290488 67784 290494
rect 67638 290456 67694 290465
rect 67732 290430 67784 290436
rect 67638 290391 67694 290400
rect 67652 289882 67680 290391
rect 67640 289876 67692 289882
rect 67640 289818 67692 289824
rect 67548 289332 67600 289338
rect 67548 289274 67600 289280
rect 67560 287026 67588 289274
rect 67638 289096 67694 289105
rect 67638 289031 67694 289040
rect 67652 288454 67680 289031
rect 67640 288448 67692 288454
rect 68388 288425 68416 295718
rect 68756 295610 68784 296783
rect 68480 295582 68784 295610
rect 67640 288390 67692 288396
rect 68374 288416 68430 288425
rect 68374 288351 68430 288360
rect 67638 287736 67694 287745
rect 67638 287671 67694 287680
rect 67652 287094 67680 287671
rect 67640 287088 67692 287094
rect 67640 287030 67692 287036
rect 67730 287056 67786 287065
rect 67548 287020 67600 287026
rect 67730 286991 67786 287000
rect 67548 286962 67600 286968
rect 67560 286385 67588 286962
rect 67546 286376 67602 286385
rect 67546 286311 67602 286320
rect 67744 285802 67772 286991
rect 67732 285796 67784 285802
rect 67732 285738 67784 285744
rect 67640 285728 67692 285734
rect 67638 285696 67640 285705
rect 67692 285696 67694 285705
rect 67638 285631 67694 285640
rect 68282 284336 68338 284345
rect 67640 284300 67692 284306
rect 68282 284271 68338 284280
rect 67640 284242 67692 284248
rect 67652 282985 67680 284242
rect 67638 282976 67694 282985
rect 67638 282911 67694 282920
rect 67640 282872 67692 282878
rect 67640 282814 67692 282820
rect 67652 281625 67680 282814
rect 67638 281616 67694 281625
rect 67638 281551 67694 281560
rect 67730 280936 67786 280945
rect 67730 280871 67786 280880
rect 67640 280288 67692 280294
rect 67638 280256 67640 280265
rect 67692 280256 67694 280265
rect 67744 280226 67772 280871
rect 67638 280191 67694 280200
rect 67732 280220 67784 280226
rect 67732 280162 67784 280168
rect 67914 279576 67970 279585
rect 67914 279511 67970 279520
rect 67928 279478 67956 279511
rect 67916 279472 67968 279478
rect 67916 279414 67968 279420
rect 67730 278216 67786 278225
rect 67730 278151 67786 278160
rect 67638 277536 67694 277545
rect 67638 277471 67640 277480
rect 67692 277471 67694 277480
rect 67640 277442 67692 277448
rect 67744 277438 67772 278151
rect 67732 277432 67784 277438
rect 67732 277374 67784 277380
rect 67730 276856 67786 276865
rect 67730 276791 67786 276800
rect 67638 276176 67694 276185
rect 67638 276111 67640 276120
rect 67692 276111 67694 276120
rect 67640 276082 67692 276088
rect 67744 276078 67772 276791
rect 67732 276072 67784 276078
rect 67732 276014 67784 276020
rect 67638 274816 67694 274825
rect 67638 274751 67694 274760
rect 67652 274718 67680 274751
rect 67640 274712 67692 274718
rect 67640 274654 67692 274660
rect 67730 274136 67786 274145
rect 67730 274071 67786 274080
rect 67638 273456 67694 273465
rect 67638 273391 67694 273400
rect 67652 273358 67680 273391
rect 67640 273352 67692 273358
rect 67640 273294 67692 273300
rect 67744 273290 67772 274071
rect 67732 273284 67784 273290
rect 67732 273226 67784 273232
rect 67730 272776 67786 272785
rect 67730 272711 67786 272720
rect 67638 272096 67694 272105
rect 67638 272031 67694 272040
rect 67652 271930 67680 272031
rect 67744 271998 67772 272711
rect 67732 271992 67784 271998
rect 67732 271934 67784 271940
rect 67640 271924 67692 271930
rect 67640 271866 67692 271872
rect 67732 271856 67784 271862
rect 67732 271798 67784 271804
rect 67638 271416 67694 271425
rect 67638 271351 67694 271360
rect 67652 270570 67680 271351
rect 67744 270745 67772 271798
rect 67730 270736 67786 270745
rect 67730 270671 67786 270680
rect 67640 270564 67692 270570
rect 67640 270506 67692 270512
rect 67638 270056 67694 270065
rect 67638 269991 67694 270000
rect 67652 269142 67680 269991
rect 68190 269376 68246 269385
rect 68190 269311 68246 269320
rect 68204 269210 68232 269311
rect 68192 269204 68244 269210
rect 68192 269146 68244 269152
rect 67640 269136 67692 269142
rect 67640 269078 67692 269084
rect 68190 268696 68246 268705
rect 68190 268631 68246 268640
rect 68204 268258 68232 268631
rect 68192 268252 68244 268258
rect 68192 268194 68244 268200
rect 67638 268016 67694 268025
rect 67638 267951 67694 267960
rect 67652 267782 67680 267951
rect 67640 267776 67692 267782
rect 67640 267718 67692 267724
rect 67640 267028 67692 267034
rect 67640 266970 67692 266976
rect 67652 266665 67680 266970
rect 67638 266656 67694 266665
rect 67638 266591 67694 266600
rect 67732 266348 67784 266354
rect 67732 266290 67784 266296
rect 67638 265976 67694 265985
rect 67638 265911 67694 265920
rect 67652 264994 67680 265911
rect 67744 265305 67772 266290
rect 67730 265296 67786 265305
rect 67730 265231 67786 265240
rect 67640 264988 67692 264994
rect 67640 264930 67692 264936
rect 67730 264616 67786 264625
rect 67730 264551 67786 264560
rect 67638 263936 67694 263945
rect 67638 263871 67694 263880
rect 67652 263702 67680 263871
rect 67640 263696 67692 263702
rect 67640 263638 67692 263644
rect 67744 263634 67772 264551
rect 67732 263628 67784 263634
rect 67732 263570 67784 263576
rect 67730 263256 67786 263265
rect 67730 263191 67786 263200
rect 67638 262576 67694 262585
rect 67638 262511 67694 262520
rect 67652 262342 67680 262511
rect 67640 262336 67692 262342
rect 67640 262278 67692 262284
rect 67744 262274 67772 263191
rect 67732 262268 67784 262274
rect 67732 262210 67784 262216
rect 67640 260840 67692 260846
rect 67640 260782 67692 260788
rect 67652 260545 67680 260782
rect 67638 260536 67694 260545
rect 67638 260471 67694 260480
rect 68098 259856 68154 259865
rect 68098 259791 68154 259800
rect 67730 259176 67786 259185
rect 67730 259111 67786 259120
rect 67638 258496 67694 258505
rect 67638 258431 67694 258440
rect 67652 258126 67680 258431
rect 67744 258194 67772 259111
rect 67732 258188 67784 258194
rect 67732 258130 67784 258136
rect 67640 258120 67692 258126
rect 67640 258062 67692 258068
rect 67638 257136 67694 257145
rect 67638 257071 67694 257080
rect 67652 256834 67680 257071
rect 67640 256828 67692 256834
rect 67640 256770 67692 256776
rect 67638 256456 67694 256465
rect 67638 256391 67694 256400
rect 67652 255338 67680 256391
rect 67640 255332 67692 255338
rect 67640 255274 67692 255280
rect 67730 255096 67786 255105
rect 67730 255031 67786 255040
rect 67638 254416 67694 254425
rect 67638 254351 67694 254360
rect 67652 254046 67680 254351
rect 67640 254040 67692 254046
rect 67640 253982 67692 253988
rect 67744 253978 67772 255031
rect 67732 253972 67784 253978
rect 67732 253914 67784 253920
rect 67640 253904 67692 253910
rect 67640 253846 67692 253852
rect 67652 253745 67680 253846
rect 67638 253736 67694 253745
rect 67638 253671 67694 253680
rect 67638 253056 67694 253065
rect 67638 252991 67694 253000
rect 67652 252618 67680 252991
rect 67640 252612 67692 252618
rect 67640 252554 67692 252560
rect 67638 252376 67694 252385
rect 67638 252311 67694 252320
rect 67546 251696 67602 251705
rect 67546 251631 67602 251640
rect 67456 209160 67508 209166
rect 67456 209102 67508 209108
rect 66168 196852 66220 196858
rect 66168 196794 66220 196800
rect 64788 180192 64840 180198
rect 64788 180134 64840 180140
rect 55126 178664 55182 178673
rect 55126 178599 55182 178608
rect 66074 129296 66130 129305
rect 66074 129231 66130 129240
rect 59268 125656 59320 125662
rect 59268 125598 59320 125604
rect 59280 95062 59308 125598
rect 66088 125474 66116 129231
rect 66166 126304 66222 126313
rect 66166 126239 66222 126248
rect 66180 125662 66208 126239
rect 66168 125656 66220 125662
rect 66168 125598 66220 125604
rect 66088 125446 66208 125474
rect 65522 125216 65578 125225
rect 65522 125151 65578 125160
rect 65536 124234 65564 125151
rect 63316 124228 63368 124234
rect 63316 124170 63368 124176
rect 65524 124228 65576 124234
rect 65524 124170 65576 124176
rect 62028 122868 62080 122874
rect 62028 122810 62080 122816
rect 59268 95056 59320 95062
rect 59268 94998 59320 95004
rect 62040 93838 62068 122810
rect 62028 93832 62080 93838
rect 62028 93774 62080 93780
rect 63328 90953 63356 124170
rect 66074 123584 66130 123593
rect 66074 123519 66130 123528
rect 66088 122874 66116 123519
rect 66076 122868 66128 122874
rect 66076 122810 66128 122816
rect 66074 122632 66130 122641
rect 66074 122567 66130 122576
rect 66088 121514 66116 122567
rect 63408 121508 63460 121514
rect 63408 121450 63460 121456
rect 66076 121508 66128 121514
rect 66076 121450 66128 121456
rect 63314 90944 63370 90953
rect 63314 90879 63370 90888
rect 50988 82816 51040 82822
rect 50988 82758 51040 82764
rect 63420 75886 63448 121450
rect 66074 102368 66130 102377
rect 66074 102303 66130 102312
rect 66088 89622 66116 102303
rect 66180 94897 66208 125446
rect 67454 120864 67510 120873
rect 67454 120799 67510 120808
rect 66166 94888 66222 94897
rect 66166 94823 66222 94832
rect 67468 89690 67496 120799
rect 67560 91089 67588 251631
rect 67652 251326 67680 252311
rect 68112 251938 68140 259791
rect 68296 257281 68324 284271
rect 68480 283665 68508 295582
rect 68560 295520 68612 295526
rect 68560 295462 68612 295468
rect 68572 285025 68600 295462
rect 68836 292664 68888 292670
rect 68836 292606 68888 292612
rect 68558 285016 68614 285025
rect 68558 284951 68614 284960
rect 68466 283656 68522 283665
rect 68466 283591 68522 283600
rect 68848 279585 68876 292606
rect 68834 279576 68890 279585
rect 68834 279511 68890 279520
rect 68926 275496 68982 275505
rect 68926 275431 68982 275440
rect 68374 261216 68430 261225
rect 68374 261151 68430 261160
rect 68282 257272 68338 257281
rect 68282 257207 68338 257216
rect 68100 251932 68152 251938
rect 68100 251874 68152 251880
rect 68388 251870 68416 261151
rect 68834 255776 68890 255785
rect 68834 255711 68890 255720
rect 68376 251864 68428 251870
rect 68376 251806 68428 251812
rect 67640 251320 67692 251326
rect 67640 251262 67692 251268
rect 68742 251016 68798 251025
rect 68742 250951 68798 250960
rect 67638 250336 67694 250345
rect 67638 250271 67694 250280
rect 67652 249830 67680 250271
rect 67640 249824 67692 249830
rect 67640 249766 67692 249772
rect 67822 248976 67878 248985
rect 67822 248911 67878 248920
rect 67836 248674 67864 248911
rect 67824 248668 67876 248674
rect 67824 248610 67876 248616
rect 67730 248296 67786 248305
rect 67730 248231 67786 248240
rect 67638 247616 67694 247625
rect 67638 247551 67694 247560
rect 67652 247178 67680 247551
rect 67640 247172 67692 247178
rect 67640 247114 67692 247120
rect 67744 247110 67772 248231
rect 67732 247104 67784 247110
rect 67732 247046 67784 247052
rect 68650 246256 68706 246265
rect 68650 246191 68706 246200
rect 67638 245576 67694 245585
rect 67638 245511 67694 245520
rect 67652 244322 67680 245511
rect 67640 244316 67692 244322
rect 67640 244258 67692 244264
rect 67730 242176 67786 242185
rect 67730 242111 67786 242120
rect 67744 241534 67772 242111
rect 67732 241528 67784 241534
rect 67638 241496 67694 241505
rect 67732 241470 67784 241476
rect 67638 241431 67640 241440
rect 67692 241431 67694 241440
rect 67640 241402 67692 241408
rect 68664 232558 68692 246191
rect 68756 233889 68784 250951
rect 68742 233880 68798 233889
rect 68742 233815 68798 233824
rect 68652 232552 68704 232558
rect 68652 232494 68704 232500
rect 68848 214577 68876 255711
rect 68940 249762 68968 275431
rect 69124 258074 69152 360198
rect 69032 258046 69152 258074
rect 69032 257825 69060 258046
rect 69018 257816 69074 257825
rect 69018 257751 69074 257760
rect 69032 256766 69060 257751
rect 69020 256760 69072 256766
rect 69020 256702 69072 256708
rect 68928 249756 68980 249762
rect 68928 249698 68980 249704
rect 69110 244896 69166 244905
rect 69110 244831 69166 244840
rect 68926 244216 68982 244225
rect 68926 244151 68982 244160
rect 68834 214568 68890 214577
rect 68834 214503 68890 214512
rect 68940 185774 68968 244151
rect 69020 233980 69072 233986
rect 69020 233922 69072 233928
rect 68928 185768 68980 185774
rect 68928 185710 68980 185716
rect 69032 185706 69060 233922
rect 69124 223038 69152 244831
rect 69216 244254 69244 364414
rect 79324 361616 79376 361622
rect 79324 361558 79376 361564
rect 75920 354816 75972 354822
rect 75920 354758 75972 354764
rect 72424 344344 72476 344350
rect 72424 344286 72476 344292
rect 72436 306374 72464 344286
rect 72252 306346 72464 306374
rect 72252 304978 72280 306346
rect 75368 305108 75420 305114
rect 75368 305050 75420 305056
rect 72240 304972 72292 304978
rect 72240 304914 72292 304920
rect 70952 300144 71004 300150
rect 70952 300086 71004 300092
rect 70676 292596 70728 292602
rect 70676 292538 70728 292544
rect 70688 291924 70716 292538
rect 70964 291938 70992 300086
rect 71964 294636 72016 294642
rect 71964 294578 72016 294584
rect 71688 292528 71740 292534
rect 71688 292470 71740 292476
rect 71700 292369 71728 292470
rect 71686 292360 71742 292369
rect 71686 292295 71742 292304
rect 70964 291910 71346 291938
rect 71976 291924 72004 294578
rect 72252 291938 72280 304914
rect 74540 302252 74592 302258
rect 74540 302194 74592 302200
rect 73252 294772 73304 294778
rect 73252 294714 73304 294720
rect 72252 291910 72634 291938
rect 73264 291924 73292 294714
rect 73894 292904 73950 292913
rect 73894 292839 73950 292848
rect 73908 291924 73936 292839
rect 74552 291924 74580 302194
rect 75184 296880 75236 296886
rect 75184 296822 75236 296828
rect 75196 291924 75224 296822
rect 75380 291938 75408 305050
rect 75932 294030 75960 354758
rect 76102 300928 76158 300937
rect 76102 300863 76158 300872
rect 75920 294024 75972 294030
rect 75920 293966 75972 293972
rect 76116 291938 76144 300863
rect 78588 294160 78640 294166
rect 78588 294102 78640 294108
rect 76748 294024 76800 294030
rect 76748 293966 76800 293972
rect 76760 291938 76788 293966
rect 78600 293282 78628 294102
rect 79336 294098 79364 361558
rect 80060 356108 80112 356114
rect 80060 356050 80112 356056
rect 79692 294704 79744 294710
rect 79692 294646 79744 294652
rect 79324 294092 79376 294098
rect 79324 294034 79376 294040
rect 78588 293276 78640 293282
rect 78588 293218 78640 293224
rect 77758 292768 77814 292777
rect 77758 292703 77814 292712
rect 75380 291910 75854 291938
rect 76116 291910 76498 291938
rect 76760 291910 77142 291938
rect 77772 291924 77800 292703
rect 78402 292632 78458 292641
rect 78402 292567 78458 292576
rect 78416 291924 78444 292567
rect 79336 291938 79364 294034
rect 79074 291910 79364 291938
rect 79704 291924 79732 294646
rect 80072 291938 80100 356050
rect 82096 304298 82124 700334
rect 84292 354068 84344 354074
rect 84292 354010 84344 354016
rect 82176 307828 82228 307834
rect 82176 307770 82228 307776
rect 82084 304292 82136 304298
rect 82084 304234 82136 304240
rect 81440 299600 81492 299606
rect 81440 299542 81492 299548
rect 80980 294228 81032 294234
rect 80980 294170 81032 294176
rect 80072 291910 80362 291938
rect 80992 291924 81020 294170
rect 81452 291938 81480 299542
rect 82188 294778 82216 307770
rect 84200 297084 84252 297090
rect 84200 297026 84252 297032
rect 83556 295656 83608 295662
rect 83556 295598 83608 295604
rect 82268 295588 82320 295594
rect 82268 295530 82320 295536
rect 82176 294772 82228 294778
rect 82176 294714 82228 294720
rect 81452 291910 81650 291938
rect 82280 291924 82308 295530
rect 82912 294024 82964 294030
rect 82912 293966 82964 293972
rect 82924 291924 82952 293966
rect 83568 291924 83596 295598
rect 84212 291924 84240 297026
rect 84304 293962 84332 354010
rect 85580 306400 85632 306406
rect 85580 306342 85632 306348
rect 84384 302932 84436 302938
rect 84384 302874 84436 302880
rect 84396 299577 84424 302874
rect 84382 299568 84438 299577
rect 84382 299503 84438 299512
rect 84292 293956 84344 293962
rect 84292 293898 84344 293904
rect 84396 291938 84424 299503
rect 85592 293962 85620 306342
rect 88352 303618 88380 702406
rect 105464 700398 105492 703520
rect 105452 700392 105504 700398
rect 105452 700334 105504 700340
rect 137848 699802 137876 703520
rect 154132 702434 154160 703520
rect 153212 702406 154160 702434
rect 137848 699774 138060 699802
rect 116584 579692 116636 579698
rect 116584 579634 116636 579640
rect 111064 462392 111116 462398
rect 111064 462334 111116 462340
rect 109040 367124 109092 367130
rect 109040 367066 109092 367072
rect 101404 358828 101456 358834
rect 101404 358770 101456 358776
rect 90364 357536 90416 357542
rect 90364 357478 90416 357484
rect 90376 336054 90404 357478
rect 97264 354884 97316 354890
rect 97264 354826 97316 354832
rect 90364 336048 90416 336054
rect 90364 335990 90416 335996
rect 94504 312588 94556 312594
rect 94504 312530 94556 312536
rect 91100 307080 91152 307086
rect 91100 307022 91152 307028
rect 88340 303612 88392 303618
rect 88340 303554 88392 303560
rect 89720 302320 89772 302326
rect 89720 302262 89772 302268
rect 85672 299668 85724 299674
rect 85672 299610 85724 299616
rect 85212 293956 85264 293962
rect 85212 293898 85264 293904
rect 85580 293956 85632 293962
rect 85580 293898 85632 293904
rect 85224 291938 85252 293898
rect 85684 291938 85712 299610
rect 88064 298308 88116 298314
rect 88064 298250 88116 298256
rect 86500 293956 86552 293962
rect 86500 293898 86552 293904
rect 86512 291938 86540 293898
rect 87420 293276 87472 293282
rect 87420 293218 87472 293224
rect 84396 291910 84870 291938
rect 85224 291910 85514 291938
rect 85684 291910 86158 291938
rect 86512 291910 86802 291938
rect 87432 291924 87460 293218
rect 88076 291924 88104 298250
rect 88708 298240 88760 298246
rect 88708 298182 88760 298188
rect 89350 298208 89406 298217
rect 88720 291924 88748 298182
rect 89350 298143 89406 298152
rect 89364 291924 89392 298143
rect 89732 291938 89760 302262
rect 90272 300960 90324 300966
rect 90272 300902 90324 300908
rect 90284 291938 90312 300902
rect 91112 291938 91140 307022
rect 92848 299804 92900 299810
rect 92848 299746 92900 299752
rect 92572 295452 92624 295458
rect 92572 295394 92624 295400
rect 91928 294296 91980 294302
rect 91928 294238 91980 294244
rect 89732 291910 90022 291938
rect 90284 291910 90666 291938
rect 91112 291910 91310 291938
rect 91940 291924 91968 294238
rect 92584 291924 92612 295394
rect 92860 291938 92888 299746
rect 94516 296954 94544 312530
rect 94596 303680 94648 303686
rect 94596 303622 94648 303628
rect 94504 296948 94556 296954
rect 94504 296890 94556 296896
rect 93860 294092 93912 294098
rect 93860 294034 93912 294040
rect 92860 291910 93242 291938
rect 93872 291924 93900 294034
rect 94516 291924 94544 296890
rect 94608 294710 94636 303622
rect 97080 296812 97132 296818
rect 97080 296754 97132 296760
rect 97092 296714 97120 296754
rect 97276 296714 97304 354826
rect 98644 336048 98696 336054
rect 98644 335990 98696 335996
rect 97092 296686 97304 296714
rect 95146 296032 95202 296041
rect 95146 295967 95202 295976
rect 94596 294704 94648 294710
rect 94596 294646 94648 294652
rect 95160 291924 95188 295967
rect 96434 294128 96490 294137
rect 96434 294063 96490 294072
rect 95790 293992 95846 294001
rect 95790 293927 95846 293936
rect 95804 291924 95832 293927
rect 96448 291924 96476 294063
rect 97092 291924 97120 296686
rect 97724 295724 97776 295730
rect 97724 295666 97776 295672
rect 97736 291924 97764 295666
rect 98656 292602 98684 335990
rect 100024 318844 100076 318850
rect 100024 318786 100076 318792
rect 98736 303748 98788 303754
rect 98736 303690 98788 303696
rect 98748 293282 98776 303690
rect 100036 301510 100064 318786
rect 100024 301504 100076 301510
rect 100024 301446 100076 301452
rect 99380 299872 99432 299878
rect 99380 299814 99432 299820
rect 99012 297016 99064 297022
rect 99012 296958 99064 296964
rect 98736 293276 98788 293282
rect 98736 293218 98788 293224
rect 98644 292596 98696 292602
rect 98644 292538 98696 292544
rect 98656 291938 98684 292538
rect 98394 291910 98684 291938
rect 99024 291924 99052 296958
rect 99392 291938 99420 299814
rect 101416 294166 101444 358770
rect 107660 357536 107712 357542
rect 107660 357478 107712 357484
rect 104164 332648 104216 332654
rect 104164 332590 104216 332596
rect 104176 303618 104204 332590
rect 106280 330540 106332 330546
rect 106280 330482 106332 330488
rect 106292 306374 106320 330482
rect 107672 306374 107700 357478
rect 106292 306346 106872 306374
rect 107672 306346 108344 306374
rect 104164 303612 104216 303618
rect 104164 303554 104216 303560
rect 104440 303612 104492 303618
rect 104440 303554 104492 303560
rect 103704 301028 103756 301034
rect 103704 300970 103756 300976
rect 102232 298444 102284 298450
rect 102232 298386 102284 298392
rect 101404 294160 101456 294166
rect 101404 294102 101456 294108
rect 101416 291938 101444 294102
rect 99392 291910 99682 291938
rect 100970 291922 101352 291938
rect 100970 291916 101364 291922
rect 100970 291910 101312 291916
rect 101416 291910 101614 291938
rect 102244 291924 102272 298386
rect 102876 292800 102928 292806
rect 102876 292742 102928 292748
rect 102888 291924 102916 292742
rect 103716 291938 103744 300970
rect 104452 291938 104480 303554
rect 106740 298376 106792 298382
rect 106740 298318 106792 298324
rect 104898 297392 104954 297401
rect 104898 297327 104954 297336
rect 104912 296041 104940 297327
rect 104898 296032 104954 296041
rect 104898 295967 104954 295976
rect 106094 295352 106150 295361
rect 106094 295287 106150 295296
rect 105452 294160 105504 294166
rect 105452 294102 105504 294108
rect 103546 291922 103652 291938
rect 103546 291916 103664 291922
rect 103546 291910 103612 291916
rect 101312 291858 101364 291864
rect 103716 291910 104190 291938
rect 104452 291910 104834 291938
rect 105464 291924 105492 294102
rect 106108 291924 106136 295287
rect 106752 291924 106780 298318
rect 106844 292074 106872 306346
rect 106924 301096 106976 301102
rect 106924 301038 106976 301044
rect 106936 294642 106964 301038
rect 106924 294636 106976 294642
rect 106924 294578 106976 294584
rect 108026 294264 108082 294273
rect 108026 294199 108082 294208
rect 106844 292046 107056 292074
rect 107028 291938 107056 292046
rect 107028 291910 107410 291938
rect 108040 291924 108068 294199
rect 108316 291938 108344 306346
rect 109052 293962 109080 367066
rect 111076 355366 111104 462334
rect 114558 358864 114614 358873
rect 114558 358799 114614 358808
rect 111156 356176 111208 356182
rect 111156 356118 111208 356124
rect 111064 355360 111116 355366
rect 111064 355302 111116 355308
rect 109132 299736 109184 299742
rect 109132 299678 109184 299684
rect 109040 293956 109092 293962
rect 109040 293898 109092 293904
rect 109144 291938 109172 299678
rect 109684 293956 109736 293962
rect 109684 293898 109736 293904
rect 109696 291938 109724 293898
rect 111168 292534 111196 356118
rect 113180 352572 113232 352578
rect 113180 352514 113232 352520
rect 111248 296812 111300 296818
rect 111248 296754 111300 296760
rect 111156 292528 111208 292534
rect 111156 292470 111208 292476
rect 108316 291910 108698 291938
rect 109144 291910 109342 291938
rect 109696 291910 109986 291938
rect 110630 291922 110920 291938
rect 111260 291924 111288 296754
rect 111892 294364 111944 294370
rect 111892 294306 111944 294312
rect 111904 291924 111932 294306
rect 112536 292868 112588 292874
rect 112536 292810 112588 292816
rect 112548 291924 112576 292810
rect 113192 291924 113220 352514
rect 113824 296744 113876 296750
rect 113824 296686 113876 296692
rect 113836 291924 113864 296686
rect 114466 294128 114522 294137
rect 114466 294063 114522 294072
rect 114480 291924 114508 294063
rect 114572 293962 114600 358799
rect 116596 312798 116624 579634
rect 122748 373312 122800 373318
rect 122748 373254 122800 373260
rect 117964 363112 118016 363118
rect 117964 363054 118016 363060
rect 116584 312792 116636 312798
rect 116584 312734 116636 312740
rect 115848 304292 115900 304298
rect 115848 304234 115900 304240
rect 115860 302190 115888 304234
rect 114744 302184 114796 302190
rect 114744 302126 114796 302132
rect 115848 302184 115900 302190
rect 115848 302126 115900 302132
rect 114560 293956 114612 293962
rect 114560 293898 114612 293904
rect 114756 291938 114784 302126
rect 116584 301504 116636 301510
rect 116584 301446 116636 301452
rect 116596 294098 116624 301446
rect 117976 300898 118004 363054
rect 120080 320884 120132 320890
rect 120080 320826 120132 320832
rect 119620 313948 119672 313954
rect 119620 313890 119672 313896
rect 117964 300892 118016 300898
rect 117964 300834 118016 300840
rect 117976 296714 118004 300834
rect 117884 296686 118004 296714
rect 115848 294092 115900 294098
rect 115848 294034 115900 294040
rect 116584 294092 116636 294098
rect 116584 294034 116636 294040
rect 115388 293956 115440 293962
rect 115388 293898 115440 293904
rect 115400 291938 115428 293898
rect 115860 293282 115888 294034
rect 115848 293276 115900 293282
rect 115848 293218 115900 293224
rect 116596 291938 116624 294034
rect 117044 292732 117096 292738
rect 117044 292674 117096 292680
rect 110630 291916 110932 291922
rect 110630 291910 110880 291916
rect 103612 291858 103664 291864
rect 114756 291910 115138 291938
rect 115400 291910 115782 291938
rect 116426 291910 116624 291938
rect 117056 291924 117084 292674
rect 117778 291952 117834 291961
rect 117714 291910 117778 291938
rect 117884 291938 117912 296686
rect 119632 292210 119660 313890
rect 119632 292182 119844 292210
rect 117884 291910 118358 291938
rect 119002 291922 119384 291938
rect 119632 291924 119660 292182
rect 119002 291916 119396 291922
rect 119002 291910 119344 291916
rect 117778 291887 117834 291896
rect 110880 291858 110932 291864
rect 119344 291858 119396 291864
rect 119712 291916 119764 291922
rect 119712 291858 119764 291864
rect 69768 291242 70058 291258
rect 69756 291236 70058 291242
rect 69808 291230 70058 291236
rect 69756 291178 69808 291184
rect 119724 267734 119752 291858
rect 119816 291310 119844 292182
rect 119804 291304 119856 291310
rect 119804 291246 119856 291252
rect 120092 268705 120120 320826
rect 121460 312792 121512 312798
rect 121460 312734 121512 312740
rect 120172 305040 120224 305046
rect 120172 304982 120224 304988
rect 120184 286385 120212 304982
rect 120724 296744 120776 296750
rect 120724 296686 120776 296692
rect 120170 286376 120226 286385
rect 120170 286311 120226 286320
rect 120078 268696 120134 268705
rect 120078 268631 120134 268640
rect 120092 267782 120120 268631
rect 120080 267776 120132 267782
rect 119724 267706 119844 267734
rect 120080 267718 120132 267724
rect 69664 249756 69716 249762
rect 69664 249698 69716 249704
rect 69204 244248 69256 244254
rect 69204 244190 69256 244196
rect 69216 243545 69244 244190
rect 69202 243536 69258 243545
rect 69202 243471 69258 243480
rect 69112 223032 69164 223038
rect 69112 222974 69164 222980
rect 69676 196722 69704 249698
rect 119816 244934 119844 267706
rect 120632 251184 120684 251190
rect 120632 251126 120684 251132
rect 120644 251025 120672 251126
rect 120170 251016 120226 251025
rect 120170 250951 120226 250960
rect 120630 251016 120686 251025
rect 120630 250951 120686 250960
rect 119804 244928 119856 244934
rect 119804 244870 119856 244876
rect 119802 242584 119858 242593
rect 119802 242519 119858 242528
rect 69846 240816 69902 240825
rect 69846 240751 69902 240760
rect 69860 240242 69888 240751
rect 69848 240236 69900 240242
rect 69848 240178 69900 240184
rect 69768 240094 70058 240122
rect 69768 233986 69796 240094
rect 70308 239420 70360 239426
rect 70308 239362 70360 239368
rect 70320 238678 70348 239362
rect 70308 238672 70360 238678
rect 70308 238614 70360 238620
rect 70688 238134 70716 240108
rect 70676 238128 70728 238134
rect 70676 238070 70728 238076
rect 69756 233980 69808 233986
rect 69756 233922 69808 233928
rect 71332 219434 71360 240108
rect 71976 219434 72004 240108
rect 72620 235890 72648 240108
rect 72608 235884 72660 235890
rect 72608 235826 72660 235832
rect 73160 229356 73212 229362
rect 73160 229298 73212 229304
rect 70412 219406 71360 219434
rect 71792 219406 72004 219434
rect 70412 205086 70440 219406
rect 70400 205080 70452 205086
rect 70400 205022 70452 205028
rect 71792 203590 71820 219406
rect 71780 203584 71832 203590
rect 71780 203526 71832 203532
rect 69664 196716 69716 196722
rect 69664 196658 69716 196664
rect 69020 185700 69072 185706
rect 69020 185642 69072 185648
rect 73172 184249 73200 229298
rect 73264 186998 73292 240108
rect 73908 229362 73936 240108
rect 73896 229356 73948 229362
rect 73896 229298 73948 229304
rect 74552 197985 74580 240108
rect 75196 238754 75224 240108
rect 75276 239964 75328 239970
rect 75276 239906 75328 239912
rect 74644 238726 75224 238754
rect 74644 210458 74672 238726
rect 75288 219434 75316 239906
rect 75840 238202 75868 240108
rect 75828 238196 75880 238202
rect 75828 238138 75880 238144
rect 75920 233980 75972 233986
rect 75920 233922 75972 233928
rect 75196 219406 75316 219434
rect 74632 210452 74684 210458
rect 74632 210394 74684 210400
rect 74538 197976 74594 197985
rect 74538 197911 74594 197920
rect 73252 186992 73304 186998
rect 73252 186934 73304 186940
rect 73158 184240 73214 184249
rect 73158 184175 73214 184184
rect 75196 181393 75224 219406
rect 75932 206310 75960 233922
rect 76484 219434 76512 240108
rect 77128 233986 77156 240108
rect 77116 233980 77168 233986
rect 77116 233922 77168 233928
rect 77300 233980 77352 233986
rect 77300 233922 77352 233928
rect 76012 219428 76512 219434
rect 76064 219406 76512 219428
rect 76012 219370 76064 219376
rect 77312 215937 77340 233922
rect 77772 221474 77800 240108
rect 78416 233986 78444 240108
rect 78404 233980 78456 233986
rect 78404 233922 78456 233928
rect 78680 233980 78732 233986
rect 78680 233922 78732 233928
rect 77760 221468 77812 221474
rect 77760 221410 77812 221416
rect 77298 215928 77354 215937
rect 77298 215863 77354 215872
rect 75920 206304 75972 206310
rect 75920 206246 75972 206252
rect 75182 181384 75238 181393
rect 75182 181319 75238 181328
rect 78692 178702 78720 233922
rect 79060 220318 79088 240108
rect 79704 233986 79732 240108
rect 80348 238754 80376 240108
rect 80072 238726 80376 238754
rect 79692 233980 79744 233986
rect 79692 233922 79744 233928
rect 79048 220312 79100 220318
rect 79048 220254 79100 220260
rect 80072 186969 80100 238726
rect 80992 219434 81020 240108
rect 81636 239306 81664 240108
rect 81452 239278 81664 239306
rect 81452 224942 81480 239278
rect 82280 238814 82308 240108
rect 81532 238808 81584 238814
rect 81532 238750 81584 238756
rect 82268 238808 82320 238814
rect 82924 238785 82952 240108
rect 82268 238750 82320 238756
rect 82910 238776 82966 238785
rect 81544 229090 81572 238750
rect 82910 238711 82966 238720
rect 83568 231742 83596 240108
rect 84212 238754 84240 240108
rect 84212 238726 84424 238754
rect 84292 233980 84344 233986
rect 84292 233922 84344 233928
rect 84108 231872 84160 231878
rect 84160 231826 84240 231854
rect 84108 231814 84160 231820
rect 83556 231736 83608 231742
rect 83556 231678 83608 231684
rect 81532 229084 81584 229090
rect 81532 229026 81584 229032
rect 81440 224936 81492 224942
rect 81440 224878 81492 224884
rect 83568 219434 83596 231678
rect 80164 219406 81020 219434
rect 83476 219406 83596 219434
rect 80164 188358 80192 219406
rect 83476 210526 83504 219406
rect 83464 210520 83516 210526
rect 83464 210462 83516 210468
rect 80152 188352 80204 188358
rect 80152 188294 80204 188300
rect 80058 186960 80114 186969
rect 80058 186895 80114 186904
rect 84212 184278 84240 231826
rect 84304 189786 84332 233922
rect 84396 210361 84424 238726
rect 84856 231878 84884 240108
rect 85500 233986 85528 240108
rect 86144 238270 86172 240108
rect 86788 238746 86816 240108
rect 87432 238754 87460 240108
rect 86776 238740 86828 238746
rect 86776 238682 86828 238688
rect 86972 238726 87460 238754
rect 86132 238264 86184 238270
rect 86132 238206 86184 238212
rect 86224 238196 86276 238202
rect 86224 238138 86276 238144
rect 85488 233980 85540 233986
rect 85488 233922 85540 233928
rect 84844 231872 84896 231878
rect 84844 231814 84896 231820
rect 86236 227730 86264 238138
rect 86788 233170 86816 238682
rect 86776 233164 86828 233170
rect 86776 233106 86828 233112
rect 86224 227724 86276 227730
rect 86224 227666 86276 227672
rect 86972 213246 87000 238726
rect 88076 221610 88104 240108
rect 88064 221604 88116 221610
rect 88064 221546 88116 221552
rect 88720 219434 88748 240108
rect 89364 238406 89392 240108
rect 90008 238754 90036 240108
rect 89732 238726 90036 238754
rect 89352 238400 89404 238406
rect 89352 238342 89404 238348
rect 88352 219406 88748 219434
rect 86960 213240 87012 213246
rect 86960 213182 87012 213188
rect 84382 210352 84438 210361
rect 84382 210287 84438 210296
rect 84292 189780 84344 189786
rect 84292 189722 84344 189728
rect 84200 184272 84252 184278
rect 84200 184214 84252 184220
rect 88352 184210 88380 219406
rect 89732 195498 89760 238726
rect 90652 219434 90680 240108
rect 91296 234530 91324 240108
rect 91940 237386 91968 240108
rect 91928 237380 91980 237386
rect 91928 237322 91980 237328
rect 91284 234524 91336 234530
rect 91284 234466 91336 234472
rect 92480 233436 92532 233442
rect 92480 233378 92532 233384
rect 89824 219406 90680 219434
rect 89824 211886 89852 219406
rect 89812 211880 89864 211886
rect 89812 211822 89864 211828
rect 89720 195492 89772 195498
rect 89720 195434 89772 195440
rect 92492 195294 92520 233378
rect 92584 227186 92612 240108
rect 93228 233442 93256 240108
rect 93872 238754 93900 240108
rect 93872 238726 93992 238754
rect 93860 233980 93912 233986
rect 93860 233922 93912 233928
rect 93216 233436 93268 233442
rect 93216 233378 93268 233384
rect 92572 227180 92624 227186
rect 92572 227122 92624 227128
rect 92480 195288 92532 195294
rect 92480 195230 92532 195236
rect 88340 184204 88392 184210
rect 88340 184146 88392 184152
rect 93872 182850 93900 233922
rect 93964 192574 93992 238726
rect 94516 233986 94544 240108
rect 95056 236700 95108 236706
rect 95056 236642 95108 236648
rect 95068 235822 95096 236642
rect 95056 235816 95108 235822
rect 95056 235758 95108 235764
rect 94504 233980 94556 233986
rect 94504 233922 94556 233928
rect 95160 219434 95188 240108
rect 95700 238264 95752 238270
rect 95700 238206 95752 238212
rect 95712 237289 95740 238206
rect 95698 237280 95754 237289
rect 95698 237215 95754 237224
rect 95804 236706 95832 240108
rect 95792 236700 95844 236706
rect 95792 236642 95844 236648
rect 96448 219434 96476 240108
rect 96526 237280 96582 237289
rect 96526 237215 96582 237224
rect 94056 219406 95188 219434
rect 95344 219406 96476 219434
rect 94056 205222 94084 219406
rect 94044 205216 94096 205222
rect 94044 205158 94096 205164
rect 93952 192568 94004 192574
rect 93952 192510 94004 192516
rect 95344 187066 95372 219406
rect 96540 199442 96568 237215
rect 96620 233980 96672 233986
rect 96620 233922 96672 233928
rect 96528 199436 96580 199442
rect 96528 199378 96580 199384
rect 96632 193866 96660 233922
rect 97092 224330 97120 240108
rect 97736 233986 97764 240108
rect 97724 233980 97776 233986
rect 97724 233922 97776 233928
rect 98380 230314 98408 240108
rect 99024 238542 99052 240108
rect 99668 238754 99696 240108
rect 99392 238726 99696 238754
rect 99012 238536 99064 238542
rect 99012 238478 99064 238484
rect 98368 230308 98420 230314
rect 98368 230250 98420 230256
rect 98644 228404 98696 228410
rect 98644 228346 98696 228352
rect 97080 224324 97132 224330
rect 97080 224266 97132 224272
rect 96620 193860 96672 193866
rect 96620 193802 96672 193808
rect 95332 187060 95384 187066
rect 95332 187002 95384 187008
rect 98656 182889 98684 228346
rect 99392 213314 99420 238726
rect 100312 228546 100340 240108
rect 100760 233980 100812 233986
rect 100760 233922 100812 233928
rect 100300 228540 100352 228546
rect 100300 228482 100352 228488
rect 99380 213308 99432 213314
rect 99380 213250 99432 213256
rect 100772 188329 100800 233922
rect 100956 219434 100984 240108
rect 101600 233986 101628 240108
rect 101588 233980 101640 233986
rect 101588 233922 101640 233928
rect 102140 233980 102192 233986
rect 102140 233922 102192 233928
rect 100864 219406 100984 219434
rect 100864 216170 100892 219406
rect 100852 216164 100904 216170
rect 100852 216106 100904 216112
rect 102152 202366 102180 233922
rect 102244 217326 102272 240108
rect 102888 233986 102916 240108
rect 103532 238678 103560 240108
rect 103520 238672 103572 238678
rect 103520 238614 103572 238620
rect 104176 237454 104204 240108
rect 104716 238672 104768 238678
rect 104716 238614 104768 238620
rect 104164 237448 104216 237454
rect 104164 237390 104216 237396
rect 102876 233980 102928 233986
rect 102876 233922 102928 233928
rect 104728 230382 104756 238614
rect 104716 230376 104768 230382
rect 104716 230318 104768 230324
rect 104820 219434 104848 240108
rect 105464 238105 105492 240108
rect 105450 238096 105506 238105
rect 105450 238031 105506 238040
rect 106108 233986 106136 240108
rect 106752 237153 106780 240108
rect 107396 238678 107424 240108
rect 108040 238754 108068 240108
rect 107672 238726 108068 238754
rect 107384 238672 107436 238678
rect 107384 238614 107436 238620
rect 106924 237448 106976 237454
rect 106924 237390 106976 237396
rect 106738 237144 106794 237153
rect 106738 237079 106794 237088
rect 104900 233980 104952 233986
rect 104900 233922 104952 233928
rect 106096 233980 106148 233986
rect 106096 233922 106148 233928
rect 103716 219406 104848 219434
rect 102232 217320 102284 217326
rect 102232 217262 102284 217268
rect 103716 209098 103744 219406
rect 103704 209092 103756 209098
rect 103704 209034 103756 209040
rect 102140 202360 102192 202366
rect 102140 202302 102192 202308
rect 104912 195362 104940 233922
rect 106936 217394 106964 237390
rect 106924 217388 106976 217394
rect 106924 217330 106976 217336
rect 104900 195356 104952 195362
rect 104900 195298 104952 195304
rect 102048 190528 102100 190534
rect 102048 190470 102100 190476
rect 100758 188320 100814 188329
rect 100758 188255 100814 188264
rect 100668 187740 100720 187746
rect 100668 187682 100720 187688
rect 98642 182880 98698 182889
rect 93860 182844 93912 182850
rect 98642 182815 98698 182824
rect 93860 182786 93912 182792
rect 97816 179444 97868 179450
rect 97816 179386 97868 179392
rect 78680 178696 78732 178702
rect 78680 178638 78732 178644
rect 97828 176905 97856 179386
rect 100680 177585 100708 187682
rect 102060 177585 102088 190470
rect 107568 189236 107620 189242
rect 107568 189178 107620 189184
rect 106188 187808 106240 187814
rect 106188 187750 106240 187756
rect 106200 177585 106228 187750
rect 107580 177585 107608 189178
rect 107672 185842 107700 238726
rect 108684 228478 108712 240108
rect 109972 238814 110000 240108
rect 109040 238808 109092 238814
rect 109040 238750 109092 238756
rect 109960 238808 110012 238814
rect 109960 238750 110012 238756
rect 108672 228472 108724 228478
rect 108672 228414 108724 228420
rect 109052 188426 109080 238750
rect 110616 238474 110644 240108
rect 111260 238754 111288 240108
rect 110984 238726 111288 238754
rect 110604 238468 110656 238474
rect 110604 238410 110656 238416
rect 110616 237862 110644 238410
rect 110604 237856 110656 237862
rect 110604 237798 110656 237804
rect 110984 219434 111012 238726
rect 111064 237856 111116 237862
rect 111064 237798 111116 237804
rect 110432 219406 111012 219434
rect 110432 206281 110460 219406
rect 110418 206272 110474 206281
rect 110418 206207 110474 206216
rect 111076 189854 111104 237798
rect 111904 220386 111932 240108
rect 112548 238066 112576 240108
rect 112536 238060 112588 238066
rect 112536 238002 112588 238008
rect 112548 237318 112576 238002
rect 112536 237312 112588 237318
rect 112536 237254 112588 237260
rect 113192 227118 113220 240108
rect 113836 235958 113864 240108
rect 114480 238746 114508 240108
rect 114468 238740 114520 238746
rect 114468 238682 114520 238688
rect 113824 235952 113876 235958
rect 113824 235894 113876 235900
rect 114560 233980 114612 233986
rect 114560 233922 114612 233928
rect 113180 227112 113232 227118
rect 113180 227054 113232 227060
rect 111892 220380 111944 220386
rect 111892 220322 111944 220328
rect 114572 214674 114600 233922
rect 115124 233102 115152 240108
rect 115768 233986 115796 240108
rect 115756 233980 115808 233986
rect 115756 233922 115808 233928
rect 115112 233096 115164 233102
rect 115112 233038 115164 233044
rect 116412 219434 116440 240108
rect 117056 239873 117084 240108
rect 117042 239864 117098 239873
rect 117042 239799 117098 239808
rect 116584 239488 116636 239494
rect 116584 239430 116636 239436
rect 115952 219406 116440 219434
rect 114560 214668 114612 214674
rect 114560 214610 114612 214616
rect 115952 198082 115980 219406
rect 116596 216034 116624 239430
rect 117700 238610 117728 240108
rect 117688 238604 117740 238610
rect 117688 238546 117740 238552
rect 117962 236600 118018 236609
rect 117962 236535 118018 236544
rect 116584 216028 116636 216034
rect 116584 215970 116636 215976
rect 117976 200705 118004 236535
rect 118344 231674 118372 240108
rect 118988 239970 119016 240108
rect 118976 239964 119028 239970
rect 118976 239906 119028 239912
rect 118608 239420 118660 239426
rect 118608 239362 118660 239368
rect 118620 238746 118648 239362
rect 118608 238740 118660 238746
rect 118608 238682 118660 238688
rect 118332 231668 118384 231674
rect 118332 231610 118384 231616
rect 119632 219434 119660 240108
rect 119816 239970 119844 242519
rect 120078 241496 120134 241505
rect 120078 241431 120134 241440
rect 119804 239964 119856 239970
rect 119804 239906 119856 239912
rect 118712 219406 119660 219434
rect 118712 204950 118740 219406
rect 118700 204944 118752 204950
rect 118700 204886 118752 204892
rect 117962 200696 118018 200705
rect 117962 200631 118018 200640
rect 115940 198076 115992 198082
rect 115940 198018 115992 198024
rect 111064 189848 111116 189854
rect 111064 189790 111116 189796
rect 118608 189168 118660 189174
rect 118608 189110 118660 189116
rect 109040 188420 109092 188426
rect 109040 188362 109092 188368
rect 107660 185836 107712 185842
rect 107660 185778 107712 185784
rect 114468 183660 114520 183666
rect 114468 183602 114520 183608
rect 112996 180940 113048 180946
rect 112996 180882 113048 180888
rect 110696 179512 110748 179518
rect 110696 179454 110748 179460
rect 109868 178288 109920 178294
rect 109868 178230 109920 178236
rect 100666 177576 100722 177585
rect 100666 177511 100722 177520
rect 102046 177576 102102 177585
rect 102046 177511 102102 177520
rect 106186 177576 106242 177585
rect 106186 177511 106242 177520
rect 107566 177576 107622 177585
rect 107566 177511 107622 177520
rect 108120 177064 108172 177070
rect 108120 177006 108172 177012
rect 97814 176896 97870 176905
rect 97814 176831 97870 176840
rect 108132 176769 108160 177006
rect 109880 176769 109908 178230
rect 110708 177177 110736 179454
rect 113008 177585 113036 180882
rect 113916 179580 113968 179586
rect 113916 179522 113968 179528
rect 112994 177576 113050 177585
rect 112994 177511 113050 177520
rect 113928 177177 113956 179522
rect 114480 177585 114508 183602
rect 116952 181008 117004 181014
rect 116952 180950 117004 180956
rect 116964 177585 116992 180950
rect 118620 177585 118648 189110
rect 119712 178016 119764 178022
rect 119712 177958 119764 177964
rect 114466 177576 114522 177585
rect 114466 177511 114522 177520
rect 116950 177576 117006 177585
rect 116950 177511 117006 177520
rect 118606 177576 118662 177585
rect 118606 177511 118662 177520
rect 110694 177168 110750 177177
rect 110694 177103 110750 177112
rect 113914 177168 113970 177177
rect 113914 177103 113970 177112
rect 119724 176769 119752 177958
rect 120092 177342 120120 241431
rect 120184 224262 120212 250951
rect 120736 245002 120764 296686
rect 120816 289876 120868 289882
rect 120816 289818 120868 289824
rect 120724 244996 120776 245002
rect 120724 244938 120776 244944
rect 120828 238814 120856 289818
rect 121472 287054 121500 312734
rect 121552 311160 121604 311166
rect 121552 311102 121604 311108
rect 121564 292534 121592 311102
rect 121552 292528 121604 292534
rect 121552 292470 121604 292476
rect 121564 291825 121592 292470
rect 121550 291816 121606 291825
rect 121550 291751 121606 291760
rect 121642 291136 121698 291145
rect 121642 291071 121698 291080
rect 121550 290456 121606 290465
rect 121550 290391 121606 290400
rect 121564 289950 121592 290391
rect 121656 290018 121684 291071
rect 121644 290012 121696 290018
rect 121644 289954 121696 289960
rect 121552 289944 121604 289950
rect 121552 289886 121604 289892
rect 121552 289808 121604 289814
rect 121550 289776 121552 289785
rect 121604 289776 121606 289785
rect 121550 289711 121606 289720
rect 121550 289096 121606 289105
rect 121550 289031 121606 289040
rect 121564 288454 121592 289031
rect 121552 288448 121604 288454
rect 121552 288390 121604 288396
rect 121734 288416 121790 288425
rect 121644 288380 121696 288386
rect 121734 288351 121790 288360
rect 121644 288322 121696 288328
rect 121656 287745 121684 288322
rect 121642 287736 121698 287745
rect 121642 287671 121698 287680
rect 121748 287094 121776 288351
rect 121736 287088 121788 287094
rect 121472 287026 121684 287054
rect 122760 287065 122788 373254
rect 128360 371272 128412 371278
rect 128360 371214 128412 371220
rect 124864 365764 124916 365770
rect 124864 365706 124916 365712
rect 124128 340944 124180 340950
rect 124128 340886 124180 340892
rect 123484 297016 123536 297022
rect 123484 296958 123536 296964
rect 121736 287030 121788 287036
rect 122746 287056 122802 287065
rect 121460 286476 121512 286482
rect 121460 286418 121512 286424
rect 121472 285705 121500 286418
rect 121458 285696 121514 285705
rect 121458 285631 121514 285640
rect 121552 285660 121604 285666
rect 121552 285602 121604 285608
rect 121458 285016 121514 285025
rect 121458 284951 121514 284960
rect 121472 284374 121500 284951
rect 121460 284368 121512 284374
rect 121564 284345 121592 285602
rect 121460 284310 121512 284316
rect 121550 284336 121606 284345
rect 121550 284271 121606 284280
rect 121458 283656 121514 283665
rect 121458 283591 121514 283600
rect 121472 282946 121500 283591
rect 121460 282940 121512 282946
rect 121460 282882 121512 282888
rect 121550 282296 121606 282305
rect 121550 282231 121606 282240
rect 121564 281654 121592 282231
rect 121552 281648 121604 281654
rect 121458 281616 121514 281625
rect 121552 281590 121604 281596
rect 121458 281551 121460 281560
rect 121512 281551 121514 281560
rect 121460 281522 121512 281528
rect 121550 280936 121606 280945
rect 121550 280871 121606 280880
rect 121564 280294 121592 280871
rect 121552 280288 121604 280294
rect 121458 280256 121514 280265
rect 121552 280230 121604 280236
rect 121458 280191 121460 280200
rect 121512 280191 121514 280200
rect 121460 280162 121512 280168
rect 121458 278896 121514 278905
rect 121458 278831 121514 278840
rect 121472 278798 121500 278831
rect 121460 278792 121512 278798
rect 121460 278734 121512 278740
rect 121458 277536 121514 277545
rect 121458 277471 121514 277480
rect 121472 277438 121500 277471
rect 121460 277432 121512 277438
rect 121460 277374 121512 277380
rect 121550 276856 121606 276865
rect 121550 276791 121606 276800
rect 121458 276176 121514 276185
rect 121564 276146 121592 276791
rect 121458 276111 121514 276120
rect 121552 276140 121604 276146
rect 121472 276078 121500 276111
rect 121552 276082 121604 276088
rect 121460 276072 121512 276078
rect 121460 276014 121512 276020
rect 121550 275496 121606 275505
rect 121550 275431 121606 275440
rect 121458 274816 121514 274825
rect 121458 274751 121460 274760
rect 121512 274751 121514 274760
rect 121460 274722 121512 274728
rect 121564 274718 121592 275431
rect 121552 274712 121604 274718
rect 121552 274654 121604 274660
rect 121460 274440 121512 274446
rect 121460 274382 121512 274388
rect 121472 274145 121500 274382
rect 121458 274136 121514 274145
rect 121458 274071 121514 274080
rect 121458 273456 121514 273465
rect 121458 273391 121514 273400
rect 121472 273290 121500 273391
rect 121460 273284 121512 273290
rect 121460 273226 121512 273232
rect 121656 272785 121684 287026
rect 122746 286991 122802 287000
rect 122760 286414 122788 286991
rect 122748 286408 122800 286414
rect 122748 286350 122800 286356
rect 121734 282976 121790 282985
rect 121734 282911 121790 282920
rect 121748 278050 121776 282911
rect 122286 279576 122342 279585
rect 122286 279511 122342 279520
rect 122194 278216 122250 278225
rect 122194 278151 122250 278160
rect 121736 278044 121788 278050
rect 121736 277986 121788 277992
rect 121642 272776 121698 272785
rect 121642 272711 121698 272720
rect 122102 272776 122158 272785
rect 122102 272711 122158 272720
rect 120908 272536 120960 272542
rect 120908 272478 120960 272484
rect 120816 238808 120868 238814
rect 120816 238750 120868 238756
rect 120920 238542 120948 272478
rect 121458 272096 121514 272105
rect 121458 272031 121514 272040
rect 121472 271930 121500 272031
rect 121460 271924 121512 271930
rect 121460 271866 121512 271872
rect 121458 271416 121514 271425
rect 121458 271351 121514 271360
rect 121472 270570 121500 271351
rect 121460 270564 121512 270570
rect 121460 270506 121512 270512
rect 121550 270056 121606 270065
rect 121550 269991 121606 270000
rect 121458 269376 121514 269385
rect 121458 269311 121514 269320
rect 121472 269210 121500 269311
rect 121460 269204 121512 269210
rect 121460 269146 121512 269152
rect 121564 269142 121592 269991
rect 121552 269136 121604 269142
rect 121552 269078 121604 269084
rect 121458 268016 121514 268025
rect 121458 267951 121514 267960
rect 121472 267850 121500 267951
rect 121460 267844 121512 267850
rect 121460 267786 121512 267792
rect 121550 267336 121606 267345
rect 121550 267271 121606 267280
rect 121458 266656 121514 266665
rect 121458 266591 121514 266600
rect 121472 266422 121500 266591
rect 121564 266490 121592 267271
rect 121552 266484 121604 266490
rect 121552 266426 121604 266432
rect 121460 266416 121512 266422
rect 121460 266358 121512 266364
rect 121550 265976 121606 265985
rect 121550 265911 121606 265920
rect 121458 265296 121514 265305
rect 121458 265231 121514 265240
rect 121472 264994 121500 265231
rect 121564 265062 121592 265911
rect 121552 265056 121604 265062
rect 121552 264998 121604 265004
rect 121460 264988 121512 264994
rect 121460 264930 121512 264936
rect 121550 263936 121606 263945
rect 121550 263871 121606 263880
rect 121564 263634 121592 263871
rect 121552 263628 121604 263634
rect 121552 263570 121604 263576
rect 121460 263560 121512 263566
rect 121460 263502 121512 263508
rect 121472 263265 121500 263502
rect 121458 263256 121514 263265
rect 121458 263191 121514 263200
rect 121458 262576 121514 262585
rect 121458 262511 121514 262520
rect 121472 262274 121500 262511
rect 121460 262268 121512 262274
rect 121460 262210 121512 262216
rect 121552 262200 121604 262206
rect 121552 262142 121604 262148
rect 121564 261225 121592 262142
rect 121642 261896 121698 261905
rect 121642 261831 121698 261840
rect 121550 261216 121606 261225
rect 121550 261151 121606 261160
rect 121656 260914 121684 261831
rect 121644 260908 121696 260914
rect 121644 260850 121696 260856
rect 121460 260840 121512 260846
rect 121460 260782 121512 260788
rect 121472 260545 121500 260782
rect 121458 260536 121514 260545
rect 121458 260471 121514 260480
rect 121458 259856 121514 259865
rect 121458 259791 121514 259800
rect 121472 259486 121500 259791
rect 121460 259480 121512 259486
rect 121460 259422 121512 259428
rect 121458 259176 121514 259185
rect 121458 259111 121514 259120
rect 121472 258126 121500 259111
rect 121460 258120 121512 258126
rect 121460 258062 121512 258068
rect 121550 257816 121606 257825
rect 121550 257751 121606 257760
rect 121458 257136 121514 257145
rect 121458 257071 121514 257080
rect 121472 256766 121500 257071
rect 121564 256834 121592 257751
rect 121552 256828 121604 256834
rect 121552 256770 121604 256776
rect 121460 256760 121512 256766
rect 121460 256702 121512 256708
rect 122116 256018 122144 272711
rect 122104 256012 122156 256018
rect 122104 255954 122156 255960
rect 120998 255912 121054 255921
rect 120998 255847 121054 255856
rect 121012 255377 121040 255847
rect 120998 255368 121054 255377
rect 120998 255303 121054 255312
rect 122102 255096 122158 255105
rect 122102 255031 122158 255040
rect 121458 254416 121514 254425
rect 121458 254351 121514 254360
rect 121472 253978 121500 254351
rect 121460 253972 121512 253978
rect 121460 253914 121512 253920
rect 121550 253736 121606 253745
rect 121550 253671 121606 253680
rect 121458 253056 121514 253065
rect 121458 252991 121514 253000
rect 121472 252618 121500 252991
rect 121564 252686 121592 253671
rect 121552 252680 121604 252686
rect 121552 252622 121604 252628
rect 121460 252612 121512 252618
rect 121460 252554 121512 252560
rect 121458 251696 121514 251705
rect 121458 251631 121514 251640
rect 121472 251258 121500 251631
rect 121460 251252 121512 251258
rect 121460 251194 121512 251200
rect 121458 250336 121514 250345
rect 121458 250271 121514 250280
rect 121472 249830 121500 250271
rect 121460 249824 121512 249830
rect 121460 249766 121512 249772
rect 121550 249656 121606 249665
rect 121550 249591 121606 249600
rect 121458 248976 121514 248985
rect 121458 248911 121514 248920
rect 121472 248470 121500 248911
rect 121564 248538 121592 249591
rect 121552 248532 121604 248538
rect 121552 248474 121604 248480
rect 121460 248464 121512 248470
rect 121460 248406 121512 248412
rect 121552 248396 121604 248402
rect 121552 248338 121604 248344
rect 121458 248296 121514 248305
rect 121458 248231 121514 248240
rect 121472 247110 121500 248231
rect 121564 248033 121592 248338
rect 121550 248024 121606 248033
rect 121550 247959 121606 247968
rect 121460 247104 121512 247110
rect 121460 247046 121512 247052
rect 121550 246936 121606 246945
rect 121550 246871 121606 246880
rect 121458 246256 121514 246265
rect 121458 246191 121514 246200
rect 121472 245750 121500 246191
rect 121460 245744 121512 245750
rect 121460 245686 121512 245692
rect 121564 245682 121592 246871
rect 121552 245676 121604 245682
rect 121552 245618 121604 245624
rect 121460 245608 121512 245614
rect 121460 245550 121512 245556
rect 121550 245576 121606 245585
rect 121472 244905 121500 245550
rect 121550 245511 121606 245520
rect 121458 244896 121514 244905
rect 121458 244831 121514 244840
rect 121564 244322 121592 245511
rect 121552 244316 121604 244322
rect 121552 244258 121604 244264
rect 121550 244216 121606 244225
rect 121550 244151 121606 244160
rect 121458 243536 121514 243545
rect 121458 243471 121514 243480
rect 121472 242962 121500 243471
rect 121564 243030 121592 244151
rect 121552 243024 121604 243030
rect 121552 242966 121604 242972
rect 121460 242956 121512 242962
rect 121460 242898 121512 242904
rect 121552 242888 121604 242894
rect 121458 242856 121514 242865
rect 121552 242830 121604 242836
rect 121458 242791 121460 242800
rect 121512 242791 121514 242800
rect 121460 242762 121512 242768
rect 121564 242185 121592 242830
rect 121550 242176 121606 242185
rect 121550 242111 121606 242120
rect 121458 240816 121514 240825
rect 121458 240751 121514 240760
rect 121472 240174 121500 240751
rect 121460 240168 121512 240174
rect 121460 240110 121512 240116
rect 121550 240136 121606 240145
rect 121550 240071 121606 240080
rect 121564 239018 121592 240071
rect 121552 239012 121604 239018
rect 121552 238954 121604 238960
rect 120908 238536 120960 238542
rect 120908 238478 120960 238484
rect 120172 224256 120224 224262
rect 120172 224198 120224 224204
rect 122116 203726 122144 255031
rect 122208 237969 122236 278151
rect 122300 267734 122328 279511
rect 122300 267706 122512 267734
rect 122484 254590 122512 267706
rect 122472 254584 122524 254590
rect 122472 254526 122524 254532
rect 122194 237960 122250 237969
rect 122194 237895 122250 237904
rect 122104 203720 122156 203726
rect 122104 203662 122156 203668
rect 123496 196790 123524 296958
rect 123668 292664 123720 292670
rect 123668 292606 123720 292612
rect 123576 286340 123628 286346
rect 123576 286282 123628 286288
rect 123588 235890 123616 286282
rect 123680 266354 123708 292606
rect 124140 286482 124168 340886
rect 124128 286476 124180 286482
rect 124128 286418 124180 286424
rect 124876 274446 124904 365706
rect 126244 360460 126296 360466
rect 126244 360402 126296 360408
rect 124956 299872 125008 299878
rect 124956 299814 125008 299820
rect 124864 274440 124916 274446
rect 124864 274382 124916 274388
rect 123668 266348 123720 266354
rect 123668 266290 123720 266296
rect 123576 235884 123628 235890
rect 123576 235826 123628 235832
rect 124968 211954 124996 299814
rect 125048 294228 125100 294234
rect 125048 294170 125100 294176
rect 125060 242214 125088 294170
rect 125138 292768 125194 292777
rect 125138 292703 125194 292712
rect 125152 284209 125180 292703
rect 125138 284200 125194 284209
rect 125138 284135 125194 284144
rect 125048 242208 125100 242214
rect 125048 242150 125100 242156
rect 126256 238474 126284 360402
rect 127716 347812 127768 347818
rect 127716 347754 127768 347760
rect 126336 295656 126388 295662
rect 126336 295598 126388 295604
rect 126244 238468 126296 238474
rect 126244 238410 126296 238416
rect 124956 211948 125008 211954
rect 124956 211890 125008 211896
rect 126348 198218 126376 295598
rect 126428 294364 126480 294370
rect 126428 294306 126480 294312
rect 126440 207738 126468 294306
rect 127624 291372 127676 291378
rect 127624 291314 127676 291320
rect 126428 207732 126480 207738
rect 126428 207674 126480 207680
rect 126336 198212 126388 198218
rect 126336 198154 126388 198160
rect 123484 196784 123536 196790
rect 123484 196726 123536 196732
rect 127636 192642 127664 291314
rect 127728 251190 127756 347754
rect 128372 273222 128400 371214
rect 130384 363044 130436 363050
rect 130384 362986 130436 362992
rect 129188 311976 129240 311982
rect 129188 311918 129240 311924
rect 129004 295724 129056 295730
rect 129004 295666 129056 295672
rect 128360 273216 128412 273222
rect 128360 273158 128412 273164
rect 128372 272542 128400 273158
rect 128360 272536 128412 272542
rect 128360 272478 128412 272484
rect 127808 265056 127860 265062
rect 127808 264998 127860 265004
rect 127716 251184 127768 251190
rect 127716 251126 127768 251132
rect 127820 240854 127848 264998
rect 127808 240848 127860 240854
rect 127808 240790 127860 240796
rect 127624 192636 127676 192642
rect 127624 192578 127676 192584
rect 128268 183592 128320 183598
rect 128268 183534 128320 183540
rect 127808 182232 127860 182238
rect 127808 182174 127860 182180
rect 122012 178152 122064 178158
rect 122012 178094 122064 178100
rect 120080 177336 120132 177342
rect 120080 177278 120132 177284
rect 122024 176769 122052 178094
rect 124956 178084 125008 178090
rect 124956 178026 125008 178032
rect 123024 176928 123076 176934
rect 123024 176870 123076 176876
rect 123036 176769 123064 176870
rect 124968 176769 124996 178026
rect 127820 177585 127848 182174
rect 127806 177576 127862 177585
rect 127806 177511 127862 177520
rect 125876 176860 125928 176866
rect 125876 176802 125928 176808
rect 125888 176769 125916 176802
rect 128280 176769 128308 183534
rect 129016 178770 129044 295666
rect 129096 278792 129148 278798
rect 129096 278734 129148 278740
rect 129108 187202 129136 278734
rect 129200 234530 129228 311918
rect 129280 295520 129332 295526
rect 129280 295462 129332 295468
rect 129292 280158 129320 295462
rect 129280 280152 129332 280158
rect 129280 280094 129332 280100
rect 129280 262268 129332 262274
rect 129280 262210 129332 262216
rect 129188 234524 129240 234530
rect 129188 234466 129240 234472
rect 129292 224398 129320 262210
rect 130396 231742 130424 362986
rect 134524 361684 134576 361690
rect 134524 361626 134576 361632
rect 130568 325712 130620 325718
rect 130568 325654 130620 325660
rect 130476 299804 130528 299810
rect 130476 299746 130528 299752
rect 130384 231736 130436 231742
rect 130384 231678 130436 231684
rect 129280 224392 129332 224398
rect 129280 224334 129332 224340
rect 129188 224324 129240 224330
rect 129188 224266 129240 224272
rect 129200 194138 129228 224266
rect 129188 194132 129240 194138
rect 129188 194074 129240 194080
rect 129096 187196 129148 187202
rect 129096 187138 129148 187144
rect 130488 181529 130516 299746
rect 130580 238678 130608 325654
rect 133144 301096 133196 301102
rect 133144 301038 133196 301044
rect 131854 298208 131910 298217
rect 131854 298143 131910 298152
rect 131764 294296 131816 294302
rect 131764 294238 131816 294244
rect 130660 249824 130712 249830
rect 130660 249766 130712 249772
rect 130568 238672 130620 238678
rect 130568 238614 130620 238620
rect 130672 196994 130700 249766
rect 131776 200870 131804 294238
rect 131868 222902 131896 298143
rect 131856 222896 131908 222902
rect 131856 222838 131908 222844
rect 131764 200864 131816 200870
rect 131764 200806 131816 200812
rect 130660 196988 130712 196994
rect 130660 196930 130712 196936
rect 133156 192506 133184 301038
rect 133236 298308 133288 298314
rect 133236 298250 133288 298256
rect 133248 210594 133276 298250
rect 134536 237386 134564 361626
rect 135260 355360 135312 355366
rect 135260 355302 135312 355308
rect 135272 354754 135300 355302
rect 135260 354748 135312 354754
rect 135260 354690 135312 354696
rect 134616 296880 134668 296886
rect 134616 296822 134668 296828
rect 134524 237380 134576 237386
rect 134524 237322 134576 237328
rect 133236 210588 133288 210594
rect 133236 210530 133288 210536
rect 134628 195566 134656 296822
rect 134708 292800 134760 292806
rect 134708 292742 134760 292748
rect 134720 199345 134748 292742
rect 134800 267844 134852 267850
rect 134800 267786 134852 267792
rect 134812 215966 134840 267786
rect 135272 239426 135300 354690
rect 137284 299668 137336 299674
rect 137284 299610 137336 299616
rect 135904 298240 135956 298246
rect 135904 298182 135956 298188
rect 135260 239420 135312 239426
rect 135260 239362 135312 239368
rect 134800 215960 134852 215966
rect 134800 215902 134852 215908
rect 134706 199336 134762 199345
rect 134706 199271 134762 199280
rect 134616 195560 134668 195566
rect 134616 195502 134668 195508
rect 133144 192500 133196 192506
rect 133144 192442 133196 192448
rect 135916 191146 135944 298182
rect 135996 291440 136048 291446
rect 135996 291382 136048 291388
rect 135904 191140 135956 191146
rect 135904 191082 135956 191088
rect 133788 189100 133840 189106
rect 133788 189042 133840 189048
rect 130474 181520 130530 181529
rect 130474 181455 130530 181464
rect 129464 180872 129516 180878
rect 129464 180814 129516 180820
rect 129004 178764 129056 178770
rect 129004 178706 129056 178712
rect 129476 177585 129504 180814
rect 133800 177585 133828 189042
rect 136008 188494 136036 291382
rect 136088 286476 136140 286482
rect 136088 286418 136140 286424
rect 136100 224262 136128 286418
rect 136088 224256 136140 224262
rect 136088 224198 136140 224204
rect 137296 191282 137324 299610
rect 137376 280288 137428 280294
rect 137376 280230 137428 280236
rect 137388 192545 137416 280230
rect 138032 235929 138060 699774
rect 142804 365832 142856 365838
rect 142804 365774 142856 365780
rect 140136 356244 140188 356250
rect 140136 356186 140188 356192
rect 138112 311908 138164 311914
rect 138112 311850 138164 311856
rect 138124 307086 138152 311850
rect 138112 307080 138164 307086
rect 138112 307022 138164 307028
rect 138756 295588 138808 295594
rect 138756 295530 138808 295536
rect 138664 290012 138716 290018
rect 138664 289954 138716 289960
rect 138018 235920 138074 235929
rect 138018 235855 138074 235864
rect 137374 192536 137430 192545
rect 137374 192471 137430 192480
rect 137284 191276 137336 191282
rect 137284 191218 137336 191224
rect 138676 188562 138704 289954
rect 138768 217462 138796 295530
rect 140044 293276 140096 293282
rect 140044 293218 140096 293224
rect 138848 270564 138900 270570
rect 138848 270506 138900 270512
rect 138756 217456 138808 217462
rect 138756 217398 138808 217404
rect 138860 209234 138888 270506
rect 138848 209228 138900 209234
rect 138848 209170 138900 209176
rect 138664 188556 138716 188562
rect 138664 188498 138716 188504
rect 135996 188488 136048 188494
rect 135996 188430 136048 188436
rect 134524 184952 134576 184958
rect 134524 184894 134576 184900
rect 134536 178022 134564 184894
rect 140056 181694 140084 293218
rect 140148 248402 140176 356186
rect 140228 306400 140280 306406
rect 140228 306342 140280 306348
rect 140136 248396 140188 248402
rect 140136 248338 140188 248344
rect 140240 240786 140268 306342
rect 141514 294128 141570 294137
rect 141514 294063 141570 294072
rect 141424 292868 141476 292874
rect 141424 292810 141476 292816
rect 140320 256828 140372 256834
rect 140320 256770 140372 256776
rect 140228 240780 140280 240786
rect 140228 240722 140280 240728
rect 140332 198150 140360 256770
rect 140320 198144 140372 198150
rect 140320 198086 140372 198092
rect 141436 189922 141464 292810
rect 141528 236706 141556 294063
rect 141516 236700 141568 236706
rect 141516 236642 141568 236648
rect 142816 235822 142844 365774
rect 144184 359100 144236 359106
rect 144184 359042 144236 359048
rect 143080 301028 143132 301034
rect 143080 300970 143132 300976
rect 142896 300960 142948 300966
rect 142896 300902 142948 300908
rect 142804 235816 142856 235822
rect 142804 235758 142856 235764
rect 142908 199578 142936 300902
rect 143092 246362 143120 300970
rect 143172 273284 143224 273290
rect 143172 273226 143224 273232
rect 143080 246356 143132 246362
rect 143080 246298 143132 246304
rect 142988 245744 143040 245750
rect 142988 245686 143040 245692
rect 142896 199572 142948 199578
rect 142896 199514 142948 199520
rect 143000 191418 143028 245686
rect 143184 242282 143212 273226
rect 143172 242276 143224 242282
rect 143172 242218 143224 242224
rect 144196 237318 144224 359042
rect 150346 357912 150402 357921
rect 150346 357847 150402 357856
rect 148324 357604 148376 357610
rect 148324 357546 148376 357552
rect 147036 305108 147088 305114
rect 147036 305050 147088 305056
rect 146944 303680 146996 303686
rect 146944 303622 146996 303628
rect 145656 298444 145708 298450
rect 145656 298386 145708 298392
rect 144368 296948 144420 296954
rect 144368 296890 144420 296896
rect 144276 289944 144328 289950
rect 144276 289886 144328 289892
rect 144184 237312 144236 237318
rect 144184 237254 144236 237260
rect 144288 214810 144316 289886
rect 144380 241233 144408 296890
rect 145564 287088 145616 287094
rect 145564 287030 145616 287036
rect 144552 247104 144604 247110
rect 144552 247046 144604 247052
rect 144366 241224 144422 241233
rect 144366 241159 144422 241168
rect 144460 240168 144512 240174
rect 144460 240110 144512 240116
rect 144276 214804 144328 214810
rect 144276 214746 144328 214752
rect 142988 191412 143040 191418
rect 142988 191354 143040 191360
rect 144472 189990 144500 240110
rect 144564 210526 144592 247046
rect 144552 210520 144604 210526
rect 144552 210462 144604 210468
rect 145576 202230 145604 287030
rect 145668 217598 145696 298386
rect 145748 269204 145800 269210
rect 145748 269146 145800 269152
rect 145656 217592 145708 217598
rect 145656 217534 145708 217540
rect 145760 206417 145788 269146
rect 145746 206408 145802 206417
rect 145746 206343 145802 206352
rect 146956 202434 146984 303622
rect 147048 245070 147076 305050
rect 147128 295384 147180 295390
rect 147128 295326 147180 295332
rect 147036 245064 147088 245070
rect 147036 245006 147088 245012
rect 147036 243024 147088 243030
rect 147036 242966 147088 242972
rect 146944 202428 146996 202434
rect 146944 202370 146996 202376
rect 145564 202224 145616 202230
rect 145564 202166 145616 202172
rect 144460 189984 144512 189990
rect 144460 189926 144512 189932
rect 141424 189916 141476 189922
rect 141424 189858 141476 189864
rect 140044 181688 140096 181694
rect 140044 181630 140096 181636
rect 147048 181490 147076 242966
rect 147140 242758 147168 295326
rect 147220 276140 147272 276146
rect 147220 276082 147272 276088
rect 147128 242752 147180 242758
rect 147128 242694 147180 242700
rect 147128 238128 147180 238134
rect 147128 238070 147180 238076
rect 147140 194002 147168 238070
rect 147232 224874 147260 276082
rect 148336 238406 148364 357546
rect 149704 303748 149756 303754
rect 149704 303690 149756 303696
rect 148416 294024 148468 294030
rect 148416 293966 148468 293972
rect 148324 238400 148376 238406
rect 148324 238342 148376 238348
rect 147220 224868 147272 224874
rect 147220 224810 147272 224816
rect 147128 193996 147180 194002
rect 147128 193938 147180 193944
rect 148428 187270 148456 293966
rect 148508 288448 148560 288454
rect 148508 288390 148560 288396
rect 148416 187264 148468 187270
rect 148416 187206 148468 187212
rect 148520 182918 148548 288390
rect 148600 263628 148652 263634
rect 148600 263570 148652 263576
rect 148612 217530 148640 263570
rect 148600 217524 148652 217530
rect 148600 217466 148652 217472
rect 149716 213382 149744 303690
rect 149888 277432 149940 277438
rect 149888 277374 149940 277380
rect 149796 245676 149848 245682
rect 149796 245618 149848 245624
rect 149704 213376 149756 213382
rect 149704 213318 149756 213324
rect 149808 191350 149836 245618
rect 149900 234054 149928 277374
rect 149888 234048 149940 234054
rect 149888 233990 149940 233996
rect 150360 219434 150388 357847
rect 153212 356726 153240 702406
rect 170324 700330 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 177948 702568 178000 702574
rect 177948 702510 178000 702516
rect 170312 700324 170364 700330
rect 170312 700266 170364 700272
rect 158628 563100 158680 563106
rect 158628 563042 158680 563048
rect 157248 359032 157300 359038
rect 157248 358974 157300 358980
rect 154028 357400 154080 357406
rect 154028 357342 154080 357348
rect 154040 356726 154068 357342
rect 153200 356720 153252 356726
rect 153200 356662 153252 356668
rect 154028 356720 154080 356726
rect 154028 356662 154080 356668
rect 155406 300928 155462 300937
rect 155406 300863 155462 300872
rect 153936 299736 153988 299742
rect 153936 299678 153988 299684
rect 151084 298376 151136 298382
rect 151084 298318 151136 298324
rect 150348 219428 150400 219434
rect 150348 219370 150400 219376
rect 150360 218754 150388 219370
rect 150348 218748 150400 218754
rect 150348 218690 150400 218696
rect 151096 198014 151124 298318
rect 151268 298172 151320 298178
rect 151268 298114 151320 298120
rect 151176 274780 151228 274786
rect 151176 274722 151228 274728
rect 151188 207874 151216 274722
rect 151280 234530 151308 298114
rect 153844 297084 153896 297090
rect 153844 297026 153896 297032
rect 152464 294160 152516 294166
rect 152464 294102 152516 294108
rect 152476 278118 152504 294102
rect 152648 291304 152700 291310
rect 152648 291246 152700 291252
rect 152554 289232 152610 289241
rect 152554 289167 152610 289176
rect 152464 278112 152516 278118
rect 152464 278054 152516 278060
rect 152464 266484 152516 266490
rect 152464 266426 152516 266432
rect 151268 234524 151320 234530
rect 151268 234466 151320 234472
rect 151176 207868 151228 207874
rect 151176 207810 151228 207816
rect 151084 198008 151136 198014
rect 151084 197950 151136 197956
rect 149796 191344 149848 191350
rect 149796 191286 149848 191292
rect 152476 188426 152504 266426
rect 152568 235278 152596 289167
rect 152660 240106 152688 291246
rect 152740 242276 152792 242282
rect 152740 242218 152792 242224
rect 152648 240100 152700 240106
rect 152648 240042 152700 240048
rect 152556 235272 152608 235278
rect 152556 235214 152608 235220
rect 152752 213450 152780 242218
rect 152740 213444 152792 213450
rect 152740 213386 152792 213392
rect 153856 203862 153884 297026
rect 153948 218958 153976 299678
rect 154026 299568 154082 299577
rect 154026 299503 154082 299512
rect 154040 240825 154068 299503
rect 155224 271924 155276 271930
rect 155224 271866 155276 271872
rect 154120 242208 154172 242214
rect 154120 242150 154172 242156
rect 154026 240816 154082 240825
rect 154026 240751 154082 240760
rect 153936 218952 153988 218958
rect 153936 218894 153988 218900
rect 153844 203856 153896 203862
rect 153844 203798 153896 203804
rect 154132 192681 154160 242150
rect 154118 192672 154174 192681
rect 154118 192607 154174 192616
rect 152464 188420 152516 188426
rect 152464 188362 152516 188368
rect 148508 182912 148560 182918
rect 148508 182854 148560 182860
rect 147036 181484 147088 181490
rect 147036 181426 147088 181432
rect 148232 178220 148284 178226
rect 148232 178162 148284 178168
rect 134524 178016 134576 178022
rect 134524 177958 134576 177964
rect 129462 177576 129518 177585
rect 129462 177511 129518 177520
rect 133786 177576 133842 177585
rect 133786 177511 133842 177520
rect 132040 176996 132092 177002
rect 132040 176938 132092 176944
rect 132052 176769 132080 176938
rect 148244 176769 148272 178162
rect 108118 176760 108174 176769
rect 108118 176695 108174 176704
rect 109866 176760 109922 176769
rect 109866 176695 109922 176704
rect 119710 176760 119766 176769
rect 119710 176695 119766 176704
rect 122010 176760 122066 176769
rect 122010 176695 122066 176704
rect 123022 176760 123078 176769
rect 123022 176695 123078 176704
rect 124954 176760 125010 176769
rect 124954 176695 125010 176704
rect 125874 176760 125930 176769
rect 125874 176695 125930 176704
rect 128266 176760 128322 176769
rect 128266 176695 128322 176704
rect 132038 176760 132094 176769
rect 132038 176695 132094 176704
rect 134430 176760 134486 176769
rect 134430 176695 134432 176704
rect 134484 176695 134486 176704
rect 135718 176760 135774 176769
rect 135718 176695 135774 176704
rect 148230 176760 148286 176769
rect 148230 176695 148286 176704
rect 134432 176666 134484 176672
rect 135732 176662 135760 176695
rect 135720 176656 135772 176662
rect 135720 176598 135772 176604
rect 120816 176180 120868 176186
rect 120816 176122 120868 176128
rect 115756 176112 115808 176118
rect 115756 176054 115808 176060
rect 104624 176044 104676 176050
rect 104624 175986 104676 175992
rect 104636 175545 104664 175986
rect 104622 175536 104678 175545
rect 104622 175471 104678 175480
rect 115768 175001 115796 176054
rect 120828 175545 120856 176122
rect 130752 175976 130804 175982
rect 155236 175953 155264 271866
rect 155316 252680 155368 252686
rect 155316 252622 155368 252628
rect 155328 185910 155356 252622
rect 155420 238066 155448 300863
rect 156604 291236 156656 291242
rect 156604 291178 156656 291184
rect 155500 274712 155552 274718
rect 155500 274654 155552 274660
rect 155408 238060 155460 238066
rect 155408 238002 155460 238008
rect 155512 226302 155540 274654
rect 155500 226296 155552 226302
rect 155500 226238 155552 226244
rect 155316 185904 155368 185910
rect 155316 185846 155368 185852
rect 156616 181558 156644 291178
rect 156696 280220 156748 280226
rect 156696 280162 156748 280168
rect 156708 183122 156736 280162
rect 156788 240848 156840 240854
rect 156788 240790 156840 240796
rect 156800 225690 156828 240790
rect 156788 225684 156840 225690
rect 156788 225626 156840 225632
rect 157260 187338 157288 358974
rect 158536 307896 158588 307902
rect 158536 307838 158588 307844
rect 157984 299600 158036 299606
rect 157984 299542 158036 299548
rect 157340 298104 157392 298110
rect 157340 298046 157392 298052
rect 157352 297401 157380 298046
rect 157338 297392 157394 297401
rect 157338 297327 157394 297336
rect 157248 187332 157300 187338
rect 157248 187274 157300 187280
rect 156696 183116 156748 183122
rect 156696 183058 156748 183064
rect 156604 181552 156656 181558
rect 156604 181494 156656 181500
rect 157996 180130 158024 299542
rect 158076 244996 158128 245002
rect 158076 244938 158128 244944
rect 158088 195430 158116 244938
rect 158548 196625 158576 307838
rect 158640 298110 158668 563042
rect 166908 456816 166960 456822
rect 166908 456758 166960 456764
rect 160836 404388 160888 404394
rect 160836 404330 160888 404336
rect 160742 356144 160798 356153
rect 160742 356079 160798 356088
rect 160008 300824 160060 300830
rect 160008 300766 160060 300772
rect 160020 299538 160048 300766
rect 160008 299532 160060 299538
rect 160008 299474 160060 299480
rect 158628 298104 158680 298110
rect 158628 298046 158680 298052
rect 159364 296812 159416 296818
rect 159364 296754 159416 296760
rect 158628 294024 158680 294030
rect 158628 293966 158680 293972
rect 158640 242826 158668 293966
rect 158628 242820 158680 242826
rect 158628 242762 158680 242768
rect 159376 220250 159404 296754
rect 160020 262138 160048 299474
rect 160008 262132 160060 262138
rect 160008 262074 160060 262080
rect 160008 259548 160060 259554
rect 160008 259490 160060 259496
rect 159456 256760 159508 256766
rect 159456 256702 159508 256708
rect 159468 235890 159496 256702
rect 159456 235884 159508 235890
rect 159456 235826 159508 235832
rect 159548 235340 159600 235346
rect 159548 235282 159600 235288
rect 159364 220244 159416 220250
rect 159364 220186 159416 220192
rect 159560 216102 159588 235282
rect 159548 216096 159600 216102
rect 159548 216038 159600 216044
rect 160020 202298 160048 259490
rect 160756 242894 160784 356079
rect 160848 300830 160876 404330
rect 162768 360528 162820 360534
rect 162768 360470 162820 360476
rect 162122 354920 162178 354929
rect 162122 354855 162178 354864
rect 161572 334620 161624 334626
rect 161572 334562 161624 334568
rect 161584 330546 161612 334562
rect 161572 330540 161624 330546
rect 161572 330482 161624 330488
rect 160836 300824 160888 300830
rect 160836 300766 160888 300772
rect 160834 291952 160890 291961
rect 160834 291887 160890 291896
rect 160744 242888 160796 242894
rect 160744 242830 160796 242836
rect 160848 217394 160876 291887
rect 161388 267844 161440 267850
rect 161388 267786 161440 267792
rect 161020 248532 161072 248538
rect 161020 248474 161072 248480
rect 160928 242820 160980 242826
rect 160928 242762 160980 242768
rect 160940 223582 160968 242762
rect 161032 237318 161060 248474
rect 161020 237312 161072 237318
rect 161020 237254 161072 237260
rect 160928 223576 160980 223582
rect 160928 223518 160980 223524
rect 160744 217388 160796 217394
rect 160744 217330 160796 217336
rect 160836 217388 160888 217394
rect 160836 217330 160888 217336
rect 160756 206378 160784 217330
rect 160744 206372 160796 206378
rect 160744 206314 160796 206320
rect 160008 202292 160060 202298
rect 160008 202234 160060 202240
rect 158534 196616 158590 196625
rect 158534 196551 158590 196560
rect 158076 195424 158128 195430
rect 158076 195366 158128 195372
rect 161400 184385 161428 267786
rect 162136 245614 162164 354855
rect 162216 302252 162268 302258
rect 162216 302194 162268 302200
rect 162124 245608 162176 245614
rect 162124 245550 162176 245556
rect 162228 221678 162256 302194
rect 162676 278112 162728 278118
rect 162676 278054 162728 278060
rect 162688 277438 162716 278054
rect 162676 277432 162728 277438
rect 162676 277374 162728 277380
rect 162308 244928 162360 244934
rect 162308 244870 162360 244876
rect 162216 221672 162268 221678
rect 162216 221614 162268 221620
rect 162320 199510 162348 244870
rect 162688 228410 162716 277374
rect 162676 228404 162728 228410
rect 162676 228346 162728 228352
rect 162308 199504 162360 199510
rect 162308 199446 162360 199452
rect 161386 184376 161442 184385
rect 161386 184311 161442 184320
rect 162780 180334 162808 360470
rect 166264 314696 166316 314702
rect 166264 314638 166316 314644
rect 166276 311982 166304 314638
rect 166264 311976 166316 311982
rect 166264 311918 166316 311924
rect 164976 307828 165028 307834
rect 164976 307770 165028 307776
rect 163596 302320 163648 302326
rect 163596 302262 163648 302268
rect 163504 266416 163556 266422
rect 163504 266358 163556 266364
rect 163516 184414 163544 266358
rect 163608 221513 163636 302262
rect 164884 281648 164936 281654
rect 164884 281590 164936 281596
rect 163688 267776 163740 267782
rect 163688 267718 163740 267724
rect 163700 241466 163728 267718
rect 163688 241460 163740 241466
rect 163688 241402 163740 241408
rect 163688 228540 163740 228546
rect 163688 228482 163740 228488
rect 163594 221504 163650 221513
rect 163594 221439 163650 221448
rect 163700 214742 163728 228482
rect 163688 214736 163740 214742
rect 163688 214678 163740 214684
rect 163504 184408 163556 184414
rect 163504 184350 163556 184356
rect 162768 180328 162820 180334
rect 162768 180270 162820 180276
rect 157984 180124 158036 180130
rect 157984 180066 158036 180072
rect 162768 178288 162820 178294
rect 162768 178230 162820 178236
rect 158996 176792 159048 176798
rect 158994 176760 158996 176769
rect 159048 176760 159050 176769
rect 158994 176695 159050 176704
rect 162780 176254 162808 178230
rect 164896 177410 164924 281590
rect 164988 224330 165016 307770
rect 166276 306374 166304 311918
rect 166276 306346 166396 306374
rect 166264 292732 166316 292738
rect 166264 292674 166316 292680
rect 165068 269136 165120 269142
rect 165068 269078 165120 269084
rect 165080 228546 165108 269078
rect 165068 228540 165120 228546
rect 165068 228482 165120 228488
rect 164976 224324 165028 224330
rect 164976 224266 165028 224272
rect 166276 211993 166304 292674
rect 166368 237386 166396 306346
rect 166920 299470 166948 456758
rect 174728 361752 174780 361758
rect 174728 361694 174780 361700
rect 167644 360392 167696 360398
rect 167644 360334 167696 360340
rect 166448 299464 166500 299470
rect 166448 299406 166500 299412
rect 166908 299464 166960 299470
rect 166908 299406 166960 299412
rect 166460 298761 166488 299406
rect 166446 298752 166502 298761
rect 166446 298687 166502 298696
rect 167656 288386 167684 360334
rect 170404 360324 170456 360330
rect 170404 360266 170456 360272
rect 169024 355020 169076 355026
rect 169024 354962 169076 354968
rect 167736 295452 167788 295458
rect 167736 295394 167788 295400
rect 167644 288380 167696 288386
rect 167644 288322 167696 288328
rect 167748 282878 167776 295394
rect 168288 291236 168340 291242
rect 168288 291178 168340 291184
rect 167828 284368 167880 284374
rect 167828 284310 167880 284316
rect 167736 282872 167788 282878
rect 167736 282814 167788 282820
rect 167644 281580 167696 281586
rect 167644 281522 167696 281528
rect 166540 276072 166592 276078
rect 166540 276014 166592 276020
rect 166448 251252 166500 251258
rect 166448 251194 166500 251200
rect 166356 237380 166408 237386
rect 166356 237322 166408 237328
rect 166262 211984 166318 211993
rect 166262 211919 166318 211928
rect 166356 179580 166408 179586
rect 166356 179522 166408 179528
rect 166264 179512 166316 179518
rect 166264 179454 166316 179460
rect 164884 177404 164936 177410
rect 164884 177346 164936 177352
rect 165252 177064 165304 177070
rect 165252 177006 165304 177012
rect 162768 176248 162820 176254
rect 162768 176190 162820 176196
rect 130752 175918 130804 175924
rect 155222 175944 155278 175953
rect 130764 175545 130792 175918
rect 155222 175879 155278 175888
rect 120814 175536 120870 175545
rect 120814 175471 120870 175480
rect 130750 175536 130806 175545
rect 130750 175471 130806 175480
rect 115754 174992 115810 175001
rect 115754 174927 115810 174936
rect 67638 128072 67694 128081
rect 67638 128007 67694 128016
rect 67652 93809 67680 128007
rect 67730 100736 67786 100745
rect 67730 100671 67786 100680
rect 67638 93800 67694 93809
rect 67638 93735 67694 93744
rect 67546 91080 67602 91089
rect 67546 91015 67602 91024
rect 67456 89684 67508 89690
rect 67456 89626 67508 89632
rect 66076 89616 66128 89622
rect 66076 89558 66128 89564
rect 67744 86970 67772 100671
rect 165264 173194 165292 177006
rect 165436 176996 165488 177002
rect 165436 176938 165488 176944
rect 165448 174554 165476 176938
rect 165528 176928 165580 176934
rect 165528 176870 165580 176876
rect 165540 174593 165568 176870
rect 165526 174584 165582 174593
rect 165436 174548 165488 174554
rect 165526 174519 165582 174528
rect 165436 174490 165488 174496
rect 165252 173188 165304 173194
rect 165252 173130 165304 173136
rect 166276 162858 166304 179454
rect 166368 164218 166396 179522
rect 166460 177342 166488 251194
rect 166552 203794 166580 276014
rect 166540 203788 166592 203794
rect 166540 203730 166592 203736
rect 166540 181008 166592 181014
rect 166540 180950 166592 180956
rect 166448 177336 166500 177342
rect 166448 177278 166500 177284
rect 166448 176112 166500 176118
rect 166448 176054 166500 176060
rect 166460 165578 166488 176054
rect 166552 167006 166580 180950
rect 167656 178838 167684 281522
rect 167736 278044 167788 278050
rect 167736 277986 167788 277992
rect 167748 194070 167776 277986
rect 167840 231130 167868 284310
rect 167828 231124 167880 231130
rect 167828 231066 167880 231072
rect 167736 194064 167788 194070
rect 167736 194006 167788 194012
rect 167736 187808 167788 187814
rect 167736 187750 167788 187756
rect 167644 178832 167696 178838
rect 167644 178774 167696 178780
rect 167644 176180 167696 176186
rect 167644 176122 167696 176128
rect 167656 168366 167684 176122
rect 167644 168360 167696 168366
rect 167644 168302 167696 168308
rect 166540 167000 166592 167006
rect 166540 166942 166592 166948
rect 166448 165572 166500 165578
rect 166448 165514 166500 165520
rect 166356 164212 166408 164218
rect 166356 164154 166408 164160
rect 166264 162852 166316 162858
rect 166264 162794 166316 162800
rect 167748 160070 167776 187750
rect 167828 180940 167880 180946
rect 167828 180882 167880 180888
rect 167840 164150 167868 180882
rect 168300 177546 168328 291178
rect 169036 263566 169064 354962
rect 169024 263560 169076 263566
rect 169024 263502 169076 263508
rect 170416 260846 170444 360266
rect 174636 357740 174688 357746
rect 174636 357682 174688 357688
rect 174544 356380 174596 356386
rect 174544 356322 174596 356328
rect 171876 356312 171928 356318
rect 171876 356254 171928 356260
rect 171784 355088 171836 355094
rect 171784 355030 171836 355036
rect 170496 292596 170548 292602
rect 170496 292538 170548 292544
rect 170404 260840 170456 260846
rect 170404 260782 170456 260788
rect 169024 259480 169076 259486
rect 169024 259422 169076 259428
rect 168288 177540 168340 177546
rect 168288 177482 168340 177488
rect 169036 177478 169064 259422
rect 169208 256012 169260 256018
rect 169208 255954 169260 255960
rect 169116 254584 169168 254590
rect 169116 254526 169168 254532
rect 169128 180266 169156 254526
rect 169220 235822 169248 255954
rect 170404 253972 170456 253978
rect 170404 253914 170456 253920
rect 169208 235816 169260 235822
rect 169208 235758 169260 235764
rect 170416 219026 170444 253914
rect 170508 238542 170536 292538
rect 171796 262206 171824 355030
rect 171888 285666 171916 356254
rect 173808 321632 173860 321638
rect 173808 321574 173860 321580
rect 173164 309188 173216 309194
rect 173164 309130 173216 309136
rect 173176 302190 173204 309130
rect 173164 302184 173216 302190
rect 173164 302126 173216 302132
rect 172060 294092 172112 294098
rect 172060 294034 172112 294040
rect 171968 286408 172020 286414
rect 171968 286350 172020 286356
rect 171876 285660 171928 285666
rect 171876 285602 171928 285608
rect 171784 262200 171836 262206
rect 171784 262142 171836 262148
rect 170588 260908 170640 260914
rect 170588 260850 170640 260856
rect 170496 238536 170548 238542
rect 170496 238478 170548 238484
rect 170600 235414 170628 260850
rect 171876 258120 171928 258126
rect 171876 258062 171928 258068
rect 171784 245064 171836 245070
rect 171784 245006 171836 245012
rect 170680 244316 170732 244322
rect 170680 244258 170732 244264
rect 170588 235408 170640 235414
rect 170588 235350 170640 235356
rect 170692 229770 170720 244258
rect 170680 229764 170732 229770
rect 170680 229706 170732 229712
rect 170404 219020 170456 219026
rect 170404 218962 170456 218968
rect 170404 187740 170456 187746
rect 170404 187682 170456 187688
rect 169300 183660 169352 183666
rect 169300 183602 169352 183608
rect 169116 180260 169168 180266
rect 169116 180202 169168 180208
rect 169208 179444 169260 179450
rect 169208 179386 169260 179392
rect 169024 177472 169076 177478
rect 169024 177414 169076 177420
rect 169114 177032 169170 177041
rect 169114 176967 169170 176976
rect 167920 176860 167972 176866
rect 167920 176802 167972 176808
rect 167932 171086 167960 176802
rect 169024 176044 169076 176050
rect 169024 175986 169076 175992
rect 168010 171592 168066 171601
rect 168010 171527 168066 171536
rect 168024 171154 168052 171527
rect 168012 171148 168064 171154
rect 168012 171090 168064 171096
rect 167920 171080 167972 171086
rect 167920 171022 167972 171028
rect 167828 164144 167880 164150
rect 167828 164086 167880 164092
rect 167736 160064 167788 160070
rect 167736 160006 167788 160012
rect 169036 160002 169064 175986
rect 169128 169046 169156 176967
rect 169116 169040 169168 169046
rect 169116 168982 169168 168988
rect 169024 159996 169076 160002
rect 169024 159938 169076 159944
rect 169220 155922 169248 179386
rect 169312 165510 169340 183602
rect 169300 165504 169352 165510
rect 169300 165446 169352 165452
rect 170416 157350 170444 187682
rect 170494 175400 170550 175409
rect 170494 175335 170550 175344
rect 170404 157344 170456 157350
rect 170404 157286 170456 157292
rect 169208 155916 169260 155922
rect 169208 155858 169260 155864
rect 170508 155854 170536 175335
rect 170496 155848 170548 155854
rect 170496 155790 170548 155796
rect 167644 146328 167696 146334
rect 167644 146270 167696 146276
rect 166264 138032 166316 138038
rect 166264 137974 166316 137980
rect 165528 95940 165580 95946
rect 165528 95882 165580 95888
rect 102046 94752 102102 94761
rect 102046 94687 102102 94696
rect 113730 94752 113786 94761
rect 113730 94687 113786 94696
rect 115478 94752 115534 94761
rect 115478 94687 115534 94696
rect 133142 94752 133198 94761
rect 133142 94687 133198 94696
rect 102060 93906 102088 94687
rect 113744 94042 113772 94687
rect 113732 94036 113784 94042
rect 113732 93978 113784 93984
rect 115492 93974 115520 94687
rect 133156 94110 133184 94687
rect 133144 94104 133196 94110
rect 133144 94046 133196 94052
rect 115480 93968 115532 93974
rect 115480 93910 115532 93916
rect 102048 93900 102100 93906
rect 102048 93842 102100 93848
rect 134430 93664 134486 93673
rect 134430 93599 134486 93608
rect 151726 93664 151782 93673
rect 151726 93599 151782 93608
rect 110142 93528 110198 93537
rect 110142 93463 110198 93472
rect 118054 93528 118110 93537
rect 118054 93463 118110 93472
rect 119526 93528 119582 93537
rect 119526 93463 119582 93472
rect 110156 93226 110184 93463
rect 118068 93294 118096 93463
rect 118056 93288 118108 93294
rect 118056 93230 118108 93236
rect 110144 93220 110196 93226
rect 110144 93162 110196 93168
rect 119540 93158 119568 93463
rect 134444 93362 134472 93599
rect 151740 93430 151768 93599
rect 151728 93424 151780 93430
rect 151728 93366 151780 93372
rect 134432 93356 134484 93362
rect 134432 93298 134484 93304
rect 128174 93256 128230 93265
rect 128174 93191 128230 93200
rect 119528 93152 119580 93158
rect 119528 93094 119580 93100
rect 88984 92472 89036 92478
rect 74814 92440 74870 92449
rect 74814 92375 74870 92384
rect 85762 92440 85818 92449
rect 85762 92375 85818 92384
rect 88062 92440 88118 92449
rect 88062 92375 88118 92384
rect 88982 92440 88984 92449
rect 89036 92440 89038 92449
rect 88982 92375 89038 92384
rect 100574 92440 100630 92449
rect 100574 92375 100630 92384
rect 109222 92440 109278 92449
rect 109222 92375 109278 92384
rect 112166 92440 112222 92449
rect 112166 92375 112222 92384
rect 115478 92440 115534 92449
rect 115478 92375 115534 92384
rect 116766 92440 116822 92449
rect 116766 92375 116822 92384
rect 119710 92440 119766 92449
rect 119710 92375 119766 92384
rect 125874 92440 125930 92449
rect 125874 92375 125930 92384
rect 126518 92440 126574 92449
rect 126518 92375 126574 92384
rect 74828 91186 74856 92375
rect 85486 91216 85542 91225
rect 74816 91180 74868 91186
rect 85486 91151 85542 91160
rect 74816 91122 74868 91128
rect 67732 86964 67784 86970
rect 67732 86906 67784 86912
rect 73160 76560 73212 76566
rect 73160 76502 73212 76508
rect 63408 75880 63460 75886
rect 63408 75822 63460 75828
rect 64880 71052 64932 71058
rect 64880 70994 64932 71000
rect 53840 69692 53892 69698
rect 53840 69634 53892 69640
rect 49698 62792 49754 62801
rect 49698 62727 49754 62736
rect 49712 16574 49740 62727
rect 52460 24132 52512 24138
rect 52460 24074 52512 24080
rect 52472 16574 52500 24074
rect 53852 16574 53880 69634
rect 57980 68332 58032 68338
rect 57980 68274 58032 68280
rect 56598 55856 56654 55865
rect 56598 55791 56654 55800
rect 55220 26988 55272 26994
rect 55220 26930 55272 26936
rect 55232 16574 55260 26930
rect 56612 16574 56640 55791
rect 57992 16574 58020 68274
rect 63500 57248 63552 57254
rect 63500 57190 63552 57196
rect 62118 44840 62174 44849
rect 62118 44775 62174 44784
rect 60740 36644 60792 36650
rect 60740 36586 60792 36592
rect 60752 16574 60780 36586
rect 62132 16574 62160 44775
rect 63512 16574 63540 57190
rect 64892 16574 64920 70994
rect 69020 66904 69072 66910
rect 69020 66846 69072 66852
rect 67640 35216 67692 35222
rect 67640 35158 67692 35164
rect 66258 25528 66314 25537
rect 66258 25463 66314 25472
rect 66272 16574 66300 25463
rect 49712 16546 50200 16574
rect 52472 16546 53328 16574
rect 53852 16546 54984 16574
rect 55232 16546 56088 16574
rect 56612 16546 56824 16574
rect 57992 16546 58480 16574
rect 60752 16546 61608 16574
rect 62132 16546 63264 16574
rect 63512 16546 64368 16574
rect 64892 16546 65104 16574
rect 66272 16546 66760 16574
rect 48964 6860 49016 6866
rect 48964 6802 49016 6808
rect 48964 4820 49016 4826
rect 48964 4762 49016 4768
rect 48976 480 49004 4762
rect 50172 480 50200 16546
rect 51080 11824 51132 11830
rect 51080 11766 51132 11772
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 47830 -960 47942 326
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51092 354 51120 11766
rect 52550 4856 52606 4865
rect 52550 4791 52606 4800
rect 52564 480 52592 4791
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53300 354 53328 16546
rect 54956 480 54984 16546
rect 56060 480 56088 16546
rect 53718 354 53830 480
rect 53300 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 58452 480 58480 16546
rect 60832 3528 60884 3534
rect 60832 3470 60884 3476
rect 59636 2100 59688 2106
rect 59636 2042 59688 2048
rect 59648 480 59676 2042
rect 60844 480 60872 3470
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61580 354 61608 16546
rect 63236 480 63264 16546
rect 64340 480 64368 16546
rect 61998 354 62110 480
rect 61580 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66732 480 66760 16546
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 35158
rect 69032 6914 69060 66846
rect 71780 65544 71832 65550
rect 71780 65486 71832 65492
rect 70400 58676 70452 58682
rect 70400 58618 70452 58624
rect 69112 22840 69164 22846
rect 69112 22782 69164 22788
rect 69124 16574 69152 22782
rect 70412 16574 70440 58618
rect 71792 16574 71820 65486
rect 73172 16574 73200 76502
rect 77300 75268 77352 75274
rect 77300 75210 77352 75216
rect 74540 60104 74592 60110
rect 74540 60046 74592 60052
rect 74552 16574 74580 60046
rect 75920 18624 75972 18630
rect 75920 18566 75972 18572
rect 69124 16546 69888 16574
rect 70412 16546 71544 16574
rect 71792 16546 72648 16574
rect 73172 16546 73384 16574
rect 74552 16546 75040 16574
rect 69032 6886 69152 6914
rect 69124 480 69152 6886
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69860 354 69888 16546
rect 71516 480 71544 16546
rect 72620 480 72648 16546
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 16546
rect 75012 480 75040 16546
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 75932 354 75960 18566
rect 77312 3602 77340 75210
rect 81440 73908 81492 73914
rect 81440 73850 81492 73856
rect 78680 38004 78732 38010
rect 78680 37946 78732 37952
rect 78692 16574 78720 37946
rect 80060 19984 80112 19990
rect 80060 19926 80112 19932
rect 80072 16574 80100 19926
rect 81452 16574 81480 73850
rect 85500 73166 85528 91151
rect 85776 91118 85804 92375
rect 88076 91254 88104 92375
rect 99194 91488 99250 91497
rect 99194 91423 99250 91432
rect 95054 91352 95110 91361
rect 95054 91287 95110 91296
rect 97262 91352 97318 91361
rect 97262 91287 97318 91296
rect 99102 91352 99158 91361
rect 99102 91287 99158 91296
rect 88064 91248 88116 91254
rect 86866 91216 86922 91225
rect 88064 91190 88116 91196
rect 91006 91216 91062 91225
rect 86866 91151 86922 91160
rect 91006 91151 91062 91160
rect 92386 91216 92442 91225
rect 92386 91151 92442 91160
rect 93766 91216 93822 91225
rect 93766 91151 93822 91160
rect 85764 91112 85816 91118
rect 85764 91054 85816 91060
rect 86880 81326 86908 91151
rect 86868 81320 86920 81326
rect 86868 81262 86920 81268
rect 91020 74526 91048 91151
rect 92400 84182 92428 91151
rect 92388 84176 92440 84182
rect 92388 84118 92440 84124
rect 93780 77178 93808 91151
rect 95068 81394 95096 91287
rect 95146 91216 95202 91225
rect 95146 91151 95202 91160
rect 96158 91216 96214 91225
rect 96158 91151 96214 91160
rect 95056 81388 95108 81394
rect 95056 81330 95108 81336
rect 95160 80034 95188 91151
rect 96172 86873 96200 91151
rect 96158 86864 96214 86873
rect 96158 86799 96214 86808
rect 97276 85270 97304 91287
rect 97906 91216 97962 91225
rect 97906 91151 97962 91160
rect 97264 85264 97316 85270
rect 97264 85206 97316 85212
rect 95148 80028 95200 80034
rect 95148 79970 95200 79976
rect 97920 78674 97948 91151
rect 99116 84114 99144 91287
rect 99104 84108 99156 84114
rect 99104 84050 99156 84056
rect 99208 79762 99236 91423
rect 99286 91216 99342 91225
rect 100482 91216 100538 91225
rect 99286 91151 99342 91160
rect 100024 91180 100076 91186
rect 99196 79756 99248 79762
rect 99196 79698 99248 79704
rect 97908 78668 97960 78674
rect 97908 78610 97960 78616
rect 99300 78441 99328 91151
rect 100588 91186 100616 92375
rect 101862 91624 101918 91633
rect 101862 91559 101918 91568
rect 100482 91151 100538 91160
rect 100576 91180 100628 91186
rect 100024 91122 100076 91128
rect 99286 78432 99342 78441
rect 99286 78367 99342 78376
rect 100036 77246 100064 91122
rect 100496 88194 100524 91151
rect 100576 91122 100628 91128
rect 101876 89486 101904 91559
rect 107014 91352 107070 91361
rect 107014 91287 107070 91296
rect 102046 91216 102102 91225
rect 102046 91151 102102 91160
rect 103426 91216 103482 91225
rect 103426 91151 103482 91160
rect 104346 91216 104402 91225
rect 104346 91151 104402 91160
rect 104622 91216 104678 91225
rect 104622 91151 104678 91160
rect 105726 91216 105782 91225
rect 105726 91151 105782 91160
rect 106186 91216 106242 91225
rect 106186 91151 106242 91160
rect 101864 89480 101916 89486
rect 101864 89422 101916 89428
rect 100484 88188 100536 88194
rect 100484 88130 100536 88136
rect 102060 79830 102088 91151
rect 103440 84046 103468 91151
rect 104360 85338 104388 91151
rect 104636 85542 104664 91151
rect 104624 85536 104676 85542
rect 104624 85478 104676 85484
rect 105740 85406 105768 91151
rect 105728 85400 105780 85406
rect 105728 85342 105780 85348
rect 104348 85332 104400 85338
rect 104348 85274 104400 85280
rect 106200 84153 106228 91151
rect 107028 86737 107056 91287
rect 107566 91216 107622 91225
rect 107566 91151 107622 91160
rect 107842 91216 107898 91225
rect 107842 91151 107898 91160
rect 108946 91216 109002 91225
rect 108946 91151 109002 91160
rect 107014 86728 107070 86737
rect 107014 86663 107070 86672
rect 106186 84144 106242 84153
rect 106186 84079 106242 84088
rect 103428 84040 103480 84046
rect 103428 83982 103480 83988
rect 102048 79824 102100 79830
rect 102048 79766 102100 79772
rect 100024 77240 100076 77246
rect 100024 77182 100076 77188
rect 93768 77172 93820 77178
rect 93768 77114 93820 77120
rect 107580 75818 107608 91151
rect 107856 86834 107884 91151
rect 107844 86828 107896 86834
rect 107844 86770 107896 86776
rect 108960 82550 108988 91151
rect 109236 89554 109264 92375
rect 111064 91248 111116 91254
rect 110326 91216 110382 91225
rect 110326 91151 110382 91160
rect 110970 91216 111026 91225
rect 111064 91190 111116 91196
rect 111430 91216 111486 91225
rect 110970 91151 111026 91160
rect 109224 89548 109276 89554
rect 109224 89490 109276 89496
rect 110340 82686 110368 91151
rect 110984 88233 111012 91151
rect 110970 88224 111026 88233
rect 110970 88159 111026 88168
rect 110328 82680 110380 82686
rect 110328 82622 110380 82628
rect 108948 82544 109000 82550
rect 108948 82486 109000 82492
rect 107568 75812 107620 75818
rect 107568 75754 107620 75760
rect 103520 75200 103572 75206
rect 103520 75142 103572 75148
rect 91008 74520 91060 74526
rect 91008 74462 91060 74468
rect 85488 73160 85540 73166
rect 85488 73102 85540 73108
rect 85580 72480 85632 72486
rect 85580 72422 85632 72428
rect 82820 62824 82872 62830
rect 82820 62766 82872 62772
rect 82832 16574 82860 62766
rect 84200 28348 84252 28354
rect 84200 28290 84252 28296
rect 78692 16546 79272 16574
rect 80072 16546 80928 16574
rect 81452 16546 81664 16574
rect 82832 16546 83320 16574
rect 77392 14544 77444 14550
rect 77392 14486 77444 14492
rect 77300 3596 77352 3602
rect 77300 3538 77352 3544
rect 77404 480 77432 14486
rect 78220 3596 78272 3602
rect 78220 3538 78272 3544
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78232 354 78260 3538
rect 78558 354 78670 480
rect 78232 326 78670 354
rect 79244 354 79272 16546
rect 80900 480 80928 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83292 480 83320 16546
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 28290
rect 85592 16574 85620 72422
rect 88340 71120 88392 71126
rect 88340 71062 88392 71068
rect 86960 24200 87012 24206
rect 86960 24142 87012 24148
rect 86972 16574 87000 24142
rect 88352 16574 88380 71062
rect 92480 69760 92532 69766
rect 92480 69702 92532 69708
rect 89720 60036 89772 60042
rect 89720 59978 89772 59984
rect 89732 16574 89760 59978
rect 91100 21480 91152 21486
rect 91100 21422 91152 21428
rect 91112 16574 91140 21422
rect 85592 16546 85712 16574
rect 86972 16546 87552 16574
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 91112 16546 91600 16574
rect 85684 480 85712 16546
rect 86868 6180 86920 6186
rect 86868 6122 86920 6128
rect 86880 480 86908 6122
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87524 354 87552 16546
rect 89180 480 89208 16546
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 69702
rect 95240 68400 95292 68406
rect 95240 68342 95292 68348
rect 93860 58744 93912 58750
rect 93860 58686 93912 58692
rect 93872 6914 93900 58686
rect 93952 33856 94004 33862
rect 93952 33798 94004 33804
rect 93964 16574 93992 33798
rect 95252 16574 95280 68342
rect 99380 66972 99432 66978
rect 99380 66914 99432 66920
rect 96620 57316 96672 57322
rect 96620 57258 96672 57264
rect 96632 16574 96660 57258
rect 99392 16574 99420 66914
rect 100760 55888 100812 55894
rect 100760 55830 100812 55836
rect 93964 16546 94728 16574
rect 95252 16546 95832 16574
rect 96632 16546 97488 16574
rect 99392 16546 99880 16574
rect 93872 6886 93992 6914
rect 93964 480 93992 6886
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94700 354 94728 16546
rect 95118 354 95230 480
rect 94700 326 95230 354
rect 95804 354 95832 16546
rect 97460 480 97488 16546
rect 98184 11756 98236 11762
rect 98184 11698 98236 11704
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 11698
rect 99852 480 99880 16546
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 55830
rect 102140 29708 102192 29714
rect 102140 29650 102192 29656
rect 102152 6914 102180 29650
rect 102232 20052 102284 20058
rect 102232 19994 102284 20000
rect 102244 16574 102272 19994
rect 103532 16574 103560 75142
rect 111076 73098 111104 91190
rect 111430 91151 111486 91160
rect 111444 88262 111472 91151
rect 112180 90982 112208 92375
rect 113086 91216 113142 91225
rect 113086 91151 113142 91160
rect 114466 91216 114522 91225
rect 114466 91151 114522 91160
rect 112168 90976 112220 90982
rect 112168 90918 112220 90924
rect 111432 88256 111484 88262
rect 111432 88198 111484 88204
rect 113100 82618 113128 91151
rect 113088 82612 113140 82618
rect 113088 82554 113140 82560
rect 114480 81190 114508 91151
rect 115492 90914 115520 92375
rect 116780 92274 116808 92375
rect 116768 92268 116820 92274
rect 116768 92210 116820 92216
rect 119724 92138 119752 92375
rect 125888 92342 125916 92375
rect 125876 92336 125928 92342
rect 125876 92278 125928 92284
rect 119712 92132 119764 92138
rect 119712 92074 119764 92080
rect 122838 91488 122894 91497
rect 122838 91423 122894 91432
rect 122102 91352 122158 91361
rect 122102 91287 122158 91296
rect 115846 91216 115902 91225
rect 117226 91216 117282 91225
rect 115846 91151 115902 91160
rect 116584 91180 116636 91186
rect 115480 90908 115532 90914
rect 115480 90850 115532 90856
rect 115860 85202 115888 91151
rect 117226 91151 117282 91160
rect 118238 91216 118294 91225
rect 118238 91151 118294 91160
rect 120446 91216 120502 91225
rect 120446 91151 120502 91160
rect 121366 91216 121422 91225
rect 121366 91151 121422 91160
rect 116584 91122 116636 91128
rect 115848 85196 115900 85202
rect 115848 85138 115900 85144
rect 114468 81184 114520 81190
rect 114468 81126 114520 81132
rect 116596 79966 116624 91122
rect 117240 81258 117268 91151
rect 118252 86766 118280 91151
rect 118240 86760 118292 86766
rect 118240 86702 118292 86708
rect 120460 85474 120488 91151
rect 120448 85468 120500 85474
rect 120448 85410 120500 85416
rect 121380 83910 121408 91151
rect 122116 86902 122144 91287
rect 122746 91216 122802 91225
rect 122746 91151 122802 91160
rect 122104 86896 122156 86902
rect 122104 86838 122156 86844
rect 121368 83904 121420 83910
rect 121368 83846 121420 83852
rect 117228 81252 117280 81258
rect 117228 81194 117280 81200
rect 116584 79960 116636 79966
rect 116584 79902 116636 79908
rect 122760 79898 122788 91151
rect 122852 89418 122880 91423
rect 124034 91352 124090 91361
rect 124034 91287 124090 91296
rect 125414 91352 125470 91361
rect 125414 91287 125470 91296
rect 122840 89412 122892 89418
rect 122840 89354 122892 89360
rect 124048 88058 124076 91287
rect 124126 91216 124182 91225
rect 124126 91151 124182 91160
rect 124036 88052 124088 88058
rect 124036 87994 124088 88000
rect 124140 82754 124168 91151
rect 124128 82748 124180 82754
rect 124128 82690 124180 82696
rect 122748 79892 122800 79898
rect 122748 79834 122800 79840
rect 125428 78538 125456 91287
rect 125506 91216 125562 91225
rect 125506 91151 125562 91160
rect 125520 78606 125548 91151
rect 126532 90846 126560 92375
rect 126794 91216 126850 91225
rect 126794 91151 126850 91160
rect 126520 90840 126572 90846
rect 126520 90782 126572 90788
rect 126808 83978 126836 91151
rect 128188 91050 128216 93191
rect 165540 92478 165568 95882
rect 165528 92472 165580 92478
rect 130750 92440 130806 92449
rect 130750 92375 130752 92384
rect 130804 92375 130806 92384
rect 151542 92440 151598 92449
rect 151542 92375 151598 92384
rect 152922 92440 152978 92449
rect 165528 92414 165580 92420
rect 152922 92375 152978 92384
rect 130752 92346 130804 92352
rect 151556 92206 151584 92375
rect 151544 92200 151596 92206
rect 151544 92142 151596 92148
rect 151358 92032 151414 92041
rect 151358 91967 151414 91976
rect 132222 91624 132278 91633
rect 132222 91559 132278 91568
rect 129646 91216 129702 91225
rect 129646 91151 129702 91160
rect 129004 91112 129056 91118
rect 129004 91054 129056 91060
rect 128176 91044 128228 91050
rect 128176 90986 128228 90992
rect 126796 83972 126848 83978
rect 126796 83914 126848 83920
rect 125508 78600 125560 78606
rect 125508 78542 125560 78548
rect 125416 78532 125468 78538
rect 125416 78474 125468 78480
rect 129016 77110 129044 91054
rect 129660 81122 129688 91151
rect 132236 89350 132264 91559
rect 136454 91216 136510 91225
rect 136454 91151 136510 91160
rect 132224 89344 132276 89350
rect 132224 89286 132276 89292
rect 136468 88126 136496 91151
rect 151372 90710 151400 91967
rect 152936 90778 152964 92375
rect 166276 92138 166304 137974
rect 166448 125656 166500 125662
rect 166448 125598 166500 125604
rect 166356 124228 166408 124234
rect 166356 124170 166408 124176
rect 166264 92132 166316 92138
rect 166264 92074 166316 92080
rect 152924 90772 152976 90778
rect 152924 90714 152976 90720
rect 151360 90704 151412 90710
rect 151360 90646 151412 90652
rect 166368 89418 166396 124170
rect 166460 90846 166488 125598
rect 167552 111920 167604 111926
rect 167552 111862 167604 111868
rect 167564 110129 167592 111862
rect 167550 110120 167606 110129
rect 167550 110055 167606 110064
rect 166540 98048 166592 98054
rect 166540 97990 166592 97996
rect 166448 90840 166500 90846
rect 166448 90782 166500 90788
rect 166356 89412 166408 89418
rect 166356 89354 166408 89360
rect 136456 88120 136508 88126
rect 136456 88062 136508 88068
rect 166552 81326 166580 97990
rect 167656 93362 167684 146270
rect 171796 141438 171824 245006
rect 171888 235346 171916 258062
rect 171876 235340 171928 235346
rect 171876 235282 171928 235288
rect 171980 233034 172008 286350
rect 172072 276010 172100 294034
rect 173162 293992 173218 294001
rect 173162 293927 173218 293936
rect 172060 276004 172112 276010
rect 172060 275946 172112 275952
rect 172428 249824 172480 249830
rect 172428 249766 172480 249772
rect 171968 233028 172020 233034
rect 171968 232970 172020 232976
rect 171876 189236 171928 189242
rect 171876 189178 171928 189184
rect 171888 161430 171916 189178
rect 172440 183054 172468 249766
rect 172428 183048 172480 183054
rect 172428 182990 172480 182996
rect 171876 161424 171928 161430
rect 171876 161366 171928 161372
rect 171876 153264 171928 153270
rect 171876 153206 171928 153212
rect 171784 141432 171836 141438
rect 171784 141374 171836 141380
rect 170496 138100 170548 138106
rect 170496 138042 170548 138048
rect 167736 137284 167788 137290
rect 167736 137226 167788 137232
rect 167748 111926 167776 137226
rect 169024 135312 169076 135318
rect 169024 135254 169076 135260
rect 167828 118720 167880 118726
rect 167828 118662 167880 118668
rect 167736 111920 167788 111926
rect 167736 111862 167788 111868
rect 167736 111784 167788 111790
rect 167734 111752 167736 111761
rect 167788 111752 167790 111761
rect 167734 111687 167790 111696
rect 167736 108996 167788 109002
rect 167736 108938 167788 108944
rect 167748 108769 167776 108938
rect 167734 108760 167790 108769
rect 167734 108695 167790 108704
rect 167736 106344 167788 106350
rect 167736 106286 167788 106292
rect 167644 93356 167696 93362
rect 167644 93298 167696 93304
rect 166540 81320 166592 81326
rect 166540 81262 166592 81268
rect 129648 81116 129700 81122
rect 129648 81058 129700 81064
rect 167748 77178 167776 106286
rect 167840 90914 167868 118662
rect 167920 117360 167972 117366
rect 167920 117302 167972 117308
rect 167932 93226 167960 117302
rect 167920 93220 167972 93226
rect 167920 93162 167972 93168
rect 169036 90982 169064 135254
rect 170404 127016 170456 127022
rect 170404 126958 170456 126964
rect 169116 120148 169168 120154
rect 169116 120090 169168 120096
rect 169024 90976 169076 90982
rect 169024 90918 169076 90924
rect 167828 90908 167880 90914
rect 167828 90850 167880 90856
rect 169128 85202 169156 120090
rect 169208 110492 169260 110498
rect 169208 110434 169260 110440
rect 169116 85196 169168 85202
rect 169116 85138 169168 85144
rect 169220 84114 169248 110434
rect 169300 97300 169352 97306
rect 169300 97242 169352 97248
rect 169312 92313 169340 97242
rect 169298 92304 169354 92313
rect 169298 92239 169354 92248
rect 169208 84108 169260 84114
rect 169208 84050 169260 84056
rect 170416 79762 170444 126958
rect 170508 93294 170536 138042
rect 171784 129804 171836 129810
rect 171784 129746 171836 129752
rect 170588 109064 170640 109070
rect 170588 109006 170640 109012
rect 170496 93288 170548 93294
rect 170496 93230 170548 93236
rect 170600 85270 170628 109006
rect 170680 100020 170732 100026
rect 170680 99962 170732 99968
rect 170692 92274 170720 99962
rect 171796 93906 171824 129746
rect 171784 93900 171836 93906
rect 171784 93842 171836 93848
rect 171888 93430 171916 153206
rect 171968 144968 172020 144974
rect 171968 144910 172020 144916
rect 171876 93424 171928 93430
rect 171876 93366 171928 93372
rect 170680 92268 170732 92274
rect 170680 92210 170732 92216
rect 171980 89350 172008 144910
rect 172060 113212 172112 113218
rect 172060 113154 172112 113160
rect 171968 89344 172020 89350
rect 171968 89286 172020 89292
rect 170588 85264 170640 85270
rect 170588 85206 170640 85212
rect 172072 84046 172100 113154
rect 173176 92478 173204 293927
rect 173256 252612 173308 252618
rect 173256 252554 173308 252560
rect 173268 189854 173296 252554
rect 173348 248464 173400 248470
rect 173348 248406 173400 248412
rect 173360 236774 173388 248406
rect 173348 236768 173400 236774
rect 173348 236710 173400 236716
rect 173256 189848 173308 189854
rect 173256 189790 173308 189796
rect 173256 132524 173308 132530
rect 173256 132466 173308 132472
rect 173164 92472 173216 92478
rect 173164 92414 173216 92420
rect 172060 84040 172112 84046
rect 172060 83982 172112 83988
rect 173268 82550 173296 132466
rect 173348 118788 173400 118794
rect 173348 118730 173400 118736
rect 173360 94042 173388 118730
rect 173348 94036 173400 94042
rect 173348 93978 173400 93984
rect 173256 82544 173308 82550
rect 173256 82486 173308 82492
rect 170404 79756 170456 79762
rect 170404 79698 170456 79704
rect 167736 77172 167788 77178
rect 167736 77114 167788 77120
rect 129004 77104 129056 77110
rect 129004 77046 129056 77052
rect 111064 73092 111116 73098
rect 111064 73034 111116 73040
rect 106280 65612 106332 65618
rect 106280 65554 106332 65560
rect 106292 16574 106320 65554
rect 110420 64252 110472 64258
rect 110420 64194 110472 64200
rect 107660 42152 107712 42158
rect 107660 42094 107712 42100
rect 107672 16574 107700 42094
rect 102244 16546 103376 16574
rect 103532 16546 104112 16574
rect 106292 16546 106504 16574
rect 107672 16546 108160 16574
rect 102152 6886 102272 6914
rect 102244 480 102272 6886
rect 103348 480 103376 16546
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105728 15972 105780 15978
rect 105728 15914 105780 15920
rect 105740 480 105768 15914
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108132 480 108160 16546
rect 109040 13116 109092 13122
rect 109040 13058 109092 13064
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109052 354 109080 13058
rect 110432 6914 110460 64194
rect 114560 61464 114612 61470
rect 114560 61406 114612 61412
rect 113180 57384 113232 57390
rect 113180 57326 113232 57332
rect 110512 54596 110564 54602
rect 110512 54538 110564 54544
rect 110524 16574 110552 54538
rect 111800 32428 111852 32434
rect 111800 32370 111852 32376
rect 111812 16574 111840 32370
rect 113192 16574 113220 57326
rect 114572 16574 114600 61406
rect 117320 51876 117372 51882
rect 117320 51818 117372 51824
rect 110524 16546 111656 16574
rect 111812 16546 112392 16574
rect 113192 16546 114048 16574
rect 114572 16546 114784 16574
rect 110432 6886 110552 6914
rect 110524 480 110552 6886
rect 111628 480 111656 16546
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 114020 480 114048 16546
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116400 7676 116452 7682
rect 116400 7618 116452 7624
rect 116412 480 116440 7618
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 51818
rect 121460 50448 121512 50454
rect 121460 50390 121512 50396
rect 118700 49088 118752 49094
rect 118700 49030 118752 49036
rect 118712 16574 118740 49030
rect 120080 47660 120132 47666
rect 120080 47602 120132 47608
rect 120092 16574 120120 47602
rect 121472 16574 121500 50390
rect 124220 46300 124272 46306
rect 124220 46242 124272 46248
rect 124232 16574 124260 46242
rect 128360 17264 128412 17270
rect 128360 17206 128412 17212
rect 128372 16574 128400 17206
rect 118712 16546 118832 16574
rect 120092 16546 120672 16574
rect 121472 16546 122328 16574
rect 124232 16546 124720 16574
rect 128372 16546 128952 16574
rect 118804 480 118832 16546
rect 119896 3596 119948 3602
rect 119896 3538 119948 3544
rect 119908 480 119936 3538
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 122300 480 122328 16546
rect 123484 6248 123536 6254
rect 123484 6190 123536 6196
rect 123496 480 123524 6190
rect 124692 480 124720 16546
rect 125876 3664 125928 3670
rect 125876 3606 125928 3612
rect 125888 480 125916 3606
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 16546
rect 173820 13190 173848 321574
rect 174556 289814 174584 356322
rect 174648 344350 174676 357682
rect 174740 351218 174768 361694
rect 175924 354952 175976 354958
rect 175924 354894 175976 354900
rect 174728 351212 174780 351218
rect 174728 351154 174780 351160
rect 174636 344344 174688 344350
rect 174636 344286 174688 344292
rect 175188 342304 175240 342310
rect 175188 342246 175240 342252
rect 174544 289808 174596 289814
rect 174544 289750 174596 289756
rect 174544 282940 174596 282946
rect 174544 282882 174596 282888
rect 174556 238814 174584 282882
rect 174636 246356 174688 246362
rect 174636 246298 174688 246304
rect 174544 238808 174596 238814
rect 174544 238750 174596 238756
rect 174648 233986 174676 246298
rect 174636 233980 174688 233986
rect 174636 233922 174688 233928
rect 173898 175944 173954 175953
rect 173898 175879 173954 175888
rect 173808 13184 173860 13190
rect 173808 13126 173860 13132
rect 173912 3670 173940 175879
rect 174544 128376 174596 128382
rect 174544 128318 174596 128324
rect 174556 79830 174584 128318
rect 174636 112464 174688 112470
rect 174636 112406 174688 112412
rect 174648 92177 174676 112406
rect 174634 92168 174690 92177
rect 174634 92103 174690 92112
rect 174544 79824 174596 79830
rect 174544 79766 174596 79772
rect 175200 6322 175228 342246
rect 175936 292534 175964 354894
rect 176658 354376 176714 354385
rect 176658 354311 176714 354320
rect 176672 354006 176700 354311
rect 176660 354000 176712 354006
rect 176660 353942 176712 353948
rect 177856 353320 177908 353326
rect 177856 353262 177908 353268
rect 176566 352200 176622 352209
rect 176566 352135 176622 352144
rect 176474 336560 176530 336569
rect 176474 336495 176530 336504
rect 176014 292632 176070 292641
rect 176014 292567 176070 292576
rect 175924 292528 175976 292534
rect 175924 292470 175976 292476
rect 176028 238678 176056 292567
rect 176382 263800 176438 263809
rect 176382 263735 176438 263744
rect 176016 238672 176068 238678
rect 176016 238614 176068 238620
rect 176396 89078 176424 263735
rect 176384 89072 176436 89078
rect 176384 89014 176436 89020
rect 176488 27062 176516 336495
rect 176476 27056 176528 27062
rect 176476 26998 176528 27004
rect 176580 11898 176608 352135
rect 176658 348120 176714 348129
rect 176658 348055 176714 348064
rect 176672 347818 176700 348055
rect 176660 347812 176712 347818
rect 176660 347754 176712 347760
rect 176658 343360 176714 343369
rect 176658 343295 176714 343304
rect 176672 342310 176700 343295
rect 176660 342304 176712 342310
rect 176660 342246 176712 342252
rect 176658 341320 176714 341329
rect 176658 341255 176714 341264
rect 176672 340950 176700 341255
rect 176660 340944 176712 340950
rect 176660 340886 176712 340892
rect 176660 332648 176712 332654
rect 176658 332616 176660 332625
rect 176712 332616 176714 332625
rect 176658 332551 176714 332560
rect 176660 321632 176712 321638
rect 176658 321600 176660 321609
rect 176712 321600 176714 321609
rect 176658 321535 176714 321544
rect 177762 318880 177818 318889
rect 177762 318815 177818 318824
rect 176658 314800 176714 314809
rect 176658 314735 176714 314744
rect 176672 314702 176700 314735
rect 176660 314696 176712 314702
rect 176660 314638 176712 314644
rect 176658 310040 176714 310049
rect 176658 309975 176714 309984
rect 176672 309194 176700 309975
rect 176660 309188 176712 309194
rect 176660 309130 176712 309136
rect 176658 308000 176714 308009
rect 176658 307935 176714 307944
rect 176672 307902 176700 307935
rect 176660 307896 176712 307902
rect 176660 307838 176712 307844
rect 176658 305960 176714 305969
rect 176658 305895 176714 305904
rect 176672 305046 176700 305895
rect 176660 305040 176712 305046
rect 176660 304982 176712 304988
rect 177670 301200 177726 301209
rect 177670 301135 177726 301144
rect 176660 299464 176712 299470
rect 176660 299406 176712 299412
rect 176672 299305 176700 299406
rect 176658 299296 176714 299305
rect 176658 299231 176714 299240
rect 176660 298104 176712 298110
rect 176660 298046 176712 298052
rect 176672 297265 176700 298046
rect 176658 297256 176714 297265
rect 176658 297191 176714 297200
rect 176658 295080 176714 295089
rect 176658 295015 176714 295024
rect 176672 294030 176700 295015
rect 176660 294024 176712 294030
rect 176660 293966 176712 293972
rect 176658 292360 176714 292369
rect 176658 292295 176714 292304
rect 176672 291242 176700 292295
rect 176660 291236 176712 291242
rect 176660 291178 176712 291184
rect 176658 290320 176714 290329
rect 176658 290255 176714 290264
rect 176672 289882 176700 290255
rect 176660 289876 176712 289882
rect 176660 289818 176712 289824
rect 176660 282872 176712 282878
rect 176660 282814 176712 282820
rect 176672 281625 176700 282814
rect 176658 281616 176714 281625
rect 176658 281551 176714 281560
rect 176752 280152 176804 280158
rect 176752 280094 176804 280100
rect 176764 279585 176792 280094
rect 176750 279576 176806 279585
rect 176750 279511 176806 279520
rect 176658 277536 176714 277545
rect 176658 277471 176714 277480
rect 176672 277438 176700 277471
rect 176660 277432 176712 277438
rect 176660 277374 176712 277380
rect 176660 276004 176712 276010
rect 176660 275946 176712 275952
rect 176672 274825 176700 275946
rect 176658 274816 176714 274825
rect 176658 274751 176714 274760
rect 176660 273216 176712 273222
rect 176660 273158 176712 273164
rect 176672 272785 176700 273158
rect 176658 272776 176714 272785
rect 176658 272711 176714 272720
rect 176658 268560 176714 268569
rect 176658 268495 176714 268504
rect 176672 267850 176700 268495
rect 176660 267844 176712 267850
rect 176660 267786 176712 267792
rect 176660 266348 176712 266354
rect 176660 266290 176712 266296
rect 176672 265985 176700 266290
rect 176658 265976 176714 265985
rect 176658 265911 176714 265920
rect 176660 262132 176712 262138
rect 176660 262074 176712 262080
rect 176672 261905 176700 262074
rect 176658 261896 176714 261905
rect 176658 261831 176714 261840
rect 176658 259720 176714 259729
rect 176658 259655 176714 259664
rect 176672 259554 176700 259655
rect 176660 259548 176712 259554
rect 176660 259490 176712 259496
rect 176842 254960 176898 254969
rect 176842 254895 176898 254904
rect 176856 254153 176884 254895
rect 176842 254144 176898 254153
rect 176842 254079 176898 254088
rect 176658 250880 176714 250889
rect 176658 250815 176714 250824
rect 176672 249830 176700 250815
rect 176660 249824 176712 249830
rect 176660 249766 176712 249772
rect 176844 242752 176896 242758
rect 176844 242694 176896 242700
rect 176856 242185 176884 242694
rect 176842 242176 176898 242185
rect 176842 242111 176898 242120
rect 177684 151094 177712 301135
rect 177672 151088 177724 151094
rect 177672 151030 177724 151036
rect 177776 140078 177804 318815
rect 177868 286385 177896 353262
rect 177960 334665 177988 702510
rect 193220 700392 193272 700398
rect 193220 700334 193272 700340
rect 189724 683188 189776 683194
rect 189724 683130 189776 683136
rect 179328 630692 179380 630698
rect 179328 630634 179380 630640
rect 179052 374672 179104 374678
rect 179052 374614 179104 374620
rect 177946 334656 178002 334665
rect 177946 334591 177948 334600
rect 178000 334591 178002 334600
rect 177948 334562 178000 334568
rect 177960 334531 177988 334562
rect 179064 316034 179092 374614
rect 179144 370524 179196 370530
rect 179144 370466 179196 370472
rect 178972 316006 179092 316034
rect 178972 312769 179000 316006
rect 178958 312760 179014 312769
rect 178958 312695 179014 312704
rect 178972 311914 179000 312695
rect 178960 311908 179012 311914
rect 178960 311850 179012 311856
rect 177946 303920 178002 303929
rect 177946 303855 178002 303864
rect 177854 286376 177910 286385
rect 177854 286311 177856 286320
rect 177908 286311 177910 286320
rect 177856 286282 177908 286288
rect 177868 286251 177896 286282
rect 177854 270600 177910 270609
rect 177854 270535 177910 270544
rect 177764 140072 177816 140078
rect 177764 140014 177816 140020
rect 177304 136672 177356 136678
rect 177304 136614 177356 136620
rect 177316 93974 177344 136614
rect 177396 111852 177448 111858
rect 177396 111794 177448 111800
rect 177304 93968 177356 93974
rect 177304 93910 177356 93916
rect 177408 89486 177436 111794
rect 177396 89480 177448 89486
rect 177396 89422 177448 89428
rect 177868 80782 177896 270535
rect 177856 80776 177908 80782
rect 177856 80718 177908 80724
rect 177960 65686 177988 303855
rect 179050 279576 179106 279585
rect 179050 279511 179106 279520
rect 178684 264988 178736 264994
rect 178684 264930 178736 264936
rect 178696 95198 178724 264930
rect 179064 220114 179092 279511
rect 179156 245993 179184 370466
rect 179236 362976 179288 362982
rect 179236 362918 179288 362924
rect 179248 288289 179276 362918
rect 179234 288280 179290 288289
rect 179234 288215 179290 288224
rect 179340 254969 179368 630634
rect 179420 377460 179472 377466
rect 179420 377402 179472 377408
rect 179432 257009 179460 377402
rect 189736 371890 189764 683130
rect 189724 371884 189776 371890
rect 189724 371826 189776 371832
rect 190460 364540 190512 364546
rect 190460 364482 190512 364488
rect 179880 364404 179932 364410
rect 179880 364346 179932 364352
rect 179788 357672 179840 357678
rect 179788 357614 179840 357620
rect 179602 355056 179658 355065
rect 179602 354991 179658 355000
rect 179616 352578 179644 354991
rect 179800 354074 179828 357614
rect 179788 354068 179840 354074
rect 179788 354010 179840 354016
rect 179892 353326 179920 364346
rect 190472 364334 190500 364482
rect 190472 364306 191236 364334
rect 189998 363080 190054 363089
rect 189998 363015 190054 363024
rect 184940 359032 184992 359038
rect 184940 358974 184992 358980
rect 181628 358896 181680 358902
rect 181628 358838 181680 358844
rect 181640 355042 181668 358838
rect 182914 357776 182970 357785
rect 182914 357711 182970 357720
rect 181332 355014 181668 355042
rect 182928 355042 182956 357711
rect 184952 355042 184980 358974
rect 187424 358080 187476 358086
rect 187424 358022 187476 358028
rect 187436 355042 187464 358022
rect 190012 355042 190040 363015
rect 182928 355014 183264 355042
rect 184952 355014 185196 355042
rect 187128 355014 187464 355042
rect 189704 355014 190040 355042
rect 191208 355042 191236 364306
rect 193232 357610 193260 700334
rect 195888 376032 195940 376038
rect 195888 375974 195940 375980
rect 195900 368966 195928 375974
rect 201512 373318 201540 702986
rect 209780 702636 209832 702642
rect 209780 702578 209832 702584
rect 206284 702500 206336 702506
rect 206284 702442 206336 702448
rect 202880 474768 202932 474774
rect 202880 474710 202932 474716
rect 201500 373312 201552 373318
rect 201500 373254 201552 373260
rect 198740 371884 198792 371890
rect 198740 371826 198792 371832
rect 194600 368960 194652 368966
rect 194600 368902 194652 368908
rect 195888 368960 195940 368966
rect 195888 368902 195940 368908
rect 194612 368626 194640 368902
rect 194600 368620 194652 368626
rect 194600 368562 194652 368568
rect 194612 364334 194640 368562
rect 194612 364306 195100 364334
rect 193220 357604 193272 357610
rect 193220 357546 193272 357552
rect 193232 355042 193260 357546
rect 195072 355042 195100 364306
rect 197728 360528 197780 360534
rect 197728 360470 197780 360476
rect 197740 355042 197768 360470
rect 198752 355094 198780 371826
rect 201592 360460 201644 360466
rect 201592 360402 201644 360408
rect 198740 355088 198792 355094
rect 191208 355014 191636 355042
rect 193232 355014 193568 355042
rect 195072 355014 195500 355042
rect 197740 355014 198076 355042
rect 198740 355030 198792 355036
rect 199660 355088 199712 355094
rect 201604 355042 201632 360402
rect 202892 355298 202920 474710
rect 206296 356153 206324 702442
rect 206376 371272 206428 371278
rect 206376 371214 206428 371220
rect 206388 358086 206416 371214
rect 209044 369164 209096 369170
rect 209044 369106 209096 369112
rect 209056 364334 209084 369106
rect 208780 364306 209084 364334
rect 209792 364334 209820 702578
rect 218992 700330 219020 703520
rect 235184 700398 235212 703520
rect 235172 700392 235224 700398
rect 235172 700334 235224 700340
rect 218980 700324 219032 700330
rect 218980 700266 219032 700272
rect 267660 697678 267688 703520
rect 283852 702434 283880 703520
rect 282932 702406 283880 702434
rect 266360 697672 266412 697678
rect 266360 697614 266412 697620
rect 267648 697672 267700 697678
rect 267648 697614 267700 697620
rect 211804 697604 211856 697610
rect 211804 697546 211856 697552
rect 209792 364306 209912 364334
rect 206376 358080 206428 358086
rect 206376 358022 206428 358028
rect 208780 356386 208808 364306
rect 208768 356380 208820 356386
rect 208768 356322 208820 356328
rect 206282 356144 206338 356153
rect 206282 356079 206338 356088
rect 202880 355292 202932 355298
rect 202880 355234 202932 355240
rect 203846 355292 203898 355298
rect 203846 355234 203898 355240
rect 199712 355036 200008 355042
rect 199660 355030 200008 355036
rect 199672 355014 200008 355030
rect 201604 355014 201940 355042
rect 202892 355026 202920 355234
rect 203858 355028 203886 355234
rect 206296 355042 206324 356079
rect 208780 355042 208808 356322
rect 202880 355020 202932 355026
rect 206296 355014 206448 355042
rect 208380 355014 208808 355042
rect 209884 355042 209912 364306
rect 211816 357678 211844 697546
rect 220084 378208 220136 378214
rect 220084 378150 220136 378156
rect 220096 369170 220124 378150
rect 266372 377466 266400 697614
rect 278044 470620 278096 470626
rect 278044 470562 278096 470568
rect 266360 377460 266412 377466
rect 266360 377402 266412 377408
rect 220084 369164 220136 369170
rect 220084 369106 220136 369112
rect 254584 367124 254636 367130
rect 254584 367066 254636 367072
rect 242900 364472 242952 364478
rect 242900 364414 242952 364420
rect 242912 364334 242940 364414
rect 242912 364306 243400 364334
rect 214472 363112 214524 363118
rect 214472 363054 214524 363060
rect 211804 357672 211856 357678
rect 211804 357614 211856 357620
rect 211816 355042 211844 357614
rect 214484 355042 214512 363054
rect 237472 361752 237524 361758
rect 233790 361720 233846 361729
rect 237472 361694 237524 361700
rect 233790 361655 233846 361664
rect 225420 360460 225472 360466
rect 225420 360402 225472 360408
rect 220268 360256 220320 360262
rect 220268 360198 220320 360204
rect 218334 357640 218390 357649
rect 217048 357604 217100 357610
rect 218334 357575 218390 357584
rect 217048 357546 217100 357552
rect 217060 355042 217088 357546
rect 209884 355014 210312 355042
rect 211816 355014 212244 355042
rect 214484 355014 214820 355042
rect 216752 355014 217088 355042
rect 218348 355042 218376 357575
rect 220280 355042 220308 360198
rect 223488 357672 223540 357678
rect 223488 357614 223540 357620
rect 223500 355042 223528 357614
rect 225432 355042 225460 360402
rect 231214 357912 231270 357921
rect 231214 357847 231270 357856
rect 227350 357504 227406 357513
rect 227350 357439 227406 357448
rect 227364 355042 227392 357439
rect 228822 356144 228878 356153
rect 228822 356079 228878 356088
rect 218348 355014 218684 355042
rect 220280 355014 220616 355042
rect 223192 355014 223528 355042
rect 225124 355014 225460 355042
rect 227056 355014 227392 355042
rect 202880 354962 202932 354968
rect 209884 354929 209912 355014
rect 209870 354920 209926 354929
rect 209870 354855 209926 354864
rect 228836 354770 228864 356079
rect 231228 355042 231256 357847
rect 233804 355042 233832 361655
rect 231228 355014 231564 355042
rect 233496 355014 233832 355042
rect 235080 354952 235132 354958
rect 237484 354906 237512 361694
rect 242808 357808 242860 357814
rect 242808 357750 242860 357756
rect 241520 357740 241572 357746
rect 241520 357682 241572 357688
rect 240046 356280 240102 356289
rect 240046 356215 240102 356224
rect 240060 355042 240088 356215
rect 239936 355014 240088 355042
rect 241532 355042 241560 357682
rect 242820 357406 242848 357750
rect 242808 357400 242860 357406
rect 242808 357342 242860 357348
rect 243372 355042 243400 364306
rect 245844 361616 245896 361622
rect 245844 361558 245896 361564
rect 241532 355014 241868 355042
rect 243372 355014 243800 355042
rect 235132 354900 235428 354906
rect 235080 354894 235428 354900
rect 235092 354878 235428 354894
rect 237360 354878 237512 354906
rect 245856 354770 245884 361558
rect 254596 360262 254624 367066
rect 276020 365832 276072 365838
rect 276020 365774 276072 365780
rect 276032 364334 276060 365774
rect 276032 364306 276888 364334
rect 273536 361752 273588 361758
rect 273536 361694 273588 361700
rect 256792 361684 256844 361690
rect 256792 361626 256844 361632
rect 254400 360256 254452 360262
rect 254400 360198 254452 360204
rect 254584 360256 254636 360262
rect 254584 360198 254636 360204
rect 250534 357640 250590 357649
rect 250534 357575 250590 357584
rect 247960 356244 248012 356250
rect 247960 356186 248012 356192
rect 247972 355042 248000 356186
rect 250548 355042 250576 357575
rect 252468 356244 252520 356250
rect 252468 356186 252520 356192
rect 252480 355042 252508 356186
rect 254412 355042 254440 360198
rect 247972 355014 248308 355042
rect 250240 355014 250576 355042
rect 252172 355014 252508 355042
rect 254104 355014 254440 355042
rect 256804 354958 256832 361626
rect 269028 357876 269080 357882
rect 269028 357818 269080 357824
rect 260748 357740 260800 357746
rect 260748 357682 260800 357688
rect 258908 356380 258960 356386
rect 258908 356322 258960 356328
rect 258920 355042 258948 356322
rect 260760 355042 260788 357682
rect 265164 357468 265216 357474
rect 265164 357410 265216 357416
rect 258612 355014 258948 355042
rect 260544 355014 260788 355042
rect 256792 354952 256844 354958
rect 256680 354900 256792 354906
rect 256680 354894 256844 354900
rect 256680 354878 256832 354894
rect 256804 354829 256832 354878
rect 228836 354742 228988 354770
rect 245732 354742 245884 354770
rect 262218 354784 262274 354793
rect 265176 354770 265204 357410
rect 269040 355042 269068 357818
rect 270500 357808 270552 357814
rect 270500 357750 270552 357756
rect 268916 355014 269068 355042
rect 270512 355042 270540 357750
rect 273548 356318 273576 361694
rect 273536 356312 273588 356318
rect 273536 356254 273588 356260
rect 270512 355014 270848 355042
rect 273548 354906 273576 356254
rect 276860 355042 276888 364306
rect 278056 361758 278084 470562
rect 282932 362234 282960 702406
rect 300136 699718 300164 703520
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 301504 702704 301556 702710
rect 301504 702646 301556 702652
rect 300124 699712 300176 699718
rect 300124 699654 300176 699660
rect 297364 683188 297416 683194
rect 297364 683130 297416 683136
rect 295616 368552 295668 368558
rect 295616 368494 295668 368500
rect 287060 365764 287112 365770
rect 287060 365706 287112 365712
rect 287072 364334 287100 365706
rect 287072 364306 287192 364334
rect 282920 362228 282972 362234
rect 282920 362170 282972 362176
rect 278044 361752 278096 361758
rect 278044 361694 278096 361700
rect 279332 360392 279384 360398
rect 279332 360334 279384 360340
rect 275356 355026 275692 355042
rect 275356 355020 275704 355026
rect 275356 355014 275652 355020
rect 276860 355014 277288 355042
rect 275652 354962 275704 354968
rect 273424 354878 273576 354906
rect 279344 354770 279372 360334
rect 283380 359100 283432 359106
rect 283380 359042 283432 359048
rect 282092 358964 282144 358970
rect 282092 358906 282144 358912
rect 282104 355042 282132 358906
rect 281796 355014 282132 355042
rect 283392 355042 283420 359042
rect 287164 357474 287192 364306
rect 295340 363044 295392 363050
rect 295340 362986 295392 362992
rect 291844 360324 291896 360330
rect 291844 360266 291896 360272
rect 291752 357672 291804 357678
rect 291752 357614 291804 357620
rect 289452 357536 289504 357542
rect 289452 357478 289504 357484
rect 290464 357536 290516 357542
rect 290464 357478 290516 357484
rect 287152 357468 287204 357474
rect 287152 357410 287204 357416
rect 285956 356312 286008 356318
rect 285956 356254 286008 356260
rect 285968 355042 285996 356254
rect 283392 355014 283728 355042
rect 285660 355014 285996 355042
rect 287164 355042 287192 357410
rect 289464 356046 289492 357478
rect 289452 356040 289504 356046
rect 289452 355982 289504 355988
rect 290476 355042 290504 357478
rect 287164 355014 287592 355042
rect 290168 355014 290504 355042
rect 262274 354742 262476 354770
rect 265052 354742 265204 354770
rect 266648 354754 266984 354770
rect 266636 354748 266984 354754
rect 262218 354719 262274 354728
rect 266688 354742 266984 354748
rect 279220 354754 279556 354770
rect 279220 354748 279568 354754
rect 279220 354742 279516 354748
rect 266636 354690 266688 354696
rect 279516 354690 279568 354696
rect 291764 354657 291792 357614
rect 291856 355042 291884 360266
rect 294144 358828 294196 358834
rect 294144 358770 294196 358776
rect 293316 357468 293368 357474
rect 293316 357410 293368 357416
rect 291856 355014 293172 355042
rect 293040 354884 293092 354890
rect 293040 354826 293092 354832
rect 291750 354648 291806 354657
rect 291750 354583 291806 354592
rect 179880 353320 179932 353326
rect 179880 353262 179932 353268
rect 179604 352572 179656 352578
rect 179604 352514 179656 352520
rect 179510 351928 179566 351937
rect 179510 351863 179566 351872
rect 179524 325757 179552 351863
rect 293052 330449 293080 354826
rect 293144 351218 293172 355014
rect 293328 354006 293356 357410
rect 294052 354816 294104 354822
rect 294052 354758 294104 354764
rect 293316 354000 293368 354006
rect 293316 353942 293368 353948
rect 293958 352336 294014 352345
rect 293958 352271 294014 352280
rect 293132 351212 293184 351218
rect 293132 351154 293184 351160
rect 293038 330440 293094 330449
rect 293038 330375 293094 330384
rect 179510 325748 179566 325757
rect 179510 325683 179512 325692
rect 179564 325683 179566 325692
rect 179512 325654 179564 325660
rect 179510 316908 179566 316917
rect 179510 316843 179566 316852
rect 179418 257000 179474 257009
rect 179418 256935 179474 256944
rect 179326 254960 179382 254969
rect 179326 254895 179382 254904
rect 179418 252920 179474 252929
rect 179418 252855 179474 252864
rect 179234 248160 179290 248169
rect 179234 248095 179290 248104
rect 179142 245984 179198 245993
rect 179142 245919 179198 245928
rect 179052 220108 179104 220114
rect 179052 220050 179104 220056
rect 178776 121508 178828 121514
rect 178776 121450 178828 121456
rect 178684 95192 178736 95198
rect 178684 95134 178736 95140
rect 178788 93158 178816 121450
rect 178776 93152 178828 93158
rect 178776 93094 178828 93100
rect 177948 65680 178000 65686
rect 177948 65622 178000 65628
rect 179248 51814 179276 248095
rect 179326 244080 179382 244089
rect 179326 244015 179382 244024
rect 179236 51808 179288 51814
rect 179236 51750 179288 51756
rect 176568 11892 176620 11898
rect 176568 11834 176620 11840
rect 175188 6316 175240 6322
rect 175188 6258 175240 6264
rect 173900 3664 173952 3670
rect 173900 3606 173952 3612
rect 179340 2174 179368 244015
rect 179432 10402 179460 252855
rect 179524 243001 179552 316843
rect 293130 301336 293186 301345
rect 293130 301271 293186 301280
rect 293038 287464 293094 287473
rect 293038 287399 293094 287408
rect 179510 242992 179566 243001
rect 179510 242927 179566 242936
rect 179696 242956 179748 242962
rect 179696 242898 179748 242904
rect 179708 240378 179736 242898
rect 188342 240680 188398 240689
rect 182824 240644 182876 240650
rect 188342 240615 188398 240624
rect 182824 240586 182876 240592
rect 179696 240372 179748 240378
rect 179696 240314 179748 240320
rect 179800 240230 180044 240258
rect 179800 240122 179828 240230
rect 179524 240094 179828 240122
rect 179880 240168 179932 240174
rect 179880 240110 179932 240116
rect 179524 28422 179552 240094
rect 179892 231742 179920 240110
rect 180812 240094 181976 240122
rect 179880 231736 179932 231742
rect 179880 231678 179932 231684
rect 180064 124296 180116 124302
rect 180064 124238 180116 124244
rect 180076 88058 180104 124238
rect 180064 88052 180116 88058
rect 180064 87994 180116 88000
rect 180812 33998 180840 240094
rect 182836 225758 182864 240586
rect 183572 240094 183908 240122
rect 184952 240094 185840 240122
rect 182824 225752 182876 225758
rect 182824 225694 182876 225700
rect 182824 146396 182876 146402
rect 182824 146338 182876 146344
rect 181444 113280 181496 113286
rect 181444 113222 181496 113228
rect 181456 85338 181484 113222
rect 182836 94110 182864 146338
rect 183008 130416 183060 130422
rect 183008 130358 183060 130364
rect 182916 114572 182968 114578
rect 182916 114514 182968 114520
rect 182824 94104 182876 94110
rect 182824 94046 182876 94052
rect 181444 85332 181496 85338
rect 181444 85274 181496 85280
rect 182928 75818 182956 114514
rect 183020 92342 183048 130358
rect 183008 92336 183060 92342
rect 183008 92278 183060 92284
rect 182916 75812 182968 75818
rect 182916 75754 182968 75760
rect 180800 33992 180852 33998
rect 180800 33934 180852 33940
rect 179512 28416 179564 28422
rect 179512 28358 179564 28364
rect 183572 21554 183600 240094
rect 184204 153332 184256 153338
rect 184204 153274 184256 153280
rect 184216 90710 184244 153274
rect 184204 90704 184256 90710
rect 184204 90646 184256 90652
rect 184952 76634 184980 240094
rect 187758 239850 187786 240108
rect 187712 239822 187786 239850
rect 186964 234048 187016 234054
rect 186964 233990 187016 233996
rect 186976 175953 187004 233990
rect 187056 176792 187108 176798
rect 187056 176734 187108 176740
rect 186962 175944 187018 175953
rect 186962 175879 187018 175888
rect 187068 149054 187096 176734
rect 187056 149048 187108 149054
rect 187056 148990 187108 148996
rect 185584 122868 185636 122874
rect 185584 122810 185636 122816
rect 185596 83910 185624 122810
rect 186964 121576 187016 121582
rect 186964 121518 187016 121524
rect 185676 114640 185728 114646
rect 185676 114582 185728 114588
rect 185688 85406 185716 114582
rect 186976 86766 187004 121518
rect 187056 116000 187108 116006
rect 187056 115942 187108 115948
rect 187068 86834 187096 115942
rect 187056 86828 187108 86834
rect 187056 86770 187108 86776
rect 186964 86760 187016 86766
rect 186964 86702 187016 86708
rect 185676 85400 185728 85406
rect 185676 85342 185728 85348
rect 185584 83904 185636 83910
rect 185584 83846 185636 83852
rect 184940 76628 184992 76634
rect 184940 76570 184992 76576
rect 187712 24342 187740 239822
rect 188356 237182 188384 240615
rect 279864 240366 280016 240394
rect 190012 240094 190348 240122
rect 191944 240094 192280 240122
rect 193232 240094 194212 240122
rect 195992 240094 196144 240122
rect 190012 239057 190040 240094
rect 189998 239048 190054 239057
rect 189998 238983 190054 238992
rect 190012 238746 190040 238983
rect 190000 238740 190052 238746
rect 190000 238682 190052 238688
rect 189724 238060 189776 238066
rect 189724 238002 189776 238008
rect 188344 237176 188396 237182
rect 188344 237118 188396 237124
rect 189736 205154 189764 238002
rect 191944 237250 191972 240094
rect 191932 237244 191984 237250
rect 191932 237186 191984 237192
rect 192484 236768 192536 236774
rect 192484 236710 192536 236716
rect 189908 205216 189960 205222
rect 189908 205158 189960 205164
rect 189724 205148 189776 205154
rect 189724 205090 189776 205096
rect 189816 189168 189868 189174
rect 189816 189110 189868 189116
rect 189724 187332 189776 187338
rect 189724 187274 189776 187280
rect 188344 143608 188396 143614
rect 188344 143550 188396 143556
rect 188356 91050 188384 143550
rect 188436 127084 188488 127090
rect 188436 127026 188488 127032
rect 188344 91044 188396 91050
rect 188344 90986 188396 90992
rect 188448 78674 188476 127026
rect 188436 78668 188488 78674
rect 188436 78610 188488 78616
rect 189736 32502 189764 187274
rect 189828 166938 189856 189110
rect 189920 182986 189948 205158
rect 192496 196926 192524 236710
rect 192484 196920 192536 196926
rect 192484 196862 192536 196868
rect 192482 184376 192538 184385
rect 192482 184311 192538 184320
rect 189908 182980 189960 182986
rect 189908 182922 189960 182928
rect 189816 166932 189868 166938
rect 189816 166874 189868 166880
rect 191104 151836 191156 151842
rect 191104 151778 191156 151784
rect 189816 133952 189868 133958
rect 189816 133894 189868 133900
rect 189828 82686 189856 133894
rect 189908 116068 189960 116074
rect 189908 116010 189960 116016
rect 189920 89554 189948 116010
rect 191116 90778 191144 151778
rect 191196 102196 191248 102202
rect 191196 102138 191248 102144
rect 191104 90772 191156 90778
rect 191104 90714 191156 90720
rect 189908 89548 189960 89554
rect 189908 89490 189960 89496
rect 189816 82680 189868 82686
rect 189816 82622 189868 82628
rect 191208 75886 191236 102138
rect 191196 75880 191248 75886
rect 191196 75822 191248 75828
rect 189724 32496 189776 32502
rect 189724 32438 189776 32444
rect 187700 24336 187752 24342
rect 187700 24278 187752 24284
rect 183560 21548 183612 21554
rect 183560 21490 183612 21496
rect 192496 16046 192524 184311
rect 192576 118856 192628 118862
rect 192576 118798 192628 118804
rect 192588 82618 192616 118798
rect 192668 110560 192720 110566
rect 192668 110502 192720 110508
rect 192680 88194 192708 110502
rect 192668 88188 192720 88194
rect 192668 88130 192720 88136
rect 192576 82612 192628 82618
rect 192576 82554 192628 82560
rect 193232 17338 193260 240094
rect 195992 238542 196020 240094
rect 198706 239850 198734 240108
rect 200132 240094 200652 240122
rect 201512 240094 202584 240122
rect 204516 240094 204944 240122
rect 198706 239822 198780 239850
rect 195980 238536 196032 238542
rect 195980 238478 196032 238484
rect 198004 235408 198056 235414
rect 198004 235350 198056 235356
rect 196716 233912 196768 233918
rect 196716 233854 196768 233860
rect 196728 194206 196756 233854
rect 198016 207942 198044 235350
rect 198004 207936 198056 207942
rect 198004 207878 198056 207884
rect 198002 196616 198058 196625
rect 198002 196551 198058 196560
rect 196716 194200 196768 194206
rect 196716 194142 196768 194148
rect 196622 193896 196678 193905
rect 196622 193831 196678 193840
rect 195980 176724 196032 176730
rect 195980 176666 196032 176672
rect 195992 175234 196020 176666
rect 195980 175228 196032 175234
rect 195980 175170 196032 175176
rect 193956 145036 194008 145042
rect 193956 144978 194008 144984
rect 193864 135380 193916 135386
rect 193864 135322 193916 135328
rect 193876 81190 193904 135322
rect 193968 92410 193996 144978
rect 195244 142180 195296 142186
rect 195244 142122 195296 142128
rect 194048 104916 194100 104922
rect 194048 104858 194100 104864
rect 193956 92404 194008 92410
rect 193956 92346 194008 92352
rect 193864 81184 193916 81190
rect 193864 81126 193916 81132
rect 194060 74526 194088 104858
rect 195256 83978 195284 142122
rect 195244 83972 195296 83978
rect 195244 83914 195296 83920
rect 194048 74520 194100 74526
rect 194048 74462 194100 74468
rect 193220 17332 193272 17338
rect 193220 17274 193272 17280
rect 192484 16040 192536 16046
rect 192484 15982 192536 15988
rect 179420 10396 179472 10402
rect 179420 10338 179472 10344
rect 196636 3670 196664 193831
rect 196716 178152 196768 178158
rect 196716 178094 196768 178100
rect 196728 168298 196756 178094
rect 196716 168292 196768 168298
rect 196716 168234 196768 168240
rect 196808 145580 196860 145586
rect 196808 145522 196860 145528
rect 196716 120216 196768 120222
rect 196716 120158 196768 120164
rect 196728 81258 196756 120158
rect 196820 109002 196848 145522
rect 196808 108996 196860 109002
rect 196808 108938 196860 108944
rect 196900 104984 196952 104990
rect 196900 104926 196952 104932
rect 196808 98116 196860 98122
rect 196808 98058 196860 98064
rect 196716 81252 196768 81258
rect 196716 81194 196768 81200
rect 196820 77110 196848 98058
rect 196912 94897 196940 104926
rect 196898 94888 196954 94897
rect 196898 94823 196954 94832
rect 196808 77104 196860 77110
rect 196808 77046 196860 77052
rect 198016 9110 198044 196551
rect 198096 147688 198148 147694
rect 198096 147630 198148 147636
rect 198108 88126 198136 147630
rect 198188 99408 198240 99414
rect 198188 99350 198240 99356
rect 198096 88120 198148 88126
rect 198096 88062 198148 88068
rect 198200 73098 198228 99350
rect 198752 80714 198780 239822
rect 199384 107704 199436 107710
rect 199384 107646 199436 107652
rect 199396 81394 199424 107646
rect 199476 103556 199528 103562
rect 199476 103498 199528 103504
rect 199488 95062 199516 103498
rect 199476 95056 199528 95062
rect 199476 94998 199528 95004
rect 199384 81388 199436 81394
rect 199384 81330 199436 81336
rect 198740 80708 198792 80714
rect 198740 80650 198792 80656
rect 198188 73092 198240 73098
rect 198188 73034 198240 73040
rect 200132 29782 200160 240094
rect 201512 33930 201540 240094
rect 204916 238513 204944 240094
rect 207078 239850 207106 240108
rect 207032 239822 207106 239850
rect 208412 240094 209024 240122
rect 210620 240094 210956 240122
rect 212552 240094 212888 240122
rect 215312 240094 215464 240122
rect 217060 240094 217396 240122
rect 218992 240094 219328 240122
rect 220832 240094 221260 240122
rect 204902 238504 204958 238513
rect 204902 238439 204958 238448
rect 203616 190528 203668 190534
rect 203616 190470 203668 190476
rect 203524 180328 203576 180334
rect 203524 180270 203576 180276
rect 202144 177540 202196 177546
rect 202144 177482 202196 177488
rect 201500 33924 201552 33930
rect 201500 33866 201552 33872
rect 200120 29776 200172 29782
rect 200120 29718 200172 29724
rect 198004 9104 198056 9110
rect 198004 9046 198056 9052
rect 202156 3738 202184 177482
rect 202236 131164 202288 131170
rect 202236 131106 202288 131112
rect 202248 85542 202276 131106
rect 202328 103624 202380 103630
rect 202328 103566 202380 103572
rect 202340 90953 202368 103566
rect 202326 90944 202382 90953
rect 202326 90879 202382 90888
rect 202236 85536 202288 85542
rect 202236 85478 202288 85484
rect 203536 6390 203564 180270
rect 203628 158710 203656 190470
rect 203616 158704 203668 158710
rect 203616 158646 203668 158652
rect 203616 151904 203668 151910
rect 203616 151846 203668 151852
rect 203628 92206 203656 151846
rect 203708 117428 203760 117434
rect 203708 117370 203760 117376
rect 203616 92200 203668 92206
rect 203616 92142 203668 92148
rect 203720 88262 203748 117370
rect 204916 89010 204944 238439
rect 206284 228540 206336 228546
rect 206284 228482 206336 228488
rect 206296 188630 206324 228482
rect 206284 188624 206336 188630
rect 206284 188566 206336 188572
rect 206468 182232 206520 182238
rect 206468 182174 206520 182180
rect 206284 178220 206336 178226
rect 206284 178162 206336 178168
rect 206296 150414 206324 178162
rect 206376 176248 206428 176254
rect 206376 176190 206428 176196
rect 206388 162790 206416 176190
rect 206480 171018 206508 182174
rect 206560 180872 206612 180878
rect 206560 180814 206612 180820
rect 206572 172514 206600 180814
rect 206560 172508 206612 172514
rect 206560 172450 206612 172456
rect 206468 171012 206520 171018
rect 206468 170954 206520 170960
rect 206376 162784 206428 162790
rect 206376 162726 206428 162732
rect 206284 150408 206336 150414
rect 206284 150350 206336 150356
rect 204996 143676 205048 143682
rect 204996 143618 205048 143624
rect 204904 89004 204956 89010
rect 204904 88946 204956 88952
rect 203708 88256 203760 88262
rect 203708 88198 203760 88204
rect 203616 87644 203668 87650
rect 203616 87586 203668 87592
rect 203524 6384 203576 6390
rect 203524 6326 203576 6332
rect 202144 3732 202196 3738
rect 202144 3674 202196 3680
rect 196624 3664 196676 3670
rect 196624 3606 196676 3612
rect 203628 3534 203656 87586
rect 205008 81122 205036 143618
rect 206284 140820 206336 140826
rect 206284 140762 206336 140768
rect 204996 81116 205048 81122
rect 204996 81058 205048 81064
rect 206296 78538 206324 140762
rect 206376 139460 206428 139466
rect 206376 139402 206428 139408
rect 206388 86902 206416 139402
rect 206468 100768 206520 100774
rect 206468 100710 206520 100716
rect 206376 86896 206428 86902
rect 206376 86838 206428 86844
rect 206284 78532 206336 78538
rect 206284 78474 206336 78480
rect 206480 73166 206508 100710
rect 207032 83502 207060 239822
rect 207664 150476 207716 150482
rect 207664 150418 207716 150424
rect 207676 111790 207704 150418
rect 207664 111784 207716 111790
rect 207664 111726 207716 111732
rect 207664 107772 207716 107778
rect 207664 107714 207716 107720
rect 207020 83496 207072 83502
rect 207020 83438 207072 83444
rect 207676 80034 207704 107714
rect 207756 102264 207808 102270
rect 207756 102206 207808 102212
rect 207768 93838 207796 102206
rect 207848 96688 207900 96694
rect 207848 96630 207900 96636
rect 207756 93832 207808 93838
rect 207756 93774 207808 93780
rect 207860 89622 207888 96630
rect 207848 89616 207900 89622
rect 207848 89558 207900 89564
rect 207664 80028 207716 80034
rect 207664 79970 207716 79976
rect 206468 73160 206520 73166
rect 206468 73102 206520 73108
rect 208412 24274 208440 240094
rect 210620 233170 210648 240094
rect 210608 233164 210660 233170
rect 210608 233106 210660 233112
rect 210424 214804 210476 214810
rect 210424 214746 210476 214752
rect 210436 178906 210464 214746
rect 211068 190120 211120 190126
rect 211068 190062 211120 190068
rect 210608 184952 210660 184958
rect 210608 184894 210660 184900
rect 210424 178900 210476 178906
rect 210424 178842 210476 178848
rect 210516 171148 210568 171154
rect 210516 171090 210568 171096
rect 210424 151088 210476 151094
rect 210424 151030 210476 151036
rect 209044 141432 209096 141438
rect 209044 141374 209096 141380
rect 209056 93838 209084 141374
rect 209044 93832 209096 93838
rect 209044 93774 209096 93780
rect 208400 24268 208452 24274
rect 208400 24210 208452 24216
rect 210436 3534 210464 151030
rect 210528 150346 210556 171090
rect 210620 166870 210648 184894
rect 210608 166864 210660 166870
rect 210608 166806 210660 166812
rect 210516 150340 210568 150346
rect 210516 150282 210568 150288
rect 210516 140888 210568 140894
rect 210516 140830 210568 140836
rect 210528 82754 210556 140830
rect 210516 82748 210568 82754
rect 210516 82690 210568 82696
rect 211080 11966 211108 190062
rect 211804 150544 211856 150550
rect 211804 150486 211856 150492
rect 211816 137290 211844 150486
rect 211804 137284 211856 137290
rect 211804 137226 211856 137232
rect 211896 125724 211948 125730
rect 211896 125666 211948 125672
rect 211804 106412 211856 106418
rect 211804 106354 211856 106360
rect 211816 84182 211844 106354
rect 211804 84176 211856 84182
rect 211804 84118 211856 84124
rect 211804 79348 211856 79354
rect 211804 79290 211856 79296
rect 211068 11960 211120 11966
rect 211068 11902 211120 11908
rect 203616 3528 203668 3534
rect 203616 3470 203668 3476
rect 210424 3528 210476 3534
rect 210424 3470 210476 3476
rect 211816 3466 211844 79290
rect 211908 78606 211936 125666
rect 211988 123412 212040 123418
rect 211988 123354 212040 123360
rect 212000 79898 212028 123354
rect 211988 79892 212040 79898
rect 211988 79834 212040 79840
rect 211896 78600 211948 78606
rect 211896 78542 211948 78548
rect 212552 14618 212580 240094
rect 215312 238814 215340 240094
rect 215300 238808 215352 238814
rect 215300 238750 215352 238756
rect 217060 237454 217088 240094
rect 215944 237448 215996 237454
rect 215944 237390 215996 237396
rect 217048 237448 217100 237454
rect 217048 237390 217100 237396
rect 214564 221672 214616 221678
rect 214564 221614 214616 221620
rect 214576 184385 214604 221614
rect 214656 189100 214708 189106
rect 214656 189042 214708 189048
rect 214562 184376 214618 184385
rect 214562 184311 214618 184320
rect 213920 176656 213972 176662
rect 213920 176598 213972 176604
rect 213932 175681 213960 176598
rect 214012 175976 214064 175982
rect 214012 175918 214064 175924
rect 213918 175672 213974 175681
rect 213918 175607 213974 175616
rect 213920 175228 213972 175234
rect 213920 175170 213972 175176
rect 213932 175001 213960 175170
rect 213918 174992 213974 175001
rect 213918 174927 213974 174936
rect 213920 174548 213972 174554
rect 213920 174490 213972 174496
rect 213932 173641 213960 174490
rect 213918 173632 213974 173641
rect 213918 173567 213974 173576
rect 214024 172961 214052 175918
rect 214668 174321 214696 189042
rect 214748 183592 214800 183598
rect 214748 183534 214800 183540
rect 214654 174312 214710 174321
rect 214654 174247 214710 174256
rect 214288 173188 214340 173194
rect 214288 173130 214340 173136
rect 214010 172952 214066 172961
rect 214010 172887 214066 172896
rect 213920 172508 213972 172514
rect 213920 172450 213972 172456
rect 213932 172281 213960 172450
rect 213918 172272 213974 172281
rect 213918 172207 213974 172216
rect 214300 171134 214328 173130
rect 214760 171601 214788 183534
rect 214932 178084 214984 178090
rect 214932 178026 214984 178032
rect 214746 171592 214802 171601
rect 214746 171527 214802 171536
rect 214300 171106 214604 171134
rect 214012 171080 214064 171086
rect 213918 171048 213974 171057
rect 214012 171022 214064 171028
rect 213918 170983 213920 170992
rect 213972 170983 213974 170992
rect 213920 170954 213972 170960
rect 214024 170377 214052 171022
rect 214010 170368 214066 170377
rect 214010 170303 214066 170312
rect 214012 168360 214064 168366
rect 213918 168328 213974 168337
rect 214012 168302 214064 168308
rect 213918 168263 213920 168272
rect 213972 168263 213974 168272
rect 213920 168234 213972 168240
rect 214024 167657 214052 168302
rect 214010 167648 214066 167657
rect 214010 167583 214066 167592
rect 214012 167000 214064 167006
rect 214012 166942 214064 166948
rect 214102 166968 214158 166977
rect 213920 166932 213972 166938
rect 213920 166874 213972 166880
rect 213932 166433 213960 166874
rect 213918 166424 213974 166433
rect 213918 166359 213974 166368
rect 214024 165753 214052 166942
rect 214102 166903 214158 166912
rect 214116 166870 214144 166903
rect 214104 166864 214156 166870
rect 214104 166806 214156 166812
rect 214010 165744 214066 165753
rect 214010 165679 214066 165688
rect 213920 165572 213972 165578
rect 213920 165514 213972 165520
rect 213932 165073 213960 165514
rect 214012 165504 214064 165510
rect 214012 165446 214064 165452
rect 213918 165064 213974 165073
rect 213918 164999 213974 165008
rect 214024 164393 214052 165446
rect 214010 164384 214066 164393
rect 214010 164319 214066 164328
rect 213920 164212 213972 164218
rect 213920 164154 213972 164160
rect 213932 163713 213960 164154
rect 214012 164144 214064 164150
rect 214012 164086 214064 164092
rect 213918 163704 213974 163713
rect 213918 163639 213974 163648
rect 214024 163033 214052 164086
rect 214010 163024 214066 163033
rect 214010 162959 214066 162968
rect 213920 162852 213972 162858
rect 213920 162794 213972 162800
rect 213932 162353 213960 162794
rect 214012 162784 214064 162790
rect 214012 162726 214064 162732
rect 213918 162344 213974 162353
rect 213918 162279 213974 162288
rect 214024 161809 214052 162726
rect 214010 161800 214066 161809
rect 214010 161735 214066 161744
rect 213920 161424 213972 161430
rect 213920 161366 213972 161372
rect 213932 160449 213960 161366
rect 214576 161129 214604 171106
rect 214944 169697 214972 178026
rect 214930 169688 214986 169697
rect 214930 169623 214986 169632
rect 214656 169040 214708 169046
rect 214656 168982 214708 168988
rect 214562 161120 214618 161129
rect 214562 161055 214618 161064
rect 214102 160712 214158 160721
rect 214102 160647 214158 160656
rect 213918 160440 213974 160449
rect 213918 160375 213974 160384
rect 213920 160064 213972 160070
rect 213920 160006 213972 160012
rect 213932 159769 213960 160006
rect 214012 159996 214064 160002
rect 214012 159938 214064 159944
rect 213918 159760 213974 159769
rect 213918 159695 213974 159704
rect 214024 159089 214052 159938
rect 214010 159080 214066 159089
rect 214010 159015 214066 159024
rect 213920 158704 213972 158710
rect 213920 158646 213972 158652
rect 213932 157729 213960 158646
rect 213918 157720 213974 157729
rect 213918 157655 213974 157664
rect 213920 157344 213972 157350
rect 213920 157286 213972 157292
rect 213932 156505 213960 157286
rect 214116 157185 214144 160647
rect 214668 158409 214696 168982
rect 214654 158400 214710 158409
rect 214654 158335 214710 158344
rect 214102 157176 214158 157185
rect 214102 157111 214158 157120
rect 213918 156496 213974 156505
rect 213918 156431 213974 156440
rect 214012 155916 214064 155922
rect 214012 155858 214064 155864
rect 213920 155848 213972 155854
rect 213918 155816 213920 155825
rect 213972 155816 213974 155825
rect 213918 155751 213974 155760
rect 214024 155145 214052 155858
rect 214010 155136 214066 155145
rect 214010 155071 214066 155080
rect 214010 154456 214066 154465
rect 214010 154391 214066 154400
rect 213918 153776 213974 153785
rect 213918 153711 213974 153720
rect 213932 153270 213960 153711
rect 214024 153338 214052 154391
rect 214012 153332 214064 153338
rect 214012 153274 214064 153280
rect 213920 153264 213972 153270
rect 213920 153206 213972 153212
rect 213918 153096 213974 153105
rect 213918 153031 213974 153040
rect 213932 151910 213960 153031
rect 214010 152552 214066 152561
rect 214010 152487 214066 152496
rect 213920 151904 213972 151910
rect 213920 151846 213972 151852
rect 214024 151842 214052 152487
rect 214378 151872 214434 151881
rect 214012 151836 214064 151842
rect 214378 151807 214434 151816
rect 214012 151778 214064 151784
rect 214010 151192 214066 151201
rect 214010 151127 214066 151136
rect 214024 150550 214052 151127
rect 214012 150544 214064 150550
rect 213918 150512 213974 150521
rect 214012 150486 214064 150492
rect 213918 150447 213920 150456
rect 213972 150447 213974 150456
rect 213920 150418 213972 150424
rect 214012 150408 214064 150414
rect 214012 150350 214064 150356
rect 213920 150340 213972 150346
rect 213920 150282 213972 150288
rect 213932 149161 213960 150282
rect 214024 149841 214052 150350
rect 214010 149832 214066 149841
rect 214010 149767 214066 149776
rect 213918 149152 213974 149161
rect 213918 149087 213974 149096
rect 213920 149048 213972 149054
rect 213920 148990 213972 148996
rect 213932 148481 213960 148990
rect 213918 148472 213974 148481
rect 213918 148407 213974 148416
rect 213918 147928 213974 147937
rect 213918 147863 213974 147872
rect 213932 147694 213960 147863
rect 213920 147688 213972 147694
rect 213920 147630 213972 147636
rect 214010 147248 214066 147257
rect 214010 147183 214066 147192
rect 213918 146568 213974 146577
rect 213918 146503 213974 146512
rect 213932 146402 213960 146503
rect 213920 146396 213972 146402
rect 213920 146338 213972 146344
rect 214024 146334 214052 147183
rect 214012 146328 214064 146334
rect 214012 146270 214064 146276
rect 214010 145888 214066 145897
rect 214010 145823 214066 145832
rect 213918 145208 213974 145217
rect 213918 145143 213974 145152
rect 213932 145042 213960 145143
rect 213920 145036 213972 145042
rect 213920 144978 213972 144984
rect 214024 144974 214052 145823
rect 214392 145586 214420 151807
rect 214380 145580 214432 145586
rect 214380 145522 214432 145528
rect 214012 144968 214064 144974
rect 214012 144910 214064 144916
rect 214010 144528 214066 144537
rect 214010 144463 214066 144472
rect 213918 143848 213974 143857
rect 213918 143783 213974 143792
rect 213932 143614 213960 143783
rect 214024 143682 214052 144463
rect 214012 143676 214064 143682
rect 214012 143618 214064 143624
rect 213920 143608 213972 143614
rect 213920 143550 213972 143556
rect 213918 143304 213974 143313
rect 213918 143239 213974 143248
rect 213932 142186 213960 143239
rect 214746 142624 214802 142633
rect 214746 142559 214802 142568
rect 213920 142180 213972 142186
rect 213920 142122 213972 142128
rect 213918 141944 213974 141953
rect 213918 141879 213974 141888
rect 213932 140826 213960 141879
rect 214010 141264 214066 141273
rect 214010 141199 214066 141208
rect 214024 140894 214052 141199
rect 214012 140888 214064 140894
rect 214012 140830 214064 140836
rect 213920 140820 213972 140826
rect 213920 140762 213972 140768
rect 213918 140584 213974 140593
rect 213918 140519 213974 140528
rect 213182 139904 213238 139913
rect 213182 139839 213238 139848
rect 213196 85474 213224 139839
rect 213932 139466 213960 140519
rect 213920 139460 213972 139466
rect 213920 139402 213972 139408
rect 214010 139224 214066 139233
rect 214010 139159 214066 139168
rect 213918 138680 213974 138689
rect 213918 138615 213974 138624
rect 213932 138106 213960 138615
rect 213920 138100 213972 138106
rect 213920 138042 213972 138048
rect 214024 138038 214052 139159
rect 214012 138032 214064 138038
rect 214012 137974 214064 137980
rect 214654 138000 214710 138009
rect 214654 137935 214710 137944
rect 213918 137320 213974 137329
rect 213918 137255 213974 137264
rect 213932 136678 213960 137255
rect 213920 136672 213972 136678
rect 213920 136614 213972 136620
rect 214562 136640 214618 136649
rect 214562 136575 214618 136584
rect 214010 135960 214066 135969
rect 214010 135895 214066 135904
rect 214024 135386 214052 135895
rect 214012 135380 214064 135386
rect 214012 135322 214064 135328
rect 213920 135312 213972 135318
rect 213918 135280 213920 135289
rect 213972 135280 213974 135289
rect 213918 135215 213974 135224
rect 213920 133952 213972 133958
rect 213918 133920 213920 133929
rect 213972 133920 213974 133929
rect 213918 133855 213974 133864
rect 213918 133376 213974 133385
rect 213918 133311 213974 133320
rect 213932 132530 213960 133311
rect 213920 132524 213972 132530
rect 213920 132466 213972 132472
rect 213918 131336 213974 131345
rect 213918 131271 213974 131280
rect 213932 131170 213960 131271
rect 213920 131164 213972 131170
rect 213920 131106 213972 131112
rect 213918 129976 213974 129985
rect 213918 129911 213974 129920
rect 213932 129810 213960 129911
rect 213920 129804 213972 129810
rect 213920 129746 213972 129752
rect 213918 129296 213974 129305
rect 213918 129231 213974 129240
rect 213932 128382 213960 129231
rect 213920 128376 213972 128382
rect 213920 128318 213972 128324
rect 214010 128072 214066 128081
rect 214010 128007 214066 128016
rect 213918 127392 213974 127401
rect 213918 127327 213974 127336
rect 213932 127090 213960 127327
rect 213920 127084 213972 127090
rect 213920 127026 213972 127032
rect 214024 127022 214052 128007
rect 214012 127016 214064 127022
rect 214012 126958 214064 126964
rect 213918 126712 213974 126721
rect 213918 126647 213974 126656
rect 213932 125662 213960 126647
rect 214470 126032 214526 126041
rect 214470 125967 214526 125976
rect 214484 125730 214512 125967
rect 214472 125724 214524 125730
rect 214472 125666 214524 125672
rect 213920 125656 213972 125662
rect 213920 125598 213972 125604
rect 214010 125352 214066 125361
rect 214010 125287 214066 125296
rect 213918 124672 213974 124681
rect 213918 124607 213974 124616
rect 213932 124234 213960 124607
rect 214024 124302 214052 125287
rect 214012 124296 214064 124302
rect 214012 124238 214064 124244
rect 213920 124228 213972 124234
rect 213920 124170 213972 124176
rect 214010 124128 214066 124137
rect 214010 124063 214066 124072
rect 213918 123448 213974 123457
rect 214024 123418 214052 124063
rect 213918 123383 213974 123392
rect 214012 123412 214064 123418
rect 213932 122874 213960 123383
rect 214012 123354 214064 123360
rect 213920 122868 213972 122874
rect 213920 122810 213972 122816
rect 214010 122768 214066 122777
rect 214010 122703 214066 122712
rect 213918 122088 213974 122097
rect 213918 122023 213974 122032
rect 213932 121582 213960 122023
rect 213920 121576 213972 121582
rect 213920 121518 213972 121524
rect 214024 121514 214052 122703
rect 214012 121508 214064 121514
rect 214012 121450 214064 121456
rect 214010 121408 214066 121417
rect 214010 121343 214066 121352
rect 213918 120728 213974 120737
rect 213918 120663 213974 120672
rect 213932 120154 213960 120663
rect 214024 120222 214052 121343
rect 214012 120216 214064 120222
rect 214012 120158 214064 120164
rect 213920 120148 213972 120154
rect 213920 120090 213972 120096
rect 214102 120048 214158 120057
rect 214102 119983 214158 119992
rect 214010 119504 214066 119513
rect 214010 119439 214066 119448
rect 213920 118856 213972 118862
rect 213918 118824 213920 118833
rect 213972 118824 213974 118833
rect 214024 118794 214052 119439
rect 213918 118759 213974 118768
rect 214012 118788 214064 118794
rect 214012 118730 214064 118736
rect 214116 118726 214144 119983
rect 214104 118720 214156 118726
rect 214104 118662 214156 118668
rect 214010 118144 214066 118153
rect 214010 118079 214066 118088
rect 213918 117464 213974 117473
rect 214024 117434 214052 118079
rect 213918 117399 213974 117408
rect 214012 117428 214064 117434
rect 213932 117366 213960 117399
rect 214012 117370 214064 117376
rect 213920 117360 213972 117366
rect 213920 117302 213972 117308
rect 214010 116784 214066 116793
rect 214010 116719 214066 116728
rect 213918 116104 213974 116113
rect 214024 116074 214052 116719
rect 213918 116039 213974 116048
rect 214012 116068 214064 116074
rect 213932 116006 213960 116039
rect 214012 116010 214064 116016
rect 213920 116000 213972 116006
rect 213920 115942 213972 115948
rect 214010 115424 214066 115433
rect 214010 115359 214066 115368
rect 213918 114880 213974 114889
rect 213918 114815 213974 114824
rect 213932 114646 213960 114815
rect 213920 114640 213972 114646
rect 213920 114582 213972 114588
rect 214024 114578 214052 115359
rect 214012 114572 214064 114578
rect 214012 114514 214064 114520
rect 214010 114200 214066 114209
rect 214010 114135 214066 114144
rect 213918 113520 213974 113529
rect 213918 113455 213974 113464
rect 213932 113218 213960 113455
rect 214024 113286 214052 114135
rect 214012 113280 214064 113286
rect 214012 113222 214064 113228
rect 213920 113212 213972 113218
rect 213920 113154 213972 113160
rect 213918 112840 213974 112849
rect 213918 112775 213974 112784
rect 213932 111858 213960 112775
rect 213920 111852 213972 111858
rect 213920 111794 213972 111800
rect 214010 111480 214066 111489
rect 214010 111415 214066 111424
rect 213918 110800 213974 110809
rect 213918 110735 213974 110744
rect 213932 110498 213960 110735
rect 214024 110566 214052 111415
rect 214012 110560 214064 110566
rect 214012 110502 214064 110508
rect 213920 110492 213972 110498
rect 213920 110434 213972 110440
rect 213918 110256 213974 110265
rect 213918 110191 213974 110200
rect 213932 109070 213960 110191
rect 213920 109064 213972 109070
rect 213920 109006 213972 109012
rect 214010 108896 214066 108905
rect 214010 108831 214066 108840
rect 213918 108216 213974 108225
rect 213918 108151 213974 108160
rect 213932 107710 213960 108151
rect 214024 107778 214052 108831
rect 214012 107772 214064 107778
rect 214012 107714 214064 107720
rect 213920 107704 213972 107710
rect 213920 107646 213972 107652
rect 213918 107536 213974 107545
rect 213918 107471 213974 107480
rect 213932 106350 213960 107471
rect 214470 106856 214526 106865
rect 214470 106791 214526 106800
rect 214484 106418 214512 106791
rect 214472 106412 214524 106418
rect 214472 106354 214524 106360
rect 213920 106344 213972 106350
rect 213920 106286 213972 106292
rect 214010 106176 214066 106185
rect 214010 106111 214066 106120
rect 213918 105632 213974 105641
rect 213918 105567 213974 105576
rect 213932 104990 213960 105567
rect 213920 104984 213972 104990
rect 213920 104926 213972 104932
rect 214024 104922 214052 106111
rect 214012 104916 214064 104922
rect 214012 104858 214064 104864
rect 214010 104272 214066 104281
rect 214010 104207 214066 104216
rect 213920 103624 213972 103630
rect 213918 103592 213920 103601
rect 213972 103592 213974 103601
rect 214024 103562 214052 104207
rect 213918 103527 213974 103536
rect 214012 103556 214064 103562
rect 214012 103498 214064 103504
rect 214010 102912 214066 102921
rect 214010 102847 214066 102856
rect 214024 102270 214052 102847
rect 214012 102264 214064 102270
rect 213918 102232 213974 102241
rect 214012 102206 214064 102212
rect 213918 102167 213920 102176
rect 213972 102167 213974 102176
rect 213920 102138 213972 102144
rect 213918 101008 213974 101017
rect 213918 100943 213974 100952
rect 213932 100774 213960 100943
rect 213920 100768 213972 100774
rect 213920 100710 213972 100716
rect 214102 100328 214158 100337
rect 214102 100263 214158 100272
rect 213918 99648 213974 99657
rect 213918 99583 213974 99592
rect 213932 99414 213960 99583
rect 213920 99408 213972 99414
rect 213920 99350 213972 99356
rect 214010 98968 214066 98977
rect 214010 98903 214066 98912
rect 213918 98288 213974 98297
rect 213918 98223 213974 98232
rect 213932 98122 213960 98223
rect 213920 98116 213972 98122
rect 213920 98058 213972 98064
rect 214024 98054 214052 98903
rect 214012 98048 214064 98054
rect 214012 97990 214064 97996
rect 213918 97608 213974 97617
rect 213918 97543 213974 97552
rect 213932 96694 213960 97543
rect 213920 96688 213972 96694
rect 213920 96630 213972 96636
rect 214116 95946 214144 100263
rect 214576 97306 214604 136575
rect 214668 100026 214696 137935
rect 214760 130422 214788 142559
rect 214930 130656 214986 130665
rect 214930 130591 214986 130600
rect 214748 130416 214800 130422
rect 214748 130358 214800 130364
rect 214944 112470 214972 130591
rect 214932 112464 214984 112470
rect 214932 112406 214984 112412
rect 214746 112160 214802 112169
rect 214746 112095 214802 112104
rect 214656 100020 214708 100026
rect 214656 99962 214708 99968
rect 214564 97300 214616 97306
rect 214564 97242 214616 97248
rect 214654 96928 214710 96937
rect 214654 96863 214710 96872
rect 214562 96384 214618 96393
rect 214562 96319 214618 96328
rect 214104 95940 214156 95946
rect 214104 95882 214156 95888
rect 213184 85468 213236 85474
rect 213184 85410 213236 85416
rect 214576 77246 214604 96319
rect 214668 86970 214696 96863
rect 214656 86964 214708 86970
rect 214656 86906 214708 86912
rect 214760 79966 214788 112095
rect 214838 101552 214894 101561
rect 214838 101487 214894 101496
rect 214852 89690 214880 101487
rect 214840 89684 214892 89690
rect 214840 89626 214892 89632
rect 214748 79960 214800 79966
rect 214748 79902 214800 79908
rect 214564 77240 214616 77246
rect 214564 77182 214616 77188
rect 215956 17270 215984 237390
rect 218992 233238 219020 240094
rect 218980 233232 219032 233238
rect 218980 233174 219032 233180
rect 220084 227180 220136 227186
rect 220084 227122 220136 227128
rect 220096 183190 220124 227122
rect 220084 183184 220136 183190
rect 220084 183126 220136 183132
rect 220832 178022 220860 240094
rect 223822 239850 223850 240108
rect 224972 240094 225768 240122
rect 223822 239822 223896 239850
rect 223868 238678 223896 239822
rect 223856 238672 223908 238678
rect 223856 238614 223908 238620
rect 222844 235340 222896 235346
rect 222844 235282 222896 235288
rect 222856 184482 222884 235282
rect 223868 233238 223896 238614
rect 224132 237448 224184 237454
rect 224132 237390 224184 237396
rect 223856 233232 223908 233238
rect 223856 233174 223908 233180
rect 224144 231674 224172 237390
rect 224132 231668 224184 231674
rect 224132 231610 224184 231616
rect 224224 231124 224276 231130
rect 224224 231066 224276 231072
rect 222844 184476 222896 184482
rect 222844 184418 222896 184424
rect 224236 181626 224264 231066
rect 224224 181620 224276 181626
rect 224224 181562 224276 181568
rect 217968 178016 218020 178022
rect 217968 177958 218020 177964
rect 220820 178016 220872 178022
rect 220820 177958 220872 177964
rect 216588 177540 216640 177546
rect 216588 177482 216640 177488
rect 216036 140072 216088 140078
rect 216036 140014 216088 140020
rect 215944 17264 215996 17270
rect 215944 17206 215996 17212
rect 212540 14612 212592 14618
rect 212540 14554 212592 14560
rect 216048 3466 216076 140014
rect 216600 86290 216628 177482
rect 216588 86284 216640 86290
rect 216588 86226 216640 86232
rect 217980 17270 218008 177958
rect 224972 177546 225000 240094
rect 227686 239850 227714 240108
rect 229112 240094 229632 240122
rect 231872 240094 232208 240122
rect 233896 240094 234140 240122
rect 227686 239822 227760 239850
rect 227732 191214 227760 239822
rect 228364 206440 228416 206446
rect 228364 206382 228416 206388
rect 227720 191208 227772 191214
rect 227720 191150 227772 191156
rect 228376 181762 228404 206382
rect 229112 190058 229140 240094
rect 231872 210662 231900 240094
rect 233896 237250 233924 240094
rect 236058 239850 236086 240108
rect 236012 239822 236086 239850
rect 237392 240094 238004 240122
rect 240152 240094 240580 240122
rect 241532 240094 242512 240122
rect 244292 240094 244444 240122
rect 245672 240094 246376 240122
rect 248432 240094 248952 240122
rect 236012 238678 236040 239822
rect 236000 238672 236052 238678
rect 236000 238614 236052 238620
rect 233884 237244 233936 237250
rect 233884 237186 233936 237192
rect 233896 230314 233924 237186
rect 236012 233102 236040 238614
rect 236000 233096 236052 233102
rect 236000 233038 236052 233044
rect 233884 230308 233936 230314
rect 233884 230250 233936 230256
rect 236644 213444 236696 213450
rect 236644 213386 236696 213392
rect 231860 210656 231912 210662
rect 231860 210598 231912 210604
rect 232504 210588 232556 210594
rect 232504 210530 232556 210536
rect 231124 200796 231176 200802
rect 231124 200738 231176 200744
rect 229100 190052 229152 190058
rect 229100 189994 229152 190000
rect 228364 181756 228416 181762
rect 228364 181698 228416 181704
rect 231136 180334 231164 200738
rect 232516 185609 232544 210530
rect 232502 185600 232558 185609
rect 232502 185535 232558 185544
rect 231124 180328 231176 180334
rect 231124 180270 231176 180276
rect 236656 177682 236684 213386
rect 237392 208010 237420 240094
rect 240152 238754 240180 240094
rect 240060 238726 240180 238754
rect 240060 237454 240088 238726
rect 240048 237448 240100 237454
rect 240048 237390 240100 237396
rect 240060 233170 240088 237390
rect 240048 233164 240100 233170
rect 240048 233106 240100 233112
rect 241532 229022 241560 240094
rect 242256 236700 242308 236706
rect 242256 236642 242308 236648
rect 241520 229016 241572 229022
rect 241520 228958 241572 228964
rect 240784 222964 240836 222970
rect 240784 222906 240836 222912
rect 237380 208004 237432 208010
rect 237380 207946 237432 207952
rect 239404 207800 239456 207806
rect 239404 207742 239456 207748
rect 236644 177676 236696 177682
rect 236644 177618 236696 177624
rect 224960 177540 225012 177546
rect 224960 177482 225012 177488
rect 239416 177313 239444 207742
rect 239496 198212 239548 198218
rect 239496 198154 239548 198160
rect 239508 180169 239536 198154
rect 239494 180160 239550 180169
rect 239494 180095 239550 180104
rect 240796 178974 240824 222906
rect 242164 220312 242216 220318
rect 242164 220254 242216 220260
rect 240784 178968 240836 178974
rect 240784 178910 240836 178916
rect 242176 177546 242204 220254
rect 242268 210633 242296 236642
rect 242254 210624 242310 210633
rect 242254 210559 242310 210568
rect 243544 203856 243596 203862
rect 243544 203798 243596 203804
rect 242256 191412 242308 191418
rect 242256 191354 242308 191360
rect 242268 177614 242296 191354
rect 242256 177608 242308 177614
rect 242256 177550 242308 177556
rect 242164 177540 242216 177546
rect 242164 177482 242216 177488
rect 239402 177304 239458 177313
rect 239402 177239 239458 177248
rect 243556 175846 243584 203798
rect 244292 190126 244320 240094
rect 245672 202502 245700 240094
rect 247684 221604 247736 221610
rect 247684 221546 247736 221552
rect 246396 210520 246448 210526
rect 246396 210462 246448 210468
rect 246304 210452 246356 210458
rect 246304 210394 246356 210400
rect 245660 202496 245712 202502
rect 245660 202438 245712 202444
rect 244924 194200 244976 194206
rect 244924 194142 244976 194148
rect 244280 190120 244332 190126
rect 244280 190062 244332 190068
rect 244936 176089 244964 194142
rect 245660 183116 245712 183122
rect 245660 183058 245712 183064
rect 245672 176662 245700 183058
rect 245660 176656 245712 176662
rect 245660 176598 245712 176604
rect 244922 176080 244978 176089
rect 246316 176050 246344 210394
rect 246408 179042 246436 210462
rect 246396 179036 246448 179042
rect 246396 178978 246448 178984
rect 244922 176015 244978 176024
rect 246304 176044 246356 176050
rect 246304 175986 246356 175992
rect 247696 175982 247724 221546
rect 247776 209160 247828 209166
rect 247776 209102 247828 209108
rect 247788 177721 247816 209102
rect 248432 203862 248460 240094
rect 250870 239850 250898 240108
rect 250824 239822 250898 239850
rect 252572 240094 252816 240122
rect 254412 240094 254748 240122
rect 256712 240094 257324 240122
rect 258092 240094 259256 240122
rect 260852 240094 261188 240122
rect 262784 240094 263120 240122
rect 250824 238610 250852 239822
rect 252572 238950 252600 240094
rect 252560 238944 252612 238950
rect 252560 238886 252612 238892
rect 250812 238604 250864 238610
rect 250812 238546 250864 238552
rect 250824 238105 250852 238546
rect 250810 238096 250866 238105
rect 250810 238031 250866 238040
rect 254412 237182 254440 240094
rect 254400 237176 254452 237182
rect 254400 237118 254452 237124
rect 255964 233980 256016 233986
rect 255964 233922 256016 233928
rect 253204 225616 253256 225622
rect 253204 225558 253256 225564
rect 249800 223032 249852 223038
rect 249800 222974 249852 222980
rect 248420 203856 248472 203862
rect 248420 203798 248472 203804
rect 249064 187128 249116 187134
rect 249064 187070 249116 187076
rect 247774 177712 247830 177721
rect 247774 177647 247830 177656
rect 249076 176118 249104 187070
rect 249340 181688 249392 181694
rect 249340 181630 249392 181636
rect 249248 177676 249300 177682
rect 249248 177618 249300 177624
rect 249156 177404 249208 177410
rect 249156 177346 249208 177352
rect 249064 176112 249116 176118
rect 249064 176054 249116 176060
rect 247684 175976 247736 175982
rect 247684 175918 247736 175924
rect 243544 175840 243596 175846
rect 248052 175840 248104 175846
rect 243544 175782 243596 175788
rect 248050 175808 248052 175817
rect 248104 175808 248106 175817
rect 248050 175743 248106 175752
rect 249168 174729 249196 177346
rect 249154 174720 249210 174729
rect 249154 174655 249210 174664
rect 249260 172417 249288 177618
rect 249352 173369 249380 181630
rect 249338 173360 249394 173369
rect 249338 173295 249394 173304
rect 249246 172408 249302 172417
rect 249246 172343 249302 172352
rect 249812 138553 249840 222974
rect 252836 205080 252888 205086
rect 252836 205022 252888 205028
rect 252652 202360 252704 202366
rect 252652 202302 252704 202308
rect 250076 196988 250128 196994
rect 250076 196930 250128 196936
rect 249984 178900 250036 178906
rect 249984 178842 250036 178848
rect 249892 176656 249944 176662
rect 249892 176598 249944 176604
rect 249904 151814 249932 176598
rect 249996 171134 250024 178842
rect 250088 175273 250116 196930
rect 251180 196852 251232 196858
rect 251180 196794 251232 196800
rect 250074 175264 250130 175273
rect 250074 175199 250130 175208
rect 249996 171106 250116 171134
rect 250088 159225 250116 171106
rect 251088 159384 251140 159390
rect 251088 159326 251140 159332
rect 250074 159216 250130 159225
rect 250074 159151 250130 159160
rect 251100 154465 251128 159326
rect 251192 158817 251220 196794
rect 251272 180192 251324 180198
rect 251272 180134 251324 180140
rect 251284 159633 251312 180134
rect 252560 179036 252612 179042
rect 252560 178978 252612 178984
rect 251456 178832 251508 178838
rect 251456 178774 251508 178780
rect 251364 177472 251416 177478
rect 251364 177414 251416 177420
rect 251376 170950 251404 177414
rect 251364 170944 251416 170950
rect 251364 170886 251416 170892
rect 251364 170332 251416 170338
rect 251364 170274 251416 170280
rect 251376 170105 251404 170274
rect 251362 170096 251418 170105
rect 251362 170031 251418 170040
rect 251468 161474 251496 178774
rect 252100 173732 252152 173738
rect 252100 173674 252152 173680
rect 252112 172825 252140 173674
rect 252098 172816 252154 172825
rect 252098 172751 252154 172760
rect 252466 171864 252522 171873
rect 252466 171799 252522 171808
rect 252480 171562 252508 171799
rect 252468 171556 252520 171562
rect 252468 171498 252520 171504
rect 252572 171465 252600 178978
rect 252558 171456 252614 171465
rect 252558 171391 252614 171400
rect 252664 171134 252692 202302
rect 252744 187264 252796 187270
rect 252744 187206 252796 187212
rect 252572 171106 252692 171134
rect 251548 170944 251600 170950
rect 251732 170944 251784 170950
rect 251548 170886 251600 170892
rect 251730 170912 251732 170921
rect 251784 170912 251786 170921
rect 251376 161446 251496 161474
rect 251376 160177 251404 161446
rect 251362 160168 251418 160177
rect 251362 160103 251418 160112
rect 251270 159624 251326 159633
rect 251270 159559 251326 159568
rect 251178 158808 251234 158817
rect 251178 158743 251234 158752
rect 251560 156913 251588 170886
rect 251730 170847 251786 170856
rect 251822 170504 251878 170513
rect 251822 170439 251878 170448
rect 251836 169862 251864 170439
rect 251824 169856 251876 169862
rect 251824 169798 251876 169804
rect 252284 169720 252336 169726
rect 252284 169662 252336 169668
rect 252296 169153 252324 169662
rect 252466 169552 252522 169561
rect 252572 169538 252600 171106
rect 252522 169510 252600 169538
rect 252466 169487 252522 169496
rect 252756 169266 252784 187206
rect 252572 169238 252784 169266
rect 252282 169144 252338 169153
rect 252282 169079 252338 169088
rect 251916 168360 251968 168366
rect 251916 168302 251968 168308
rect 251928 167249 251956 168302
rect 252466 168192 252522 168201
rect 252572 168178 252600 169238
rect 252522 168150 252600 168178
rect 252466 168127 252522 168136
rect 252466 167648 252522 167657
rect 252466 167583 252522 167592
rect 252480 167278 252508 167583
rect 252468 167272 252520 167278
rect 251914 167240 251970 167249
rect 252468 167214 252520 167220
rect 251914 167175 251970 167184
rect 252100 167000 252152 167006
rect 252100 166942 252152 166948
rect 252112 166705 252140 166942
rect 252376 166796 252428 166802
rect 252376 166738 252428 166744
rect 252098 166696 252154 166705
rect 252098 166631 252154 166640
rect 252388 166433 252416 166738
rect 252468 166524 252520 166530
rect 252468 166466 252520 166472
rect 252374 166424 252430 166433
rect 252374 166359 252430 166368
rect 252480 165753 252508 166466
rect 252466 165744 252522 165753
rect 252466 165679 252522 165688
rect 252468 165572 252520 165578
rect 252468 165514 252520 165520
rect 252100 165504 252152 165510
rect 252100 165446 252152 165452
rect 251732 165436 251784 165442
rect 251732 165378 251784 165384
rect 251744 164801 251772 165378
rect 251730 164792 251786 164801
rect 251730 164727 251786 164736
rect 252112 164393 252140 165446
rect 252480 165345 252508 165514
rect 252466 165336 252522 165345
rect 252466 165271 252522 165280
rect 252098 164384 252154 164393
rect 252098 164319 252154 164328
rect 252192 164212 252244 164218
rect 252192 164154 252244 164160
rect 252204 163033 252232 164154
rect 252190 163024 252246 163033
rect 252190 162959 252246 162968
rect 252468 162852 252520 162858
rect 252468 162794 252520 162800
rect 252480 162489 252508 162794
rect 252466 162480 252522 162489
rect 252466 162415 252522 162424
rect 252848 161474 252876 205022
rect 253216 194206 253244 225558
rect 255320 216164 255372 216170
rect 255320 216106 255372 216112
rect 253204 194200 253256 194206
rect 253204 194142 253256 194148
rect 254124 192568 254176 192574
rect 254124 192510 254176 192516
rect 254032 189780 254084 189786
rect 254032 189722 254084 189728
rect 253940 176112 253992 176118
rect 253940 176054 253992 176060
rect 253952 170338 253980 176054
rect 253940 170332 253992 170338
rect 253940 170274 253992 170280
rect 253202 163976 253258 163985
rect 253202 163911 253258 163920
rect 253216 163033 253244 163911
rect 253202 163024 253258 163033
rect 253202 162959 253258 162968
rect 252572 161446 252876 161474
rect 252468 161424 252520 161430
rect 252468 161366 252520 161372
rect 252480 160585 252508 161366
rect 252466 160576 252522 160585
rect 252466 160511 252522 160520
rect 251916 158704 251968 158710
rect 251916 158646 251968 158652
rect 251928 157865 251956 158646
rect 251914 157856 251970 157865
rect 251914 157791 251970 157800
rect 252468 157344 252520 157350
rect 252466 157312 252468 157321
rect 252520 157312 252522 157321
rect 252376 157276 252428 157282
rect 252466 157247 252522 157256
rect 252376 157218 252428 157224
rect 251546 156904 251602 156913
rect 251546 156839 251602 156848
rect 252388 156369 252416 157218
rect 252374 156360 252430 156369
rect 252374 156295 252430 156304
rect 251914 155952 251970 155961
rect 251914 155887 251916 155896
rect 251968 155887 251970 155896
rect 251916 155858 251968 155864
rect 251180 155848 251232 155854
rect 251180 155790 251232 155796
rect 251192 155417 251220 155790
rect 252468 155780 252520 155786
rect 252468 155722 252520 155728
rect 251178 155408 251234 155417
rect 251178 155343 251234 155352
rect 252480 155009 252508 155722
rect 252466 155000 252522 155009
rect 252466 154935 252522 154944
rect 251640 154556 251692 154562
rect 251640 154498 251692 154504
rect 251086 154456 251142 154465
rect 251086 154391 251142 154400
rect 251652 154057 251680 154498
rect 251638 154048 251694 154057
rect 251638 153983 251694 153992
rect 252466 153504 252522 153513
rect 252572 153490 252600 161446
rect 254044 155854 254072 189722
rect 254032 155848 254084 155854
rect 254032 155790 254084 155796
rect 252522 153462 252600 153490
rect 252466 153439 252522 153448
rect 251916 153196 251968 153202
rect 251916 153138 251968 153144
rect 250534 152960 250590 152969
rect 250534 152895 250590 152904
rect 249904 151786 250024 151814
rect 249996 141409 250024 151786
rect 249982 141400 250038 141409
rect 249982 141335 250038 141344
rect 249798 138544 249854 138553
rect 249798 138479 249854 138488
rect 250444 138032 250496 138038
rect 250444 137974 250496 137980
rect 249064 136672 249116 136678
rect 249064 136614 249116 136620
rect 246948 94512 247000 94518
rect 241518 94480 241574 94489
rect 246948 94454 247000 94460
rect 241518 94415 241574 94424
rect 238760 93152 238812 93158
rect 238760 93094 238812 93100
rect 228364 91792 228416 91798
rect 228364 91734 228416 91740
rect 224224 89208 224276 89214
rect 224224 89150 224276 89156
rect 217968 17264 218020 17270
rect 217968 17206 218020 17212
rect 224236 3602 224264 89150
rect 228376 11830 228404 91734
rect 238024 86352 238076 86358
rect 238024 86294 238076 86300
rect 228364 11824 228416 11830
rect 228364 11766 228416 11772
rect 224224 3596 224276 3602
rect 224224 3538 224276 3544
rect 211804 3460 211856 3466
rect 211804 3402 211856 3408
rect 216036 3460 216088 3466
rect 216036 3402 216088 3408
rect 238036 2990 238064 86294
rect 238772 16574 238800 93094
rect 241532 16574 241560 94415
rect 242900 89140 242952 89146
rect 242900 89082 242952 89088
rect 238772 16546 239352 16574
rect 241532 16546 241744 16574
rect 235816 2984 235868 2990
rect 235816 2926 235868 2932
rect 238024 2984 238076 2990
rect 238024 2926 238076 2932
rect 179328 2168 179380 2174
rect 179328 2110 179380 2116
rect 235828 480 235856 2926
rect 239324 480 239352 16546
rect 240508 3460 240560 3466
rect 240508 3402 240560 3408
rect 240520 480 240548 3402
rect 241716 480 241744 16546
rect 242912 3534 242940 89082
rect 245660 89072 245712 89078
rect 245660 89014 245712 89020
rect 245672 16574 245700 89014
rect 245672 16546 245976 16574
rect 242900 3528 242952 3534
rect 242900 3470 242952 3476
rect 244096 3528 244148 3534
rect 244096 3470 244148 3476
rect 242898 3360 242954 3369
rect 242898 3295 242954 3304
rect 242912 480 242940 3295
rect 244108 480 244136 3470
rect 245200 3460 245252 3466
rect 245200 3402 245252 3408
rect 245212 480 245240 3402
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 16546
rect 246960 3534 246988 94454
rect 247684 80776 247736 80782
rect 247684 80718 247736 80724
rect 247040 17332 247092 17338
rect 247040 17274 247092 17280
rect 247052 16574 247080 17274
rect 247052 16546 247632 16574
rect 246948 3528 247000 3534
rect 246948 3470 247000 3476
rect 247604 480 247632 16546
rect 247696 3466 247724 80718
rect 249076 20058 249104 136614
rect 249154 97064 249210 97073
rect 249154 96999 249210 97008
rect 249168 35902 249196 96999
rect 250456 47666 250484 137974
rect 250548 136649 250576 152895
rect 251928 152153 251956 153138
rect 252376 153128 252428 153134
rect 252376 153070 252428 153076
rect 252466 153096 252522 153105
rect 252388 152697 252416 153070
rect 252466 153031 252468 153040
rect 252520 153031 252522 153040
rect 252468 153002 252520 153008
rect 252374 152688 252430 152697
rect 252374 152623 252430 152632
rect 251914 152144 251970 152153
rect 251914 152079 251970 152088
rect 253480 151836 253532 151842
rect 253480 151778 253532 151784
rect 251916 151768 251968 151774
rect 251916 151710 251968 151716
rect 252466 151736 252522 151745
rect 251928 150793 251956 151710
rect 252376 151700 252428 151706
rect 252466 151671 252522 151680
rect 252376 151642 252428 151648
rect 252388 151201 252416 151642
rect 252480 151638 252508 151671
rect 252468 151632 252520 151638
rect 252468 151574 252520 151580
rect 252374 151192 252430 151201
rect 252374 151127 252430 151136
rect 251914 150784 251970 150793
rect 251914 150719 251970 150728
rect 251180 150408 251232 150414
rect 251180 150350 251232 150356
rect 251192 149841 251220 150350
rect 252008 150340 252060 150346
rect 252008 150282 252060 150288
rect 251178 149832 251234 149841
rect 251178 149767 251234 149776
rect 252020 149297 252048 150282
rect 252468 150272 252520 150278
rect 252466 150240 252468 150249
rect 252520 150240 252522 150249
rect 252466 150175 252522 150184
rect 252006 149288 252062 149297
rect 252006 149223 252062 149232
rect 253204 149116 253256 149122
rect 253204 149058 253256 149064
rect 252468 149048 252520 149054
rect 252468 148990 252520 148996
rect 251916 148912 251968 148918
rect 251914 148880 251916 148889
rect 251968 148880 251970 148889
rect 251914 148815 251970 148824
rect 252284 148640 252336 148646
rect 252284 148582 252336 148588
rect 251916 146940 251968 146946
rect 251916 146882 251968 146888
rect 251824 146124 251876 146130
rect 251824 146066 251876 146072
rect 251836 143177 251864 146066
rect 251822 143168 251878 143177
rect 251822 143103 251878 143112
rect 250628 142860 250680 142866
rect 250628 142802 250680 142808
rect 250534 136640 250590 136649
rect 250534 136575 250590 136584
rect 250536 96688 250588 96694
rect 250536 96630 250588 96636
rect 250444 47660 250496 47666
rect 250444 47602 250496 47608
rect 249156 35896 249208 35902
rect 249156 35838 249208 35844
rect 250548 26926 250576 96630
rect 250640 93158 250668 142802
rect 251928 142154 251956 146882
rect 252100 146192 252152 146198
rect 252100 146134 252152 146140
rect 252112 145081 252140 146134
rect 252296 145625 252324 148582
rect 252480 148345 252508 148990
rect 252466 148336 252522 148345
rect 252466 148271 252522 148280
rect 252468 147620 252520 147626
rect 252468 147562 252520 147568
rect 252376 147552 252428 147558
rect 252480 147529 252508 147562
rect 252376 147494 252428 147500
rect 252466 147520 252522 147529
rect 252388 146577 252416 147494
rect 252466 147455 252522 147464
rect 252374 146568 252430 146577
rect 252374 146503 252430 146512
rect 252468 146260 252520 146266
rect 252468 146202 252520 146208
rect 252480 146033 252508 146202
rect 252466 146024 252522 146033
rect 252466 145959 252522 145968
rect 252282 145616 252338 145625
rect 252282 145551 252338 145560
rect 252284 145512 252336 145518
rect 252284 145454 252336 145460
rect 252098 145072 252154 145081
rect 252098 145007 252154 145016
rect 252100 144900 252152 144906
rect 252100 144842 252152 144848
rect 252112 143721 252140 144842
rect 252098 143712 252154 143721
rect 252098 143647 252154 143656
rect 252296 142769 252324 145454
rect 252468 144832 252520 144838
rect 252468 144774 252520 144780
rect 252480 144129 252508 144774
rect 252466 144120 252522 144129
rect 252466 144055 252522 144064
rect 252282 142760 252338 142769
rect 252282 142695 252338 142704
rect 251836 142126 251956 142154
rect 251640 135244 251692 135250
rect 251640 135186 251692 135192
rect 251652 134745 251680 135186
rect 251638 134736 251694 134745
rect 251638 134671 251694 134680
rect 251456 133884 251508 133890
rect 251456 133826 251508 133832
rect 251468 133385 251496 133826
rect 251454 133376 251510 133385
rect 251454 133311 251510 133320
rect 251548 132184 251600 132190
rect 251548 132126 251600 132132
rect 251560 131889 251588 132126
rect 251546 131880 251602 131889
rect 251546 131815 251602 131824
rect 251548 131028 251600 131034
rect 251548 130970 251600 130976
rect 251560 130937 251588 130970
rect 251546 130928 251602 130937
rect 251546 130863 251602 130872
rect 251836 130121 251864 142126
rect 252100 140752 252152 140758
rect 252100 140694 252152 140700
rect 252112 140457 252140 140694
rect 252098 140448 252154 140457
rect 252098 140383 252154 140392
rect 252284 139868 252336 139874
rect 252284 139810 252336 139816
rect 252100 137896 252152 137902
rect 252100 137838 252152 137844
rect 252112 137601 252140 137838
rect 252098 137592 252154 137601
rect 252098 137527 252154 137536
rect 252192 137148 252244 137154
rect 252192 137090 252244 137096
rect 252100 136536 252152 136542
rect 252100 136478 252152 136484
rect 252112 136241 252140 136478
rect 252098 136232 252154 136241
rect 252098 136167 252154 136176
rect 251916 135924 251968 135930
rect 251916 135866 251968 135872
rect 251822 130112 251878 130121
rect 251822 130047 251878 130056
rect 251928 129962 251956 135866
rect 252008 133748 252060 133754
rect 252008 133690 252060 133696
rect 252020 132841 252048 133690
rect 252006 132832 252062 132841
rect 252006 132767 252062 132776
rect 252204 132682 252232 137090
rect 251836 129934 251956 129962
rect 252020 132654 252232 132682
rect 251732 129736 251784 129742
rect 251732 129678 251784 129684
rect 251744 129169 251772 129678
rect 251730 129160 251786 129169
rect 251730 129095 251786 129104
rect 251836 127786 251864 129934
rect 252020 129826 252048 132654
rect 252296 131481 252324 139810
rect 252466 138000 252522 138009
rect 252376 137964 252428 137970
rect 252466 137935 252522 137944
rect 252376 137906 252428 137912
rect 252388 137057 252416 137906
rect 252480 137834 252508 137935
rect 252468 137828 252520 137834
rect 252468 137770 252520 137776
rect 252374 137048 252430 137057
rect 252374 136983 252430 136992
rect 252376 136604 252428 136610
rect 252376 136546 252428 136552
rect 252388 135697 252416 136546
rect 252468 136468 252520 136474
rect 252468 136410 252520 136416
rect 252374 135688 252430 135697
rect 252374 135623 252430 135632
rect 252480 135289 252508 136410
rect 252466 135280 252522 135289
rect 252466 135215 252522 135224
rect 252468 135176 252520 135182
rect 252468 135118 252520 135124
rect 252480 134337 252508 135118
rect 252466 134328 252522 134337
rect 252466 134263 252522 134272
rect 252468 133816 252520 133822
rect 252466 133784 252468 133793
rect 252520 133784 252522 133793
rect 252466 133719 252522 133728
rect 252468 132456 252520 132462
rect 252466 132424 252468 132433
rect 252520 132424 252522 132433
rect 252466 132359 252522 132368
rect 252282 131472 252338 131481
rect 252282 131407 252338 131416
rect 252468 131096 252520 131102
rect 252468 131038 252520 131044
rect 252480 130529 252508 131038
rect 252466 130520 252522 130529
rect 252466 130455 252522 130464
rect 251744 127758 251864 127786
rect 251928 129798 252048 129826
rect 251272 126268 251324 126274
rect 251272 126210 251324 126216
rect 251180 125384 251232 125390
rect 251178 125352 251180 125361
rect 251232 125352 251234 125361
rect 251178 125287 251234 125296
rect 251284 124817 251312 126210
rect 251270 124808 251326 124817
rect 251270 124743 251326 124752
rect 251744 123049 251772 127758
rect 251824 127628 251876 127634
rect 251824 127570 251876 127576
rect 251730 123040 251786 123049
rect 251730 122975 251786 122984
rect 251836 118833 251864 127570
rect 251928 126313 251956 129798
rect 252008 129668 252060 129674
rect 252008 129610 252060 129616
rect 252020 128625 252048 129610
rect 252468 129600 252520 129606
rect 252466 129568 252468 129577
rect 252520 129568 252522 129577
rect 252466 129503 252522 129512
rect 252006 128616 252062 128625
rect 252006 128551 252062 128560
rect 252376 128308 252428 128314
rect 252376 128250 252428 128256
rect 252008 128172 252060 128178
rect 252008 128114 252060 128120
rect 252020 127265 252048 128114
rect 252388 127673 252416 128250
rect 252468 128240 252520 128246
rect 252466 128208 252468 128217
rect 252520 128208 252522 128217
rect 252466 128143 252522 128152
rect 252374 127664 252430 127673
rect 252374 127599 252430 127608
rect 252006 127256 252062 127265
rect 252006 127191 252062 127200
rect 252192 126948 252244 126954
rect 252192 126890 252244 126896
rect 251914 126304 251970 126313
rect 251914 126239 251970 126248
rect 252204 125769 252232 126890
rect 252468 126744 252520 126750
rect 252466 126712 252468 126721
rect 252520 126712 252522 126721
rect 252466 126647 252522 126656
rect 252190 125760 252246 125769
rect 252190 125695 252246 125704
rect 252192 125588 252244 125594
rect 252192 125530 252244 125536
rect 252100 124908 252152 124914
rect 252100 124850 252152 124856
rect 252008 123480 252060 123486
rect 252112 123457 252140 124850
rect 252204 124409 252232 125530
rect 252190 124400 252246 124409
rect 252190 124335 252246 124344
rect 252468 124160 252520 124166
rect 252468 124102 252520 124108
rect 252480 124001 252508 124102
rect 252466 123992 252522 124001
rect 252466 123927 252522 123936
rect 252008 123422 252060 123428
rect 252098 123448 252154 123457
rect 251916 121440 251968 121446
rect 251916 121382 251968 121388
rect 251928 120601 251956 121382
rect 251914 120592 251970 120601
rect 251914 120527 251970 120536
rect 251822 118824 251878 118833
rect 251822 118759 251878 118768
rect 251548 118448 251600 118454
rect 251548 118390 251600 118396
rect 251560 118289 251588 118390
rect 251546 118280 251602 118289
rect 251546 118215 251602 118224
rect 251824 117972 251876 117978
rect 251824 117914 251876 117920
rect 251548 116952 251600 116958
rect 251546 116920 251548 116929
rect 251600 116920 251602 116929
rect 251546 116855 251602 116864
rect 251640 115864 251692 115870
rect 251640 115806 251692 115812
rect 251652 115433 251680 115806
rect 251638 115424 251694 115433
rect 251638 115359 251694 115368
rect 251732 113416 251784 113422
rect 251732 113358 251784 113364
rect 251744 110809 251772 113358
rect 251730 110800 251786 110809
rect 251730 110735 251786 110744
rect 251456 110424 251508 110430
rect 251456 110366 251508 110372
rect 251468 109313 251496 110366
rect 251548 110356 251600 110362
rect 251548 110298 251600 110304
rect 251560 110265 251588 110298
rect 251546 110256 251602 110265
rect 251546 110191 251602 110200
rect 251454 109304 251510 109313
rect 251454 109239 251510 109248
rect 251836 109154 251864 117914
rect 251916 116612 251968 116618
rect 251916 116554 251968 116560
rect 251928 112713 251956 116554
rect 252020 113529 252048 123422
rect 252098 123383 252154 123392
rect 252284 122868 252336 122874
rect 252284 122810 252336 122816
rect 252100 121304 252152 121310
rect 252100 121246 252152 121252
rect 252112 120193 252140 121246
rect 252098 120184 252154 120193
rect 252098 120119 252154 120128
rect 252100 118652 252152 118658
rect 252100 118594 252152 118600
rect 252112 117337 252140 118594
rect 252098 117328 252154 117337
rect 252098 117263 252154 117272
rect 252296 115977 252324 122810
rect 252468 122800 252520 122806
rect 252468 122742 252520 122748
rect 252376 122732 252428 122738
rect 252376 122674 252428 122680
rect 252388 122097 252416 122674
rect 252480 122505 252508 122742
rect 252466 122496 252522 122505
rect 252466 122431 252522 122440
rect 252374 122088 252430 122097
rect 252374 122023 252430 122032
rect 252468 121576 252520 121582
rect 252466 121544 252468 121553
rect 252520 121544 252522 121553
rect 252466 121479 252522 121488
rect 252468 121372 252520 121378
rect 252468 121314 252520 121320
rect 252480 121145 252508 121314
rect 252466 121136 252522 121145
rect 252466 121071 252522 121080
rect 252376 120080 252428 120086
rect 252376 120022 252428 120028
rect 252388 119241 252416 120022
rect 252468 120012 252520 120018
rect 252468 119954 252520 119960
rect 252480 119649 252508 119954
rect 252466 119640 252522 119649
rect 252466 119575 252522 119584
rect 252374 119232 252430 119241
rect 252374 119167 252430 119176
rect 252468 118720 252520 118726
rect 252468 118662 252520 118668
rect 252480 117881 252508 118662
rect 252466 117872 252522 117881
rect 252466 117807 252522 117816
rect 252376 117292 252428 117298
rect 252376 117234 252428 117240
rect 252388 116385 252416 117234
rect 252374 116376 252430 116385
rect 252374 116311 252430 116320
rect 252282 115968 252338 115977
rect 252282 115903 252338 115912
rect 252376 115932 252428 115938
rect 252376 115874 252428 115880
rect 252388 115025 252416 115874
rect 252374 115016 252430 115025
rect 252374 114951 252430 114960
rect 252468 114504 252520 114510
rect 252466 114472 252468 114481
rect 252520 114472 252522 114481
rect 252466 114407 252522 114416
rect 252466 114064 252522 114073
rect 252466 113999 252522 114008
rect 252480 113762 252508 113999
rect 252468 113756 252520 113762
rect 252468 113698 252520 113704
rect 252006 113520 252062 113529
rect 252006 113455 252062 113464
rect 252100 113144 252152 113150
rect 252100 113086 252152 113092
rect 252190 113112 252246 113121
rect 251914 112704 251970 112713
rect 251914 112639 251970 112648
rect 252008 112464 252060 112470
rect 252008 112406 252060 112412
rect 251916 111104 251968 111110
rect 251916 111046 251968 111052
rect 251744 109126 251864 109154
rect 251180 108928 251232 108934
rect 251178 108896 251180 108905
rect 251232 108896 251234 108905
rect 251178 108831 251234 108840
rect 251548 107432 251600 107438
rect 251548 107374 251600 107380
rect 251560 106593 251588 107374
rect 251546 106584 251602 106593
rect 251546 106519 251602 106528
rect 251180 106208 251232 106214
rect 251180 106150 251232 106156
rect 251192 106049 251220 106150
rect 251178 106040 251234 106049
rect 251178 105975 251234 105984
rect 251640 105596 251692 105602
rect 251640 105538 251692 105544
rect 251652 98025 251680 105538
rect 251744 104689 251772 109126
rect 251824 108996 251876 109002
rect 251824 108938 251876 108944
rect 251836 108361 251864 108938
rect 251822 108352 251878 108361
rect 251822 108287 251878 108296
rect 251928 107953 251956 111046
rect 251914 107944 251970 107953
rect 251914 107879 251970 107888
rect 251730 104680 251786 104689
rect 251730 104615 251786 104624
rect 252020 103737 252048 112406
rect 252112 112169 252140 113086
rect 252190 113047 252192 113056
rect 252244 113047 252246 113056
rect 252192 113018 252244 113024
rect 252098 112160 252154 112169
rect 252098 112095 252154 112104
rect 252376 111784 252428 111790
rect 252374 111752 252376 111761
rect 252428 111752 252430 111761
rect 252374 111687 252430 111696
rect 252284 111240 252336 111246
rect 252284 111182 252336 111188
rect 252192 105664 252244 105670
rect 252192 105606 252244 105612
rect 252006 103728 252062 103737
rect 252006 103663 252062 103672
rect 252204 101425 252232 105606
rect 252296 105097 252324 111182
rect 252468 110288 252520 110294
rect 252468 110230 252520 110236
rect 252480 109857 252508 110230
rect 252466 109848 252522 109857
rect 252466 109783 252522 109792
rect 253216 108934 253244 149058
rect 253388 145580 253440 145586
rect 253388 145522 253440 145528
rect 253296 141432 253348 141438
rect 253296 141374 253348 141380
rect 253308 125390 253336 141374
rect 253296 125384 253348 125390
rect 253296 125326 253348 125332
rect 253296 114572 253348 114578
rect 253296 114514 253348 114520
rect 253204 108928 253256 108934
rect 253204 108870 253256 108876
rect 252560 108316 252612 108322
rect 252560 108258 252612 108264
rect 252376 107636 252428 107642
rect 252376 107578 252428 107584
rect 252388 107001 252416 107578
rect 252468 107568 252520 107574
rect 252466 107536 252468 107545
rect 252520 107536 252522 107545
rect 252466 107471 252522 107480
rect 252374 106992 252430 107001
rect 252374 106927 252430 106936
rect 252376 105732 252428 105738
rect 252376 105674 252428 105680
rect 252388 105641 252416 105674
rect 252374 105632 252430 105641
rect 252374 105567 252430 105576
rect 252282 105088 252338 105097
rect 252282 105023 252338 105032
rect 252468 104848 252520 104854
rect 252468 104790 252520 104796
rect 252284 104168 252336 104174
rect 252480 104145 252508 104790
rect 252284 104110 252336 104116
rect 252466 104136 252522 104145
rect 252296 102785 252324 104110
rect 252466 104071 252522 104080
rect 252376 103488 252428 103494
rect 252376 103430 252428 103436
rect 252282 102776 252338 102785
rect 252282 102711 252338 102720
rect 252388 102241 252416 103430
rect 252468 103420 252520 103426
rect 252468 103362 252520 103368
rect 252480 103193 252508 103362
rect 252466 103184 252522 103193
rect 252466 103119 252522 103128
rect 252374 102232 252430 102241
rect 252374 102167 252430 102176
rect 252468 102128 252520 102134
rect 252468 102070 252520 102076
rect 252190 101416 252246 101425
rect 252190 101351 252246 101360
rect 252008 101244 252060 101250
rect 252008 101186 252060 101192
rect 252020 100473 252048 101186
rect 252480 100881 252508 102070
rect 252466 100872 252522 100881
rect 252466 100807 252522 100816
rect 252100 100700 252152 100706
rect 252100 100642 252152 100648
rect 252006 100464 252062 100473
rect 252006 100399 252062 100408
rect 252112 99521 252140 100642
rect 252468 100632 252520 100638
rect 252468 100574 252520 100580
rect 252480 99929 252508 100574
rect 252466 99920 252522 99929
rect 252466 99855 252522 99864
rect 252098 99512 252154 99521
rect 252098 99447 252154 99456
rect 252468 99340 252520 99346
rect 252468 99282 252520 99288
rect 252376 99272 252428 99278
rect 252376 99214 252428 99220
rect 252388 98569 252416 99214
rect 252480 98977 252508 99282
rect 252466 98968 252522 98977
rect 252466 98903 252522 98912
rect 252374 98560 252430 98569
rect 252374 98495 252430 98504
rect 252468 98184 252520 98190
rect 252468 98126 252520 98132
rect 251638 98016 251694 98025
rect 251638 97951 251694 97960
rect 252480 97617 252508 98126
rect 252466 97608 252522 97617
rect 252466 97543 252522 97552
rect 251178 96656 251234 96665
rect 251178 96591 251234 96600
rect 250628 93152 250680 93158
rect 250628 93094 250680 93100
rect 250536 26920 250588 26926
rect 250536 26862 250588 26868
rect 249064 20052 249116 20058
rect 249064 19994 249116 20000
rect 248420 17264 248472 17270
rect 248420 17206 248472 17212
rect 247684 3460 247736 3466
rect 247684 3402 247736 3408
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248432 354 248460 17206
rect 251192 11014 251220 96591
rect 251270 96248 251326 96257
rect 251270 96183 251326 96192
rect 251284 86358 251312 96183
rect 251824 95260 251876 95266
rect 251824 95202 251876 95208
rect 251272 86352 251324 86358
rect 251272 86294 251324 86300
rect 251272 82136 251324 82142
rect 251272 82078 251324 82084
rect 251180 11008 251232 11014
rect 251180 10950 251232 10956
rect 251284 6914 251312 82078
rect 251836 33794 251864 95202
rect 251824 33788 251876 33794
rect 251824 33730 251876 33736
rect 252572 16574 252600 108258
rect 253204 96756 253256 96762
rect 253204 96698 253256 96704
rect 253216 29646 253244 96698
rect 253308 53174 253336 114514
rect 253400 106214 253428 145522
rect 253492 113422 253520 151778
rect 254136 150414 254164 192510
rect 254860 160744 254912 160750
rect 254860 160686 254912 160692
rect 254676 155984 254728 155990
rect 254676 155926 254728 155932
rect 254584 150476 254636 150482
rect 254584 150418 254636 150424
rect 254124 150408 254176 150414
rect 254124 150350 254176 150356
rect 253480 113416 253532 113422
rect 253480 113358 253532 113364
rect 254596 110430 254624 150418
rect 254688 115870 254716 155926
rect 254768 147688 254820 147694
rect 254768 147630 254820 147636
rect 254676 115864 254728 115870
rect 254676 115806 254728 115812
rect 254584 110424 254636 110430
rect 254584 110366 254636 110372
rect 254780 107438 254808 147630
rect 254872 132190 254900 160686
rect 255332 155922 255360 216106
rect 255976 213926 256004 233922
rect 256712 222970 256740 240094
rect 257344 224392 257396 224398
rect 257344 224334 257396 224340
rect 256700 222964 256752 222970
rect 256700 222906 256752 222912
rect 255964 213920 256016 213926
rect 255964 213862 256016 213868
rect 255504 191276 255556 191282
rect 255504 191218 255556 191224
rect 255412 176044 255464 176050
rect 255412 175986 255464 175992
rect 255320 155916 255372 155922
rect 255320 155858 255372 155864
rect 255424 148918 255452 175986
rect 255516 170950 255544 191218
rect 257356 189786 257384 224334
rect 258092 215082 258120 240094
rect 260104 235272 260156 235278
rect 260104 235214 260156 235220
rect 258080 215076 258132 215082
rect 258080 215018 258132 215024
rect 258724 213920 258776 213926
rect 258724 213862 258776 213868
rect 258172 209228 258224 209234
rect 258172 209170 258224 209176
rect 257344 189780 257396 189786
rect 257344 189722 257396 189728
rect 258080 188556 258132 188562
rect 258080 188498 258132 188504
rect 256700 187196 256752 187202
rect 256700 187138 256752 187144
rect 255596 185904 255648 185910
rect 255596 185846 255648 185852
rect 255504 170944 255556 170950
rect 255504 170886 255556 170892
rect 255608 168366 255636 185846
rect 256712 173738 256740 187138
rect 256792 184340 256844 184346
rect 256792 184282 256844 184288
rect 256700 173732 256752 173738
rect 256700 173674 256752 173680
rect 255596 168360 255648 168366
rect 255596 168302 255648 168308
rect 256804 158710 256832 184282
rect 256884 178968 256936 178974
rect 256884 178910 256936 178916
rect 256896 166802 256924 178910
rect 256976 177608 257028 177614
rect 256976 177550 257028 177556
rect 256884 166796 256936 166802
rect 256884 166738 256936 166744
rect 256792 158704 256844 158710
rect 256792 158646 256844 158652
rect 255964 153264 256016 153270
rect 255964 153206 256016 153212
rect 255412 148912 255464 148918
rect 255412 148854 255464 148860
rect 254860 132184 254912 132190
rect 254860 132126 254912 132132
rect 255976 113082 256004 153206
rect 256148 146328 256200 146334
rect 256148 146270 256200 146276
rect 256056 142316 256108 142322
rect 256056 142258 256108 142264
rect 255964 113076 256016 113082
rect 255964 113018 256016 113024
rect 255964 107908 256016 107914
rect 255964 107850 256016 107856
rect 254768 107432 254820 107438
rect 254768 107374 254820 107380
rect 253388 106208 253440 106214
rect 253388 106150 253440 106156
rect 254584 100972 254636 100978
rect 254584 100914 254636 100920
rect 253296 53168 253348 53174
rect 253296 53110 253348 53116
rect 253204 29640 253256 29646
rect 253204 29582 253256 29588
rect 254596 25566 254624 100914
rect 254584 25560 254636 25566
rect 254584 25502 254636 25508
rect 254584 24336 254636 24342
rect 254584 24278 254636 24284
rect 252572 16546 253520 16574
rect 252376 11960 252428 11966
rect 252376 11902 252428 11908
rect 251192 6886 251312 6914
rect 249984 3256 250036 3262
rect 249984 3198 250036 3204
rect 249996 480 250024 3198
rect 251192 480 251220 6886
rect 252388 480 252416 11902
rect 253492 480 253520 16546
rect 254596 3602 254624 24278
rect 255976 6186 256004 107850
rect 256068 101250 256096 142258
rect 256160 105738 256188 146270
rect 256240 145648 256292 145654
rect 256240 145590 256292 145596
rect 256252 111790 256280 145590
rect 256988 145518 257016 177550
rect 257436 164892 257488 164898
rect 257436 164834 257488 164840
rect 257344 157412 257396 157418
rect 257344 157354 257396 157360
rect 256976 145512 257028 145518
rect 256976 145454 257028 145460
rect 256698 138680 256754 138689
rect 256698 138615 256754 138624
rect 256240 111784 256292 111790
rect 256240 111726 256292 111732
rect 256608 111172 256660 111178
rect 256608 111114 256660 111120
rect 256148 105732 256200 105738
rect 256148 105674 256200 105680
rect 256056 101244 256108 101250
rect 256056 101186 256108 101192
rect 256056 90364 256108 90370
rect 256056 90306 256108 90312
rect 255964 6180 256016 6186
rect 255964 6122 256016 6128
rect 254584 3596 254636 3602
rect 254584 3538 254636 3544
rect 255870 3496 255926 3505
rect 254676 3460 254728 3466
rect 255870 3431 255926 3440
rect 254676 3402 254728 3408
rect 254688 480 254716 3402
rect 255884 480 255912 3431
rect 256068 3262 256096 90306
rect 256620 3466 256648 111114
rect 256608 3460 256660 3466
rect 256608 3402 256660 3408
rect 256056 3256 256108 3262
rect 256056 3198 256108 3204
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 256712 354 256740 138615
rect 257356 118454 257384 157354
rect 257448 126750 257476 164834
rect 257526 148336 257582 148345
rect 257526 148271 257582 148280
rect 257436 126744 257488 126750
rect 257436 126686 257488 126692
rect 257344 118448 257396 118454
rect 257344 118390 257396 118396
rect 257540 116958 257568 148271
rect 258092 146130 258120 188498
rect 258184 171562 258212 209170
rect 258264 200864 258316 200870
rect 258264 200806 258316 200812
rect 258172 171556 258224 171562
rect 258172 171498 258224 171504
rect 258276 167278 258304 200806
rect 258736 188562 258764 213862
rect 260116 211818 260144 235214
rect 259460 211812 259512 211818
rect 259460 211754 259512 211760
rect 260104 211812 260156 211818
rect 260104 211754 260156 211760
rect 258724 188556 258776 188562
rect 258724 188498 258776 188504
rect 258356 183184 258408 183190
rect 258356 183126 258408 183132
rect 258264 167272 258316 167278
rect 258264 167214 258316 167220
rect 258368 166530 258396 183126
rect 258356 166524 258408 166530
rect 258356 166466 258408 166472
rect 259092 165640 259144 165646
rect 259092 165582 259144 165588
rect 258724 156052 258776 156058
rect 258724 155994 258776 156000
rect 258080 146124 258132 146130
rect 258080 146066 258132 146072
rect 258736 122874 258764 155994
rect 258908 152516 258960 152522
rect 258908 152458 258960 152464
rect 258816 136740 258868 136746
rect 258816 136682 258868 136688
rect 258724 122868 258776 122874
rect 258724 122810 258776 122816
rect 257528 116952 257580 116958
rect 257528 116894 257580 116900
rect 258724 99408 258776 99414
rect 258724 99350 258776 99356
rect 258080 83564 258132 83570
rect 258080 83506 258132 83512
rect 258092 16574 258120 83506
rect 258092 16546 258304 16574
rect 258276 480 258304 16546
rect 258736 15910 258764 99350
rect 258828 65618 258856 136682
rect 258920 121310 258948 152458
rect 258998 144120 259054 144129
rect 258998 144055 259054 144064
rect 258908 121304 258960 121310
rect 258908 121246 258960 121252
rect 259012 113762 259040 144055
rect 259104 137154 259132 165582
rect 259472 148646 259500 211754
rect 260852 206446 260880 240094
rect 262784 238882 262812 240094
rect 265682 239850 265710 240108
rect 265636 239822 265710 239850
rect 266372 240094 267628 240122
rect 269560 240094 269804 240122
rect 262220 238876 262272 238882
rect 262220 238818 262272 238824
rect 262772 238876 262824 238882
rect 262772 238818 262824 238824
rect 260840 206440 260892 206446
rect 260840 206382 260892 206388
rect 259552 205012 259604 205018
rect 259552 204954 259604 204960
rect 259564 169862 259592 204954
rect 260932 198076 260984 198082
rect 260932 198018 260984 198024
rect 260840 191344 260892 191350
rect 260840 191286 260892 191292
rect 259644 175976 259696 175982
rect 259644 175918 259696 175924
rect 259552 169856 259604 169862
rect 259552 169798 259604 169804
rect 259656 159390 259684 175918
rect 260380 169788 260432 169794
rect 260380 169730 260432 169736
rect 260104 160812 260156 160818
rect 260104 160754 260156 160760
rect 259644 159384 259696 159390
rect 259644 159326 259696 159332
rect 259460 148640 259512 148646
rect 259460 148582 259512 148588
rect 259092 137148 259144 137154
rect 259092 137090 259144 137096
rect 260116 121582 260144 160754
rect 260196 157480 260248 157486
rect 260196 157422 260248 157428
rect 260104 121576 260156 121582
rect 260104 121518 260156 121524
rect 260208 118726 260236 157422
rect 260392 139874 260420 169730
rect 260852 144838 260880 191286
rect 260944 161430 260972 198018
rect 261024 189984 261076 189990
rect 261024 189926 261076 189932
rect 261036 167006 261064 189926
rect 261668 171148 261720 171154
rect 261668 171090 261720 171096
rect 261024 167000 261076 167006
rect 261024 166942 261076 166948
rect 260932 161424 260984 161430
rect 260932 161366 260984 161372
rect 261484 154624 261536 154630
rect 261484 154566 261536 154572
rect 260840 144832 260892 144838
rect 260840 144774 260892 144780
rect 260380 139868 260432 139874
rect 260380 139810 260432 139816
rect 260288 139460 260340 139466
rect 260288 139402 260340 139408
rect 260196 118720 260248 118726
rect 260196 118662 260248 118668
rect 259000 113756 259052 113762
rect 259000 113698 259052 113704
rect 260104 113212 260156 113218
rect 260104 113154 260156 113160
rect 258816 65612 258868 65618
rect 258816 65554 258868 65560
rect 259552 32496 259604 32502
rect 259552 32438 259604 32444
rect 259564 16574 259592 32438
rect 260116 28286 260144 113154
rect 260196 100836 260248 100842
rect 260196 100778 260248 100784
rect 260208 46238 260236 100778
rect 260300 98190 260328 139402
rect 260380 124228 260432 124234
rect 260380 124170 260432 124176
rect 260288 98184 260340 98190
rect 260288 98126 260340 98132
rect 260392 89214 260420 124170
rect 261496 114510 261524 154566
rect 261576 138100 261628 138106
rect 261576 138042 261628 138048
rect 261484 114504 261536 114510
rect 261484 114446 261536 114452
rect 261484 106344 261536 106350
rect 261484 106286 261536 106292
rect 260380 89208 260432 89214
rect 260380 89150 260432 89156
rect 260196 46232 260248 46238
rect 260196 46174 260248 46180
rect 260104 28280 260156 28286
rect 260104 28222 260156 28228
rect 261496 18630 261524 106286
rect 261588 51882 261616 138042
rect 261680 133754 261708 171090
rect 262232 162081 262260 238818
rect 265636 234462 265664 239822
rect 264980 234456 265032 234462
rect 264980 234398 265032 234404
rect 265624 234456 265676 234462
rect 265624 234398 265676 234404
rect 264992 233209 265020 234398
rect 264978 233200 265034 233209
rect 264978 233135 265034 233144
rect 264336 229764 264388 229770
rect 264336 229706 264388 229712
rect 264244 215076 264296 215082
rect 264244 215018 264296 215024
rect 263600 195492 263652 195498
rect 263600 195434 263652 195440
rect 262404 194132 262456 194138
rect 262404 194074 262456 194080
rect 262312 177540 262364 177546
rect 262312 177482 262364 177488
rect 262218 162072 262274 162081
rect 262218 162007 262274 162016
rect 261760 158772 261812 158778
rect 261760 158714 261812 158720
rect 261668 133748 261720 133754
rect 261668 133690 261720 133696
rect 261772 127634 261800 158714
rect 262324 146198 262352 177482
rect 262416 169726 262444 194074
rect 262496 180328 262548 180334
rect 262496 180270 262548 180276
rect 262404 169720 262456 169726
rect 262404 169662 262456 169668
rect 262508 165442 262536 180270
rect 262864 168428 262916 168434
rect 262864 168370 262916 168376
rect 262496 165436 262548 165442
rect 262496 165378 262548 165384
rect 262312 146192 262364 146198
rect 262312 146134 262364 146140
rect 262876 129606 262904 168370
rect 263612 165510 263640 195434
rect 263692 188624 263744 188630
rect 263692 188566 263744 188572
rect 263600 165504 263652 165510
rect 263600 165446 263652 165452
rect 263704 162858 263732 188566
rect 263692 162852 263744 162858
rect 263692 162794 263744 162800
rect 262956 162172 263008 162178
rect 262956 162114 263008 162120
rect 262864 129600 262916 129606
rect 262864 129542 262916 129548
rect 261760 127628 261812 127634
rect 261760 127570 261812 127576
rect 261760 119400 261812 119406
rect 261760 119342 261812 119348
rect 261772 99278 261800 119342
rect 262864 116000 262916 116006
rect 262864 115942 262916 115948
rect 261760 99272 261812 99278
rect 261760 99214 261812 99220
rect 261668 98048 261720 98054
rect 261668 97990 261720 97996
rect 261576 51876 261628 51882
rect 261576 51818 261628 51824
rect 261576 33992 261628 33998
rect 261576 33934 261628 33940
rect 261484 18624 261536 18630
rect 261484 18566 261536 18572
rect 259564 16546 260696 16574
rect 258724 15904 258776 15910
rect 258724 15846 258776 15852
rect 259460 3528 259512 3534
rect 259460 3470 259512 3476
rect 259472 480 259500 3470
rect 260668 480 260696 16546
rect 261588 4146 261616 33934
rect 261680 21418 261708 97990
rect 261668 21412 261720 21418
rect 261668 21354 261720 21360
rect 262496 11892 262548 11898
rect 262496 11834 262548 11840
rect 261576 4140 261628 4146
rect 261576 4082 261628 4088
rect 261760 3596 261812 3602
rect 261760 3538 261812 3544
rect 261772 480 261800 3538
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 11834
rect 262876 4826 262904 115942
rect 262968 99346 262996 162114
rect 263048 153332 263100 153338
rect 263048 153274 263100 153280
rect 263060 116618 263088 153274
rect 263048 116612 263100 116618
rect 263048 116554 263100 116560
rect 262956 99340 263008 99346
rect 262956 99282 263008 99288
rect 262864 4820 262916 4826
rect 262864 4762 262916 4768
rect 264150 3360 264206 3369
rect 264256 3330 264284 215018
rect 264348 191282 264376 229706
rect 264980 198144 265032 198150
rect 264980 198086 265032 198092
rect 264336 191276 264388 191282
rect 264336 191218 264388 191224
rect 264428 173936 264480 173942
rect 264428 173878 264480 173884
rect 264336 158840 264388 158846
rect 264336 158782 264388 158788
rect 264348 120018 264376 158782
rect 264440 136474 264468 173878
rect 264992 144906 265020 198086
rect 265072 181756 265124 181762
rect 265072 181698 265124 181704
rect 265084 157282 265112 181698
rect 265624 171216 265676 171222
rect 265624 171158 265676 171164
rect 265072 157276 265124 157282
rect 265072 157218 265124 157224
rect 265072 145716 265124 145722
rect 265072 145658 265124 145664
rect 264980 144900 265032 144906
rect 264980 144842 265032 144848
rect 264428 136468 264480 136474
rect 264428 136410 264480 136416
rect 264336 120012 264388 120018
rect 264336 119954 264388 119960
rect 264336 113280 264388 113286
rect 264336 113222 264388 113228
rect 264348 50386 264376 113222
rect 264336 50380 264388 50386
rect 264336 50322 264388 50328
rect 264150 3295 264206 3304
rect 264244 3324 264296 3330
rect 264164 480 264192 3295
rect 264244 3266 264296 3272
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 265084 354 265112 145658
rect 265636 132462 265664 171158
rect 265716 162920 265768 162926
rect 265716 162862 265768 162868
rect 265624 132456 265676 132462
rect 265624 132398 265676 132404
rect 265728 124914 265756 162862
rect 265716 124908 265768 124914
rect 265716 124850 265768 124856
rect 265624 124296 265676 124302
rect 265624 124238 265676 124244
rect 265636 13122 265664 124238
rect 266372 90370 266400 240094
rect 269776 238513 269804 240094
rect 271156 240094 271492 240122
rect 273732 240094 274068 240122
rect 276000 240094 276336 240122
rect 269762 238504 269818 238513
rect 269762 238439 269818 238448
rect 269776 231713 269804 238439
rect 271156 233034 271184 240094
rect 273732 238921 273760 240094
rect 273718 238912 273774 238921
rect 273718 238847 273774 238856
rect 276308 235754 276336 240094
rect 277412 240094 277932 240122
rect 276296 235748 276348 235754
rect 276296 235690 276348 235696
rect 276664 235748 276716 235754
rect 276664 235690 276716 235696
rect 271144 233028 271196 233034
rect 271144 232970 271196 232976
rect 274640 232620 274692 232626
rect 274640 232562 274692 232568
rect 269762 231704 269818 231713
rect 269762 231639 269818 231648
rect 267740 220380 267792 220386
rect 267740 220322 267792 220328
rect 266452 217592 266504 217598
rect 266452 217534 266504 217540
rect 266464 149054 266492 217534
rect 266544 188488 266596 188494
rect 266544 188430 266596 188436
rect 266556 165578 266584 188430
rect 267096 169856 267148 169862
rect 267096 169798 267148 169804
rect 266544 165572 266596 165578
rect 266544 165514 266596 165520
rect 266452 149048 266504 149054
rect 266452 148990 266504 148996
rect 267004 131164 267056 131170
rect 267004 131106 267056 131112
rect 266360 90364 266412 90370
rect 266360 90306 266412 90312
rect 267016 57254 267044 131106
rect 267108 131034 267136 169798
rect 267752 151638 267780 220322
rect 273352 219020 273404 219026
rect 273352 218962 273404 218968
rect 270500 217524 270552 217530
rect 270500 217466 270552 217472
rect 269120 199572 269172 199578
rect 269120 199514 269172 199520
rect 267832 195560 267884 195566
rect 267832 195502 267884 195508
rect 267740 151632 267792 151638
rect 267740 151574 267792 151580
rect 267844 137834 267872 195502
rect 268384 190052 268436 190058
rect 268384 189994 268436 190000
rect 267832 137828 267884 137834
rect 267832 137770 267884 137776
rect 267096 131028 267148 131034
rect 267096 130970 267148 130976
rect 267004 57248 267056 57254
rect 267004 57190 267056 57196
rect 265624 13116 265676 13122
rect 265624 13058 265676 13064
rect 266544 6384 266596 6390
rect 266544 6326 266596 6332
rect 266556 480 266584 6326
rect 267740 3732 267792 3738
rect 267740 3674 267792 3680
rect 267752 480 267780 3674
rect 268396 3534 268424 189994
rect 269132 155786 269160 199514
rect 269212 189916 269264 189922
rect 269212 189858 269264 189864
rect 269120 155780 269172 155786
rect 269120 155722 269172 155728
rect 269224 153066 269252 189858
rect 269856 172576 269908 172582
rect 269856 172518 269908 172524
rect 269212 153060 269264 153066
rect 269212 153002 269264 153008
rect 268568 150544 268620 150550
rect 268568 150486 268620 150492
rect 268476 129804 268528 129810
rect 268476 129746 268528 129752
rect 268488 24138 268516 129746
rect 268580 110362 268608 150486
rect 269764 147756 269816 147762
rect 269764 147698 269816 147704
rect 268568 110356 268620 110362
rect 268568 110298 268620 110304
rect 269776 107574 269804 147698
rect 269868 135182 269896 172518
rect 269948 165708 270000 165714
rect 269948 165650 270000 165656
rect 269856 135176 269908 135182
rect 269856 135118 269908 135124
rect 269960 128178 269988 165650
rect 270512 164218 270540 217466
rect 273260 211948 273312 211954
rect 273260 211890 273312 211896
rect 271880 210452 271932 210458
rect 271880 210394 271932 210400
rect 270592 193928 270644 193934
rect 270592 193870 270644 193876
rect 270500 164212 270552 164218
rect 270500 164154 270552 164160
rect 270604 154562 270632 193870
rect 271236 172644 271288 172650
rect 271236 172586 271288 172592
rect 270592 154556 270644 154562
rect 270592 154498 270644 154504
rect 271144 139528 271196 139534
rect 271144 139470 271196 139476
rect 270040 133952 270092 133958
rect 270040 133894 270092 133900
rect 269948 128172 270000 128178
rect 269948 128114 270000 128120
rect 269856 127016 269908 127022
rect 269856 126958 269908 126964
rect 269764 107568 269816 107574
rect 269764 107510 269816 107516
rect 269764 98116 269816 98122
rect 269764 98058 269816 98064
rect 268476 24132 268528 24138
rect 268476 24074 268528 24080
rect 269776 7614 269804 98058
rect 269868 37942 269896 126958
rect 269948 80708 270000 80714
rect 269948 80650 270000 80656
rect 269856 37936 269908 37942
rect 269856 37878 269908 37884
rect 269764 7608 269816 7614
rect 269764 7550 269816 7556
rect 268844 4140 268896 4146
rect 268844 4082 268896 4088
rect 268384 3528 268436 3534
rect 268384 3470 268436 3476
rect 268856 480 268884 4082
rect 269960 3058 269988 80650
rect 270052 75274 270080 133894
rect 270040 75268 270092 75274
rect 270040 75210 270092 75216
rect 271156 40730 271184 139470
rect 271248 133822 271276 172586
rect 271328 164960 271380 164966
rect 271328 164902 271380 164908
rect 271236 133816 271288 133822
rect 271236 133758 271288 133764
rect 271340 131102 271368 164902
rect 271420 133204 271472 133210
rect 271420 133146 271472 133152
rect 271328 131096 271380 131102
rect 271328 131038 271380 131044
rect 271328 125656 271380 125662
rect 271328 125598 271380 125604
rect 271236 102196 271288 102202
rect 271236 102138 271288 102144
rect 271144 40724 271196 40730
rect 271144 40666 271196 40672
rect 271248 22778 271276 102138
rect 271340 61402 271368 125598
rect 271432 103426 271460 133146
rect 271420 103420 271472 103426
rect 271420 103362 271472 103368
rect 271328 61396 271380 61402
rect 271328 61338 271380 61344
rect 271236 22772 271288 22778
rect 271236 22714 271288 22720
rect 271892 16574 271920 210394
rect 271972 207664 272024 207670
rect 271972 207606 272024 207612
rect 271984 153134 272012 207606
rect 272064 192636 272116 192642
rect 272064 192578 272116 192584
rect 272076 157350 272104 192578
rect 272524 162988 272576 162994
rect 272524 162930 272576 162936
rect 272064 157344 272116 157350
rect 272064 157286 272116 157292
rect 271972 153128 272024 153134
rect 271972 153070 272024 153076
rect 272536 124166 272564 162930
rect 272616 142248 272668 142254
rect 272616 142190 272668 142196
rect 272524 124160 272576 124166
rect 272524 124102 272576 124108
rect 272524 109064 272576 109070
rect 272524 109006 272576 109012
rect 272536 55894 272564 109006
rect 272628 102134 272656 142190
rect 273272 137902 273300 211890
rect 273364 150346 273392 218962
rect 273444 203652 273496 203658
rect 273444 203594 273496 203600
rect 273352 150340 273404 150346
rect 273352 150282 273404 150288
rect 273456 146266 273484 203594
rect 273904 168496 273956 168502
rect 273904 168438 273956 168444
rect 273916 146946 273944 168438
rect 273904 146940 273956 146946
rect 273904 146882 273956 146888
rect 274180 146396 274232 146402
rect 274180 146338 274232 146344
rect 273444 146260 273496 146266
rect 273444 146202 273496 146208
rect 274088 143608 274140 143614
rect 274088 143550 274140 143556
rect 273260 137896 273312 137902
rect 273260 137838 273312 137844
rect 273904 129872 273956 129878
rect 273904 129814 273956 129820
rect 272616 102128 272668 102134
rect 272616 102070 272668 102076
rect 272524 55888 272576 55894
rect 272524 55830 272576 55836
rect 271892 16546 272472 16574
rect 271236 3460 271288 3466
rect 271236 3402 271288 3408
rect 270040 3324 270092 3330
rect 270040 3266 270092 3272
rect 269948 3052 270000 3058
rect 269948 2994 270000 3000
rect 270052 480 270080 3266
rect 271248 480 271276 3402
rect 272444 480 272472 16546
rect 273260 16040 273312 16046
rect 273260 15982 273312 15988
rect 265318 354 265430 480
rect 265084 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273272 354 273300 15982
rect 273916 9042 273944 129814
rect 273996 120148 274048 120154
rect 273996 120090 274048 120096
rect 274008 14550 274036 120090
rect 274100 103494 274128 143550
rect 274192 111246 274220 146338
rect 274180 111240 274232 111246
rect 274180 111182 274232 111188
rect 274088 103488 274140 103494
rect 274088 103430 274140 103436
rect 274180 102264 274232 102270
rect 274180 102206 274232 102212
rect 274192 73846 274220 102206
rect 274180 73840 274232 73846
rect 274180 73782 274232 73788
rect 274652 16574 274680 232562
rect 276676 227633 276704 235690
rect 277412 229090 277440 240094
rect 279988 238882 280016 240366
rect 281552 240094 282440 240122
rect 278872 238876 278924 238882
rect 278872 238818 278924 238824
rect 279976 238876 280028 238882
rect 279976 238818 280028 238824
rect 278780 232688 278832 232694
rect 278780 232630 278832 232636
rect 277400 229084 277452 229090
rect 277400 229026 277452 229032
rect 276662 227624 276718 227633
rect 276662 227559 276718 227568
rect 278044 222964 278096 222970
rect 278044 222906 278096 222912
rect 274732 217456 274784 217462
rect 274732 217398 274784 217404
rect 274744 150278 274772 217398
rect 276020 214736 276072 214742
rect 276020 214678 276072 214684
rect 274824 211880 274876 211886
rect 274824 211822 274876 211828
rect 274836 151706 274864 211822
rect 275284 167068 275336 167074
rect 275284 167010 275336 167016
rect 274824 151700 274876 151706
rect 274824 151642 274876 151648
rect 274732 150272 274784 150278
rect 274732 150214 274784 150220
rect 275296 129674 275324 167010
rect 276032 151774 276060 214678
rect 277400 213376 277452 213382
rect 277400 213318 277452 213324
rect 276112 202156 276164 202162
rect 276112 202098 276164 202104
rect 276020 151768 276072 151774
rect 276020 151710 276072 151716
rect 276124 147558 276152 202098
rect 276848 160132 276900 160138
rect 276848 160074 276900 160080
rect 276112 147552 276164 147558
rect 276112 147494 276164 147500
rect 276756 146940 276808 146946
rect 276756 146882 276808 146888
rect 275284 129668 275336 129674
rect 275284 129610 275336 129616
rect 276664 128444 276716 128450
rect 276664 128386 276716 128392
rect 275376 128376 275428 128382
rect 275376 128318 275428 128324
rect 275284 122868 275336 122874
rect 275284 122810 275336 122816
rect 275296 29714 275324 122810
rect 275388 43518 275416 128318
rect 276112 106956 276164 106962
rect 276112 106898 276164 106904
rect 275376 43512 275428 43518
rect 275376 43454 275428 43460
rect 275284 29708 275336 29714
rect 275284 29650 275336 29656
rect 276124 16574 276152 106898
rect 276676 44878 276704 128386
rect 276768 107642 276796 146882
rect 276860 121378 276888 160074
rect 277412 147626 277440 213318
rect 277400 147620 277452 147626
rect 277400 147562 277452 147568
rect 276848 121372 276900 121378
rect 276848 121314 276900 121320
rect 276756 107636 276808 107642
rect 276756 107578 276808 107584
rect 276664 44872 276716 44878
rect 276664 44814 276716 44820
rect 274652 16546 274864 16574
rect 276124 16546 276704 16574
rect 273996 14544 274048 14550
rect 273996 14486 274048 14492
rect 273904 9036 273956 9042
rect 273904 8978 273956 8984
rect 274836 480 274864 16546
rect 276020 3052 276072 3058
rect 276020 2994 276072 3000
rect 276032 480 276060 2994
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276676 354 276704 16546
rect 278056 3738 278084 222906
rect 278228 167136 278280 167142
rect 278228 167078 278280 167084
rect 278240 128246 278268 167078
rect 278320 159384 278372 159390
rect 278320 159326 278372 159332
rect 278228 128240 278280 128246
rect 278228 128182 278280 128188
rect 278136 127084 278188 127090
rect 278136 127026 278188 127032
rect 278148 10334 278176 127026
rect 278332 126954 278360 159326
rect 278320 126948 278372 126954
rect 278320 126890 278372 126896
rect 278228 121508 278280 121514
rect 278228 121450 278280 121456
rect 278240 33862 278268 121450
rect 278320 103556 278372 103562
rect 278320 103498 278372 103504
rect 278332 91798 278360 103498
rect 278320 91792 278372 91798
rect 278320 91734 278372 91740
rect 278228 33856 278280 33862
rect 278228 33798 278280 33804
rect 278792 16574 278820 232630
rect 278884 224942 278912 238818
rect 280160 227180 280212 227186
rect 280160 227122 280212 227128
rect 278872 224936 278924 224942
rect 278872 224878 278924 224884
rect 278872 218884 278924 218890
rect 278872 218826 278924 218832
rect 278884 137970 278912 218826
rect 279424 208004 279476 208010
rect 279424 207946 279476 207952
rect 278872 137964 278924 137970
rect 278872 137906 278924 137912
rect 278792 16546 279096 16574
rect 278136 10328 278188 10334
rect 278136 10270 278188 10276
rect 278044 3732 278096 3738
rect 278044 3674 278096 3680
rect 278320 3528 278372 3534
rect 278320 3470 278372 3476
rect 278332 480 278360 3470
rect 277094 354 277206 480
rect 276676 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 279436 3466 279464 207946
rect 279608 161492 279660 161498
rect 279608 161434 279660 161440
rect 279516 127152 279568 127158
rect 279516 127094 279568 127100
rect 279528 36582 279556 127094
rect 279620 122738 279648 161434
rect 279608 122732 279660 122738
rect 279608 122674 279660 122680
rect 279516 36576 279568 36582
rect 279516 36518 279568 36524
rect 280172 16574 280200 227122
rect 281552 207670 281580 240094
rect 284358 239850 284386 240108
rect 284312 239822 284386 239850
rect 285692 240094 286304 240122
rect 287072 240094 288236 240122
rect 289924 240094 290812 240122
rect 292592 240094 292744 240122
rect 283564 227112 283616 227118
rect 283564 227054 283616 227060
rect 282920 210656 282972 210662
rect 282920 210598 282972 210604
rect 281632 207868 281684 207874
rect 281632 207810 281684 207816
rect 281540 207664 281592 207670
rect 281540 207606 281592 207612
rect 281540 202428 281592 202434
rect 281540 202370 281592 202376
rect 280804 171284 280856 171290
rect 280804 171226 280856 171232
rect 280816 133890 280844 171226
rect 280988 140888 281040 140894
rect 280988 140830 281040 140836
rect 280896 136808 280948 136814
rect 280896 136750 280948 136756
rect 280804 133884 280856 133890
rect 280804 133826 280856 133832
rect 280804 120216 280856 120222
rect 280804 120158 280856 120164
rect 280816 19990 280844 120158
rect 280908 64258 280936 136750
rect 281000 100638 281028 140830
rect 281552 140758 281580 202370
rect 281644 153202 281672 207810
rect 282184 183048 282236 183054
rect 282184 182990 282236 182996
rect 281632 153196 281684 153202
rect 281632 153138 281684 153144
rect 281540 140752 281592 140758
rect 281540 140694 281592 140700
rect 280988 100632 281040 100638
rect 280988 100574 281040 100580
rect 280896 64252 280948 64258
rect 280896 64194 280948 64200
rect 280804 19984 280856 19990
rect 280804 19926 280856 19932
rect 280172 16546 280752 16574
rect 279424 3460 279476 3466
rect 279424 3402 279476 3408
rect 280724 480 280752 16546
rect 281908 3664 281960 3670
rect 281908 3606 281960 3612
rect 281920 480 281948 3606
rect 282196 3602 282224 182990
rect 282276 174004 282328 174010
rect 282276 173946 282328 173952
rect 282288 136542 282316 173946
rect 282460 145784 282512 145790
rect 282460 145726 282512 145732
rect 282276 136536 282328 136542
rect 282276 136478 282328 136484
rect 282368 135516 282420 135522
rect 282368 135458 282420 135464
rect 282276 132524 282328 132530
rect 282276 132466 282328 132472
rect 282288 60110 282316 132466
rect 282380 66978 282408 135458
rect 282472 111178 282500 145726
rect 282460 111172 282512 111178
rect 282460 111114 282512 111120
rect 282368 66972 282420 66978
rect 282368 66914 282420 66920
rect 282368 65680 282420 65686
rect 282368 65622 282420 65628
rect 282276 60104 282328 60110
rect 282276 60046 282328 60052
rect 282184 3596 282236 3602
rect 282184 3538 282236 3544
rect 282380 3534 282408 65622
rect 282932 16574 282960 210598
rect 283576 180198 283604 227054
rect 283564 180192 283616 180198
rect 283564 180134 283616 180140
rect 283564 168564 283616 168570
rect 283564 168506 283616 168512
rect 283576 129742 283604 168506
rect 283748 153400 283800 153406
rect 283748 153342 283800 153348
rect 283656 129940 283708 129946
rect 283656 129882 283708 129888
rect 283564 129736 283616 129742
rect 283564 129678 283616 129684
rect 283564 122936 283616 122942
rect 283564 122878 283616 122884
rect 282932 16546 283144 16574
rect 282368 3528 282420 3534
rect 282368 3470 282420 3476
rect 283116 480 283144 16546
rect 283576 11762 283604 122878
rect 283668 39438 283696 129882
rect 283760 123486 283788 153342
rect 283748 123480 283800 123486
rect 283748 123422 283800 123428
rect 283748 110492 283800 110498
rect 283748 110434 283800 110440
rect 283760 61470 283788 110434
rect 284312 83570 284340 239822
rect 285128 156120 285180 156126
rect 285128 156062 285180 156068
rect 284944 121576 284996 121582
rect 284944 121518 284996 121524
rect 284300 83564 284352 83570
rect 284300 83506 284352 83512
rect 283748 61464 283800 61470
rect 283748 61406 283800 61412
rect 283656 39432 283708 39438
rect 283656 39374 283708 39380
rect 284956 24206 284984 121518
rect 285140 117298 285168 156062
rect 285128 117292 285180 117298
rect 285128 117234 285180 117240
rect 285036 116068 285088 116074
rect 285036 116010 285088 116016
rect 285048 54534 285076 116010
rect 285036 54528 285088 54534
rect 285036 54470 285088 54476
rect 284944 24200 284996 24206
rect 284944 24142 284996 24148
rect 283564 11756 283616 11762
rect 283564 11698 283616 11704
rect 284300 3528 284352 3534
rect 285692 3482 285720 240094
rect 287072 231849 287100 240094
rect 287704 239420 287756 239426
rect 287704 239362 287756 239368
rect 287058 231840 287114 231849
rect 287058 231775 287114 231784
rect 287716 166297 287744 239362
rect 289820 233708 289872 233714
rect 289820 233650 289872 233656
rect 289084 206440 289136 206446
rect 289084 206382 289136 206388
rect 288072 174072 288124 174078
rect 288072 174014 288124 174020
rect 287702 166288 287758 166297
rect 287702 166223 287758 166232
rect 287796 164280 287848 164286
rect 287796 164222 287848 164228
rect 286324 139596 286376 139602
rect 286324 139538 286376 139544
rect 285770 80744 285826 80753
rect 285770 80679 285826 80688
rect 285784 16574 285812 80679
rect 286336 46306 286364 139538
rect 287808 125594 287836 164222
rect 287980 157548 288032 157554
rect 287980 157490 288032 157496
rect 287888 138168 287940 138174
rect 287888 138110 287940 138116
rect 287796 125588 287848 125594
rect 287796 125530 287848 125536
rect 287704 124364 287756 124370
rect 287704 124306 287756 124312
rect 286324 46300 286376 46306
rect 286324 46242 286376 46248
rect 285784 16546 286640 16574
rect 284300 3470 284352 3476
rect 284312 480 284340 3470
rect 285416 3454 285720 3482
rect 285416 480 285444 3454
rect 286612 480 286640 16546
rect 287716 7682 287744 124306
rect 287796 117360 287848 117366
rect 287796 117302 287848 117308
rect 287808 16574 287836 117302
rect 287900 57390 287928 138110
rect 287992 118658 288020 157490
rect 288084 136610 288112 174014
rect 288072 136604 288124 136610
rect 288072 136546 288124 136552
rect 287980 118652 288032 118658
rect 287980 118594 288032 118600
rect 287980 114640 288032 114646
rect 287980 114582 288032 114588
rect 287888 57384 287940 57390
rect 287888 57326 287940 57332
rect 287992 49026 288020 114582
rect 287980 49020 288032 49026
rect 287980 48962 288032 48968
rect 287808 16546 287928 16574
rect 287796 9104 287848 9110
rect 287796 9046 287848 9052
rect 287704 7676 287756 7682
rect 287704 7618 287756 7624
rect 287808 480 287836 9046
rect 287900 2106 287928 16546
rect 289096 3602 289124 206382
rect 289268 161560 289320 161566
rect 289268 161502 289320 161508
rect 289176 123004 289228 123010
rect 289176 122946 289228 122952
rect 289188 15978 289216 122946
rect 289280 122806 289308 161502
rect 289360 134020 289412 134026
rect 289360 133962 289412 133968
rect 289268 122800 289320 122806
rect 289268 122742 289320 122748
rect 289268 96824 289320 96830
rect 289268 96766 289320 96772
rect 289176 15972 289228 15978
rect 289176 15914 289228 15920
rect 289280 8974 289308 96766
rect 289372 72486 289400 133962
rect 289360 72480 289412 72486
rect 289360 72422 289412 72428
rect 289268 8968 289320 8974
rect 289268 8910 289320 8916
rect 288992 3596 289044 3602
rect 288992 3538 289044 3544
rect 289084 3596 289136 3602
rect 289084 3538 289136 3544
rect 287888 2100 287940 2106
rect 287888 2042 287940 2048
rect 289004 480 289032 3538
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 289832 354 289860 233650
rect 289924 230450 289952 240094
rect 292592 237454 292620 240094
rect 291844 237448 291896 237454
rect 291844 237390 291896 237396
rect 292580 237448 292632 237454
rect 292580 237390 292632 237396
rect 289912 230444 289964 230450
rect 289912 230386 289964 230392
rect 291200 203856 291252 203862
rect 291200 203798 291252 203804
rect 290464 163056 290516 163062
rect 290464 162998 290516 163004
rect 290476 135930 290504 162998
rect 290464 135924 290516 135930
rect 290464 135866 290516 135872
rect 290556 135380 290608 135386
rect 290556 135322 290608 135328
rect 290464 125724 290516 125730
rect 290464 125666 290516 125672
rect 290476 6254 290504 125666
rect 290568 68406 290596 135322
rect 290556 68400 290608 68406
rect 290556 68342 290608 68348
rect 291212 16574 291240 203798
rect 291856 108322 291884 237390
rect 291936 167204 291988 167210
rect 291936 167146 291988 167152
rect 291948 128314 291976 167146
rect 293052 145722 293080 287399
rect 293144 230382 293172 301271
rect 293222 259176 293278 259185
rect 293222 259111 293278 259120
rect 293236 232626 293264 259111
rect 293314 241904 293370 241913
rect 293314 241839 293370 241848
rect 293328 241097 293356 241839
rect 293314 241088 293370 241097
rect 293314 241023 293370 241032
rect 293224 232620 293276 232626
rect 293224 232562 293276 232568
rect 293132 230376 293184 230382
rect 293132 230318 293184 230324
rect 293040 145716 293092 145722
rect 293040 145658 293092 145664
rect 293408 144968 293460 144974
rect 293408 144910 293460 144916
rect 293224 132592 293276 132598
rect 293224 132534 293276 132540
rect 291936 128308 291988 128314
rect 291936 128250 291988 128256
rect 291936 121644 291988 121650
rect 291936 121586 291988 121592
rect 291844 108316 291896 108322
rect 291844 108258 291896 108264
rect 291844 99476 291896 99482
rect 291844 99418 291896 99424
rect 291856 47598 291884 99418
rect 291844 47592 291896 47598
rect 291844 47534 291896 47540
rect 291948 21486 291976 121586
rect 292028 107024 292080 107030
rect 292028 106966 292080 106972
rect 292040 100706 292068 106966
rect 292028 100700 292080 100706
rect 292028 100642 292080 100648
rect 293236 35222 293264 132534
rect 293316 111852 293368 111858
rect 293316 111794 293368 111800
rect 293224 35216 293276 35222
rect 293224 35158 293276 35164
rect 293328 31074 293356 111794
rect 293420 104854 293448 144910
rect 293500 105052 293552 105058
rect 293500 104994 293552 105000
rect 293408 104848 293460 104854
rect 293408 104790 293460 104796
rect 293512 71058 293540 104994
rect 293972 82142 294000 352271
rect 294064 327865 294092 354758
rect 294156 338745 294184 358770
rect 294236 356040 294288 356046
rect 294236 355982 294288 355988
rect 294142 338736 294198 338745
rect 294142 338671 294198 338680
rect 294050 327856 294106 327865
rect 294050 327791 294106 327800
rect 294050 325816 294106 325825
rect 294050 325751 294106 325760
rect 294064 210458 294092 325751
rect 294142 323096 294198 323105
rect 294142 323031 294198 323040
rect 294156 233714 294184 323031
rect 294248 303618 294276 355982
rect 295352 343602 295380 362986
rect 295432 362228 295484 362234
rect 295432 362170 295484 362176
rect 295340 343596 295392 343602
rect 295340 343538 295392 343544
rect 295338 343496 295394 343505
rect 295338 343431 295394 343440
rect 295352 342922 295380 343431
rect 295340 342916 295392 342922
rect 295340 342858 295392 342864
rect 295338 340776 295394 340785
rect 295338 340711 295394 340720
rect 295352 339522 295380 340711
rect 295340 339516 295392 339522
rect 295340 339458 295392 339464
rect 295444 334665 295472 362170
rect 295524 356176 295576 356182
rect 295524 356118 295576 356124
rect 295430 334656 295486 334665
rect 295430 334591 295486 334600
rect 295338 331936 295394 331945
rect 295338 331871 295394 331880
rect 294418 327856 294474 327865
rect 294418 327791 294474 327800
rect 294432 327146 294460 327791
rect 294420 327140 294472 327146
rect 294420 327082 294472 327088
rect 294236 303612 294288 303618
rect 294236 303554 294288 303560
rect 294248 303385 294276 303554
rect 294234 303376 294290 303385
rect 294234 303311 294290 303320
rect 295352 294658 295380 331871
rect 295444 306374 295472 334591
rect 295536 325694 295564 356118
rect 295628 354385 295656 368494
rect 296812 357740 296864 357746
rect 296812 357682 296864 357688
rect 295614 354376 295670 354385
rect 295614 354311 295670 354320
rect 296166 345536 296222 345545
rect 296166 345471 296222 345480
rect 296180 345098 296208 345471
rect 296168 345092 296220 345098
rect 296168 345034 296220 345040
rect 295616 343596 295668 343602
rect 295616 343538 295668 343544
rect 295628 336705 295656 343538
rect 295614 336696 295670 336705
rect 295614 336631 295670 336640
rect 295536 325666 295656 325694
rect 295522 321056 295578 321065
rect 295522 320991 295578 321000
rect 295536 320210 295564 320991
rect 295524 320204 295576 320210
rect 295524 320146 295576 320152
rect 295522 319016 295578 319025
rect 295522 318951 295578 318960
rect 295536 318850 295564 318951
rect 295524 318844 295576 318850
rect 295524 318786 295576 318792
rect 295628 316985 295656 325666
rect 295614 316976 295670 316985
rect 295614 316911 295670 316920
rect 295628 316742 295656 316911
rect 295616 316736 295668 316742
rect 295616 316678 295668 316684
rect 295524 314628 295576 314634
rect 295524 314570 295576 314576
rect 295536 314265 295564 314570
rect 295522 314256 295578 314265
rect 295522 314191 295578 314200
rect 295522 312216 295578 312225
rect 295522 312151 295578 312160
rect 295536 311914 295564 312151
rect 295524 311908 295576 311914
rect 295524 311850 295576 311856
rect 295522 310176 295578 310185
rect 295522 310111 295578 310120
rect 295536 309806 295564 310111
rect 295524 309800 295576 309806
rect 295524 309742 295576 309748
rect 295522 308136 295578 308145
rect 295522 308071 295578 308080
rect 295536 307834 295564 308071
rect 295524 307828 295576 307834
rect 295524 307770 295576 307776
rect 295444 306346 295564 306374
rect 295430 305416 295486 305425
rect 295430 305351 295486 305360
rect 295444 305046 295472 305351
rect 295432 305040 295484 305046
rect 295432 304982 295484 304988
rect 295430 296576 295486 296585
rect 295430 296511 295486 296520
rect 295444 295390 295472 296511
rect 295432 295384 295484 295390
rect 295432 295326 295484 295332
rect 295352 294630 295472 294658
rect 295338 294536 295394 294545
rect 295338 294471 295394 294480
rect 295352 294030 295380 294471
rect 295340 294024 295392 294030
rect 295340 293966 295392 293972
rect 295444 291938 295472 294630
rect 295352 291910 295472 291938
rect 294234 268016 294290 268025
rect 294234 267951 294290 267960
rect 294144 233708 294196 233714
rect 294144 233650 294196 233656
rect 294248 232694 294276 267951
rect 295352 250918 295380 291910
rect 295536 291802 295564 306346
rect 296626 299296 296682 299305
rect 296682 299254 296760 299282
rect 296626 299231 296682 299240
rect 295614 292496 295670 292505
rect 295614 292431 295670 292440
rect 295444 291774 295564 291802
rect 295340 250912 295392 250918
rect 295340 250854 295392 250860
rect 295338 243536 295394 243545
rect 295338 243471 295394 243480
rect 295352 242962 295380 243471
rect 295340 242956 295392 242962
rect 295340 242898 295392 242904
rect 295338 241496 295394 241505
rect 295338 241431 295394 241440
rect 294236 232688 294288 232694
rect 294236 232630 294288 232636
rect 294052 210452 294104 210458
rect 294052 210394 294104 210400
rect 294604 170400 294656 170406
rect 294604 170342 294656 170348
rect 294616 135250 294644 170342
rect 294604 135244 294656 135250
rect 294604 135186 294656 135192
rect 294696 134088 294748 134094
rect 294696 134030 294748 134036
rect 294604 118720 294656 118726
rect 294604 118662 294656 118668
rect 293960 82136 294012 82142
rect 293960 82078 294012 82084
rect 293500 71052 293552 71058
rect 293500 70994 293552 71000
rect 293316 31068 293368 31074
rect 293316 31010 293368 31016
rect 293960 28416 294012 28422
rect 293960 28358 294012 28364
rect 291936 21480 291988 21486
rect 291936 21422 291988 21428
rect 293972 16574 294000 28358
rect 294616 22846 294644 118662
rect 294708 73914 294736 134030
rect 295352 106962 295380 241431
rect 295444 231742 295472 291774
rect 295522 290456 295578 290465
rect 295522 290391 295578 290400
rect 295536 289882 295564 290391
rect 295524 289876 295576 289882
rect 295524 289818 295576 289824
rect 295524 285728 295576 285734
rect 295522 285696 295524 285705
rect 295576 285696 295578 285705
rect 295522 285631 295578 285640
rect 295522 283656 295578 283665
rect 295522 283591 295578 283600
rect 295536 282946 295564 283591
rect 295524 282940 295576 282946
rect 295524 282882 295576 282888
rect 295522 281616 295578 281625
rect 295522 281551 295524 281560
rect 295576 281551 295578 281560
rect 295524 281522 295576 281528
rect 295522 278896 295578 278905
rect 295522 278831 295578 278840
rect 295536 278798 295564 278831
rect 295524 278792 295576 278798
rect 295524 278734 295576 278740
rect 295628 277394 295656 292431
rect 295536 277366 295656 277394
rect 295536 253502 295564 277366
rect 295614 276856 295670 276865
rect 295614 276791 295670 276800
rect 295628 276078 295656 276791
rect 295616 276072 295668 276078
rect 295616 276014 295668 276020
rect 295706 274816 295762 274825
rect 295706 274751 295762 274760
rect 295614 272776 295670 272785
rect 295614 272711 295670 272720
rect 295628 271930 295656 272711
rect 295616 271924 295668 271930
rect 295616 271866 295668 271872
rect 295614 270056 295670 270065
rect 295614 269991 295670 270000
rect 295628 269142 295656 269991
rect 295616 269136 295668 269142
rect 295616 269078 295668 269084
rect 295614 265976 295670 265985
rect 295614 265911 295670 265920
rect 295628 264994 295656 265911
rect 295616 264988 295668 264994
rect 295616 264930 295668 264936
rect 295614 263936 295670 263945
rect 295614 263871 295670 263880
rect 295628 263634 295656 263871
rect 295616 263628 295668 263634
rect 295616 263570 295668 263576
rect 295614 261216 295670 261225
rect 295614 261151 295670 261160
rect 295628 260914 295656 261151
rect 295616 260908 295668 260914
rect 295616 260850 295668 260856
rect 295720 258074 295748 274751
rect 295628 258046 295748 258074
rect 295524 253496 295576 253502
rect 295524 253438 295576 253444
rect 295524 250912 295576 250918
rect 295524 250854 295576 250860
rect 295536 241466 295564 250854
rect 295524 241460 295576 241466
rect 295524 241402 295576 241408
rect 295628 235822 295656 258046
rect 295706 257136 295762 257145
rect 295706 257071 295708 257080
rect 295760 257071 295762 257080
rect 295708 257042 295760 257048
rect 295706 255096 295762 255105
rect 295706 255031 295762 255040
rect 295720 253978 295748 255031
rect 295708 253972 295760 253978
rect 295708 253914 295760 253920
rect 295708 253496 295760 253502
rect 295708 253438 295760 253444
rect 295720 240106 295748 253438
rect 296442 252376 296498 252385
rect 296442 252311 296498 252320
rect 296456 251258 296484 252311
rect 296444 251252 296496 251258
rect 296444 251194 296496 251200
rect 295798 250336 295854 250345
rect 295798 250271 295854 250280
rect 295812 249830 295840 250271
rect 295800 249824 295852 249830
rect 295800 249766 295852 249772
rect 296628 248396 296680 248402
rect 296628 248338 296680 248344
rect 296640 248305 296668 248338
rect 296626 248296 296682 248305
rect 296626 248231 296682 248240
rect 295708 240100 295760 240106
rect 295708 240042 295760 240048
rect 295616 235816 295668 235822
rect 295616 235758 295668 235764
rect 295432 231736 295484 231742
rect 295432 231678 295484 231684
rect 295984 154692 296036 154698
rect 295984 154634 296036 154640
rect 295996 115938 296024 154634
rect 296076 149728 296128 149734
rect 296076 149670 296128 149676
rect 296088 120086 296116 149670
rect 296076 120080 296128 120086
rect 296076 120022 296128 120028
rect 296168 118788 296220 118794
rect 296168 118730 296220 118736
rect 296076 116612 296128 116618
rect 296076 116554 296128 116560
rect 295984 115932 296036 115938
rect 295984 115874 296036 115880
rect 296088 113150 296116 116554
rect 296076 113144 296128 113150
rect 296076 113086 296128 113092
rect 295984 110560 296036 110566
rect 295984 110502 296036 110508
rect 295340 106956 295392 106962
rect 295340 106898 295392 106904
rect 294788 99544 294840 99550
rect 294788 99486 294840 99492
rect 294696 73908 294748 73914
rect 294696 73850 294748 73856
rect 294800 51746 294828 99486
rect 294788 51740 294840 51746
rect 294788 51682 294840 51688
rect 295996 42158 296024 110502
rect 296076 109132 296128 109138
rect 296076 109074 296128 109080
rect 296088 57322 296116 109074
rect 296180 76566 296208 118730
rect 296260 103624 296312 103630
rect 296260 103566 296312 103572
rect 296168 76560 296220 76566
rect 296168 76502 296220 76508
rect 296272 68338 296300 103566
rect 296732 89146 296760 299254
rect 296824 239426 296852 357682
rect 296902 246256 296958 246265
rect 296902 246191 296958 246200
rect 296916 245682 296944 246191
rect 296904 245676 296956 245682
rect 296904 245618 296956 245624
rect 296812 239420 296864 239426
rect 296812 239362 296864 239368
rect 296916 226302 296944 245618
rect 297376 238921 297404 683130
rect 298742 357504 298798 357513
rect 298742 357439 298798 357448
rect 298192 356108 298244 356114
rect 298192 356050 298244 356056
rect 297456 354952 297508 354958
rect 297456 354894 297508 354900
rect 297468 299470 297496 354894
rect 298098 354648 298154 354657
rect 298098 354583 298154 354592
rect 297456 299464 297508 299470
rect 297456 299406 297508 299412
rect 297362 238912 297418 238921
rect 297362 238847 297418 238856
rect 298112 228313 298140 354583
rect 298204 309806 298232 356050
rect 298192 309800 298244 309806
rect 298192 309742 298244 309748
rect 298192 257100 298244 257106
rect 298192 257042 298244 257048
rect 298204 234530 298232 257042
rect 298192 234524 298244 234530
rect 298192 234466 298244 234472
rect 298098 228304 298154 228313
rect 298098 228239 298154 228248
rect 296904 226296 296956 226302
rect 296904 226238 296956 226244
rect 297456 135448 297508 135454
rect 297456 135390 297508 135396
rect 297364 128512 297416 128518
rect 297364 128454 297416 128460
rect 296720 89140 296772 89146
rect 296720 89082 296772 89088
rect 296260 68332 296312 68338
rect 296260 68274 296312 68280
rect 296076 57316 296128 57322
rect 296076 57258 296128 57264
rect 295984 42152 296036 42158
rect 295984 42094 296036 42100
rect 297376 40798 297404 128454
rect 297468 69766 297496 135390
rect 297548 100904 297600 100910
rect 297548 100846 297600 100852
rect 297456 69760 297508 69766
rect 297456 69702 297508 69708
rect 297560 43450 297588 100846
rect 298756 80714 298784 357439
rect 299572 356380 299624 356386
rect 299572 356322 299624 356328
rect 299478 355056 299534 355065
rect 299478 354991 299534 355000
rect 299492 314634 299520 354991
rect 299480 314628 299532 314634
rect 299480 314570 299532 314576
rect 299492 313954 299520 314570
rect 299480 313948 299532 313954
rect 299480 313890 299532 313896
rect 299480 278792 299532 278798
rect 299480 278734 299532 278740
rect 298928 150612 298980 150618
rect 298928 150554 298980 150560
rect 298836 114708 298888 114714
rect 298836 114650 298888 114656
rect 298744 80708 298796 80714
rect 298744 80650 298796 80656
rect 297548 43444 297600 43450
rect 297548 43386 297600 43392
rect 297364 40792 297416 40798
rect 297364 40734 297416 40740
rect 296720 27056 296772 27062
rect 296720 26998 296772 27004
rect 294604 22840 294656 22846
rect 294604 22782 294656 22788
rect 296732 16574 296760 26998
rect 291212 16546 291424 16574
rect 293972 16546 294920 16574
rect 296732 16546 297312 16574
rect 290464 6248 290516 6254
rect 290464 6190 290516 6196
rect 291396 480 291424 16546
rect 292580 3528 292632 3534
rect 292580 3470 292632 3476
rect 293682 3496 293738 3505
rect 292592 480 292620 3470
rect 293682 3431 293738 3440
rect 293696 480 293724 3431
rect 294892 480 294920 16546
rect 296074 3496 296130 3505
rect 296074 3431 296130 3440
rect 296088 480 296116 3431
rect 297284 480 297312 16546
rect 298848 14482 298876 114650
rect 298940 110294 298968 150554
rect 298928 110288 298980 110294
rect 298928 110230 298980 110236
rect 298928 106412 298980 106418
rect 298928 106354 298980 106360
rect 298940 38010 298968 106354
rect 299020 102332 299072 102338
rect 299020 102274 299072 102280
rect 299032 53106 299060 102274
rect 299020 53100 299072 53106
rect 299020 53042 299072 53048
rect 298928 38004 298980 38010
rect 298928 37946 298980 37952
rect 298836 14476 298888 14482
rect 298836 14418 298888 14424
rect 298468 3596 298520 3602
rect 298468 3538 298520 3544
rect 298480 480 298508 3538
rect 299492 3534 299520 278734
rect 299584 94518 299612 356322
rect 299756 355020 299808 355026
rect 299756 354962 299808 354968
rect 299664 248396 299716 248402
rect 299664 248338 299716 248344
rect 299676 247081 299704 248338
rect 299662 247072 299718 247081
rect 299662 247007 299718 247016
rect 299664 242956 299716 242962
rect 299664 242898 299716 242904
rect 299676 224874 299704 242898
rect 299768 241913 299796 354962
rect 301516 342786 301544 702646
rect 305000 700392 305052 700398
rect 305000 700334 305052 700340
rect 303620 360460 303672 360466
rect 303620 360402 303672 360408
rect 301596 356244 301648 356250
rect 301596 356186 301648 356192
rect 300860 342780 300912 342786
rect 300860 342722 300912 342728
rect 301504 342780 301556 342786
rect 301504 342722 301556 342728
rect 299754 241904 299810 241913
rect 299754 241839 299810 241848
rect 300872 235958 300900 342722
rect 300952 271924 301004 271930
rect 300952 271866 301004 271872
rect 300964 241233 300992 271866
rect 300950 241224 301006 241233
rect 300950 241159 301006 241168
rect 300860 235952 300912 235958
rect 300860 235894 300912 235900
rect 299664 224868 299716 224874
rect 299664 224810 299716 224816
rect 300124 164348 300176 164354
rect 300124 164290 300176 164296
rect 300136 126274 300164 164290
rect 300768 151904 300820 151910
rect 300768 151846 300820 151852
rect 300780 149705 300808 151846
rect 300766 149696 300822 149705
rect 300766 149631 300822 149640
rect 300308 149252 300360 149258
rect 300308 149194 300360 149200
rect 300124 126268 300176 126274
rect 300124 126210 300176 126216
rect 300124 110628 300176 110634
rect 300124 110570 300176 110576
rect 299572 94512 299624 94518
rect 299572 94454 299624 94460
rect 300136 54602 300164 110570
rect 300320 109002 300348 149194
rect 301504 124432 301556 124438
rect 301504 124374 301556 124380
rect 300308 108996 300360 109002
rect 300308 108938 300360 108944
rect 300216 107772 300268 107778
rect 300216 107714 300268 107720
rect 300228 62830 300256 107714
rect 300216 62824 300268 62830
rect 300216 62766 300268 62772
rect 300124 54596 300176 54602
rect 300124 54538 300176 54544
rect 301516 32434 301544 124374
rect 301504 32428 301556 32434
rect 301504 32370 301556 32376
rect 301504 13184 301556 13190
rect 301504 13126 301556 13132
rect 299664 10396 299716 10402
rect 299664 10338 299716 10344
rect 299480 3528 299532 3534
rect 299480 3470 299532 3476
rect 299676 480 299704 10338
rect 300768 3528 300820 3534
rect 300768 3470 300820 3476
rect 300780 480 300808 3470
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 13126
rect 301608 3534 301636 356186
rect 302240 312588 302292 312594
rect 302240 312530 302292 312536
rect 302252 311914 302280 312530
rect 302240 311908 302292 311914
rect 302240 311850 302292 311856
rect 302252 227730 302280 311850
rect 302332 290488 302384 290494
rect 302332 290430 302384 290436
rect 302344 289882 302372 290430
rect 302332 289876 302384 289882
rect 302332 289818 302384 289824
rect 302344 238649 302372 289818
rect 302424 251864 302476 251870
rect 302424 251806 302476 251812
rect 302436 251258 302464 251806
rect 302424 251252 302476 251258
rect 302424 251194 302476 251200
rect 302330 238640 302386 238649
rect 302330 238575 302386 238584
rect 302436 231810 302464 251194
rect 302424 231804 302476 231810
rect 302424 231746 302476 231752
rect 302240 227724 302292 227730
rect 302240 227666 302292 227672
rect 303068 160200 303120 160206
rect 303068 160142 303120 160148
rect 301780 149184 301832 149190
rect 301780 149126 301832 149132
rect 301688 117428 301740 117434
rect 301688 117370 301740 117376
rect 301700 26994 301728 117370
rect 301792 111110 301820 149126
rect 302976 132660 303028 132666
rect 302976 132602 303028 132608
rect 302884 120284 302936 120290
rect 302884 120226 302936 120232
rect 301780 111104 301832 111110
rect 301780 111046 301832 111052
rect 301780 107704 301832 107710
rect 301780 107646 301832 107652
rect 301792 60042 301820 107646
rect 301780 60036 301832 60042
rect 301780 59978 301832 59984
rect 302896 28354 302924 120226
rect 302988 58682 303016 132602
rect 303080 121446 303108 160142
rect 303632 145790 303660 360402
rect 303712 307828 303764 307834
rect 303712 307770 303764 307776
rect 303724 234598 303752 307770
rect 305012 235754 305040 700334
rect 310520 700324 310572 700330
rect 310520 700266 310572 700272
rect 319444 700324 319496 700330
rect 319444 700266 319496 700272
rect 306472 699712 306524 699718
rect 306472 699654 306524 699660
rect 305644 320204 305696 320210
rect 305644 320146 305696 320152
rect 305092 276684 305144 276690
rect 305092 276626 305144 276632
rect 305104 276078 305132 276626
rect 305092 276072 305144 276078
rect 305092 276014 305144 276020
rect 305104 267734 305132 276014
rect 305104 267706 305224 267734
rect 305092 263628 305144 263634
rect 305092 263570 305144 263576
rect 305000 235748 305052 235754
rect 305000 235690 305052 235696
rect 303712 234592 303764 234598
rect 303712 234534 303764 234540
rect 304356 146464 304408 146470
rect 304356 146406 304408 146412
rect 303620 145784 303672 145790
rect 303620 145726 303672 145732
rect 304264 135312 304316 135318
rect 304264 135254 304316 135260
rect 303068 121440 303120 121446
rect 303068 121382 303120 121388
rect 303068 111988 303120 111994
rect 303068 111930 303120 111936
rect 302976 58676 303028 58682
rect 302976 58618 303028 58624
rect 303080 49094 303108 111930
rect 303160 109200 303212 109206
rect 303160 109142 303212 109148
rect 303172 75206 303200 109142
rect 303160 75200 303212 75206
rect 303160 75142 303212 75148
rect 304276 71126 304304 135254
rect 304368 117978 304396 146406
rect 304448 145036 304500 145042
rect 304448 144978 304500 144984
rect 304356 117972 304408 117978
rect 304356 117914 304408 117920
rect 304460 112470 304488 144978
rect 305104 142866 305132 263570
rect 305196 237289 305224 267706
rect 305656 257378 305684 320146
rect 306380 294024 306432 294030
rect 306380 293966 306432 293972
rect 305644 257372 305696 257378
rect 305644 257314 305696 257320
rect 305182 237280 305238 237289
rect 305182 237215 305238 237224
rect 305644 207936 305696 207942
rect 305644 207878 305696 207884
rect 305656 178838 305684 207878
rect 305644 178832 305696 178838
rect 305644 178774 305696 178780
rect 306392 176050 306420 293966
rect 306484 234462 306512 699654
rect 309784 590708 309836 590714
rect 309784 590650 309836 590656
rect 308404 357536 308456 357542
rect 308404 357478 308456 357484
rect 306472 234456 306524 234462
rect 306472 234398 306524 234404
rect 305644 176044 305696 176050
rect 305644 175986 305696 175992
rect 306380 176044 306432 176050
rect 306380 175986 306432 175992
rect 307576 176044 307628 176050
rect 307576 175986 307628 175992
rect 305092 142860 305144 142866
rect 305092 142802 305144 142808
rect 305656 131753 305684 175986
rect 307588 175681 307616 175986
rect 307574 175672 307630 175681
rect 307574 175607 307630 175616
rect 307114 175264 307170 175273
rect 307114 175199 307170 175208
rect 306746 174856 306802 174865
rect 306746 174791 306802 174800
rect 306760 174010 306788 174791
rect 306748 174004 306800 174010
rect 306748 173946 306800 173952
rect 306562 173632 306618 173641
rect 306562 173567 306618 173576
rect 306576 170406 306604 173567
rect 306930 173224 306986 173233
rect 306930 173159 306986 173168
rect 306944 172582 306972 173159
rect 306932 172576 306984 172582
rect 306932 172518 306984 172524
rect 306930 172272 306986 172281
rect 306930 172207 306986 172216
rect 306944 171290 306972 172207
rect 306932 171284 306984 171290
rect 306932 171226 306984 171232
rect 306746 170640 306802 170649
rect 306746 170575 306802 170584
rect 306564 170400 306616 170406
rect 306564 170342 306616 170348
rect 306760 169794 306788 170575
rect 306930 169824 306986 169833
rect 306748 169788 306800 169794
rect 306930 169759 306986 169768
rect 306748 169730 306800 169736
rect 306944 164966 306972 169759
rect 307022 165064 307078 165073
rect 307022 164999 307078 165008
rect 306932 164960 306984 164966
rect 306932 164902 306984 164908
rect 306746 163840 306802 163849
rect 306746 163775 306802 163784
rect 306760 162994 306788 163775
rect 306748 162988 306800 162994
rect 306748 162930 306800 162936
rect 306470 161664 306526 161673
rect 306470 161599 306526 161608
rect 306484 160818 306512 161599
rect 306472 160812 306524 160818
rect 306472 160754 306524 160760
rect 306562 160440 306618 160449
rect 306562 160375 306618 160384
rect 306576 152522 306604 160375
rect 306930 160032 306986 160041
rect 306930 159967 306986 159976
rect 306944 158846 306972 159967
rect 306932 158840 306984 158846
rect 306932 158782 306984 158788
rect 306930 158672 306986 158681
rect 306930 158607 306986 158616
rect 306944 157418 306972 158607
rect 306932 157412 306984 157418
rect 306932 157354 306984 157360
rect 306654 152688 306710 152697
rect 306654 152623 306710 152632
rect 306564 152516 306616 152522
rect 306564 152458 306616 152464
rect 306668 145654 306696 152623
rect 306746 150648 306802 150657
rect 306746 150583 306802 150592
rect 306760 150482 306788 150583
rect 306748 150476 306800 150482
rect 306748 150418 306800 150424
rect 306746 149832 306802 149841
rect 306746 149767 306802 149776
rect 306760 149258 306788 149767
rect 306748 149252 306800 149258
rect 306748 149194 306800 149200
rect 306656 145648 306708 145654
rect 306656 145590 306708 145596
rect 306654 143848 306710 143857
rect 306654 143783 306710 143792
rect 305734 143712 305790 143721
rect 305734 143647 305790 143656
rect 305642 131744 305698 131753
rect 305642 131679 305698 131688
rect 304448 112464 304500 112470
rect 304448 112406 304500 112412
rect 304356 111920 304408 111926
rect 304356 111862 304408 111868
rect 304264 71120 304316 71126
rect 304264 71062 304316 71068
rect 304368 50454 304396 111862
rect 304448 106480 304500 106486
rect 304448 106422 304500 106428
rect 304460 65550 304488 106422
rect 305642 104952 305698 104961
rect 305642 104887 305698 104896
rect 304540 103692 304592 103698
rect 304540 103634 304592 103640
rect 304552 69698 304580 103634
rect 304540 69692 304592 69698
rect 304540 69634 304592 69640
rect 304448 65544 304500 65550
rect 304448 65486 304500 65492
rect 304356 50448 304408 50454
rect 304356 50390 304408 50396
rect 303068 49088 303120 49094
rect 303068 49030 303120 49036
rect 305656 36650 305684 104887
rect 305748 104174 305776 143647
rect 306562 143440 306618 143449
rect 306562 143375 306618 143384
rect 306576 142361 306604 143375
rect 306010 142352 306066 142361
rect 306010 142287 306066 142296
rect 306562 142352 306618 142361
rect 306562 142287 306618 142296
rect 305826 107808 305882 107817
rect 305826 107743 305882 107752
rect 305736 104168 305788 104174
rect 305736 104110 305788 104116
rect 305734 100872 305790 100881
rect 305734 100807 305790 100816
rect 305748 39370 305776 100807
rect 305840 58750 305868 107743
rect 306024 105670 306052 142287
rect 306668 142154 306696 143783
rect 306576 142126 306696 142154
rect 306576 141409 306604 142126
rect 306930 142080 306986 142089
rect 306930 142015 306986 142024
rect 306562 141400 306618 141409
rect 306562 141335 306618 141344
rect 306944 140894 306972 142015
rect 307036 141438 307064 164999
rect 307128 162178 307156 175199
rect 307666 174448 307722 174457
rect 307666 174383 307722 174392
rect 307680 174078 307708 174383
rect 307668 174072 307720 174078
rect 307574 174040 307630 174049
rect 307668 174014 307720 174020
rect 307574 173975 307630 173984
rect 307588 173942 307616 173975
rect 307576 173936 307628 173942
rect 307576 173878 307628 173884
rect 307298 172680 307354 172689
rect 307298 172615 307300 172624
rect 307352 172615 307354 172624
rect 307300 172586 307352 172592
rect 307574 171864 307630 171873
rect 307574 171799 307630 171808
rect 307588 171154 307616 171799
rect 307666 171456 307722 171465
rect 307666 171391 307722 171400
rect 307680 171222 307708 171391
rect 307668 171216 307720 171222
rect 307668 171158 307720 171164
rect 307576 171148 307628 171154
rect 307576 171090 307628 171096
rect 307206 171048 307262 171057
rect 307206 170983 307262 170992
rect 307116 162172 307168 162178
rect 307116 162114 307168 162120
rect 307220 160750 307248 170983
rect 307666 170232 307722 170241
rect 307666 170167 307722 170176
rect 307680 169862 307708 170167
rect 307668 169856 307720 169862
rect 307668 169798 307720 169804
rect 307482 169280 307538 169289
rect 307482 169215 307538 169224
rect 307496 168502 307524 169215
rect 307574 168872 307630 168881
rect 307574 168807 307630 168816
rect 307484 168496 307536 168502
rect 307484 168438 307536 168444
rect 307588 168434 307616 168807
rect 307668 168564 307720 168570
rect 307668 168506 307720 168512
rect 307680 168473 307708 168506
rect 307666 168464 307722 168473
rect 307576 168428 307628 168434
rect 307666 168399 307722 168408
rect 307576 168370 307628 168376
rect 307482 168056 307538 168065
rect 307482 167991 307538 168000
rect 307298 167240 307354 167249
rect 307298 167175 307300 167184
rect 307352 167175 307354 167184
rect 307300 167146 307352 167152
rect 307496 167074 307524 167991
rect 307666 167648 307722 167657
rect 307666 167583 307722 167592
rect 307680 167142 307708 167583
rect 307668 167136 307720 167142
rect 307668 167078 307720 167084
rect 307484 167068 307536 167074
rect 307484 167010 307536 167016
rect 307574 166832 307630 166841
rect 307574 166767 307630 166776
rect 307482 166424 307538 166433
rect 307482 166359 307538 166368
rect 307390 165472 307446 165481
rect 307390 165407 307446 165416
rect 307300 164280 307352 164286
rect 307298 164248 307300 164257
rect 307352 164248 307354 164257
rect 307298 164183 307354 164192
rect 307300 163056 307352 163062
rect 307298 163024 307300 163033
rect 307352 163024 307354 163033
rect 307298 162959 307354 162968
rect 307208 160744 307260 160750
rect 307208 160686 307260 160692
rect 307114 159624 307170 159633
rect 307114 159559 307170 159568
rect 307128 149734 307156 159559
rect 307404 159390 307432 165407
rect 307496 164898 307524 166359
rect 307588 165714 307616 166767
rect 307666 165880 307722 165889
rect 307666 165815 307722 165824
rect 307576 165708 307628 165714
rect 307576 165650 307628 165656
rect 307680 165646 307708 165815
rect 307668 165640 307720 165646
rect 307668 165582 307720 165588
rect 307484 164892 307536 164898
rect 307484 164834 307536 164840
rect 307666 164656 307722 164665
rect 307666 164591 307722 164600
rect 307680 164354 307708 164591
rect 307668 164348 307720 164354
rect 307668 164290 307720 164296
rect 307666 163432 307722 163441
rect 307666 163367 307722 163376
rect 307680 162926 307708 163367
rect 307668 162920 307720 162926
rect 307668 162862 307720 162868
rect 307482 162480 307538 162489
rect 307482 162415 307538 162424
rect 307496 161566 307524 162415
rect 307666 162072 307722 162081
rect 307666 162007 307722 162016
rect 307484 161560 307536 161566
rect 307484 161502 307536 161508
rect 307680 161498 307708 162007
rect 307668 161492 307720 161498
rect 307668 161434 307720 161440
rect 307574 161256 307630 161265
rect 307574 161191 307630 161200
rect 307588 160138 307616 161191
rect 307666 160848 307722 160857
rect 307666 160783 307722 160792
rect 307680 160206 307708 160783
rect 307668 160200 307720 160206
rect 307668 160142 307720 160148
rect 307576 160132 307628 160138
rect 307576 160074 307628 160080
rect 307392 159384 307444 159390
rect 307392 159326 307444 159332
rect 307666 159080 307722 159089
rect 307666 159015 307722 159024
rect 307680 158778 307708 159015
rect 307668 158772 307720 158778
rect 307668 158714 307720 158720
rect 307482 158264 307538 158273
rect 307482 158199 307538 158208
rect 307496 157486 307524 158199
rect 307666 157856 307722 157865
rect 307666 157791 307722 157800
rect 307680 157554 307708 157791
rect 307668 157548 307720 157554
rect 307668 157490 307720 157496
rect 307484 157480 307536 157486
rect 307484 157422 307536 157428
rect 307482 157040 307538 157049
rect 307482 156975 307538 156984
rect 307496 156126 307524 156975
rect 307574 156632 307630 156641
rect 307574 156567 307630 156576
rect 307484 156120 307536 156126
rect 307484 156062 307536 156068
rect 307588 156058 307616 156567
rect 307666 156224 307722 156233
rect 307666 156159 307722 156168
rect 307576 156052 307628 156058
rect 307576 155994 307628 156000
rect 307680 155990 307708 156159
rect 307668 155984 307720 155990
rect 307668 155926 307720 155932
rect 307666 155680 307722 155689
rect 307666 155615 307722 155624
rect 307482 155272 307538 155281
rect 307482 155207 307538 155216
rect 307496 154630 307524 155207
rect 307680 154698 307708 155615
rect 307668 154692 307720 154698
rect 307668 154634 307720 154640
rect 307484 154624 307536 154630
rect 307484 154566 307536 154572
rect 307574 154456 307630 154465
rect 307574 154391 307630 154400
rect 307482 154048 307538 154057
rect 307482 153983 307538 153992
rect 307496 153270 307524 153983
rect 307588 153406 307616 154391
rect 307666 153640 307722 153649
rect 307666 153575 307722 153584
rect 307576 153400 307628 153406
rect 307576 153342 307628 153348
rect 307680 153338 307708 153575
rect 307668 153332 307720 153338
rect 307668 153274 307720 153280
rect 307484 153264 307536 153270
rect 307206 153232 307262 153241
rect 307484 153206 307536 153212
rect 307206 153167 307262 153176
rect 307116 149728 307168 149734
rect 307116 149670 307168 149676
rect 307114 145072 307170 145081
rect 307114 145007 307170 145016
rect 307024 141432 307076 141438
rect 307024 141374 307076 141380
rect 306932 140888 306984 140894
rect 306102 140856 306158 140865
rect 306932 140830 306984 140836
rect 306102 140791 306158 140800
rect 306012 105664 306064 105670
rect 306012 105606 306064 105612
rect 306116 105602 306144 140791
rect 306562 137456 306618 137465
rect 306562 137391 306618 137400
rect 306576 136746 306604 137391
rect 306564 136740 306616 136746
rect 306564 136682 306616 136688
rect 307128 133210 307156 145007
rect 307116 133204 307168 133210
rect 307116 133146 307168 133152
rect 307022 131880 307078 131889
rect 307022 131815 307078 131824
rect 306746 131064 306802 131073
rect 306746 130999 306802 131008
rect 306760 129810 306788 130999
rect 306748 129804 306800 129810
rect 306748 129746 306800 129752
rect 306746 127256 306802 127265
rect 306746 127191 306802 127200
rect 306760 127022 306788 127191
rect 306748 127016 306800 127022
rect 306748 126958 306800 126964
rect 306746 126848 306802 126857
rect 306746 126783 306802 126792
rect 306760 125662 306788 126783
rect 306748 125656 306800 125662
rect 306748 125598 306800 125604
rect 306746 125080 306802 125089
rect 306746 125015 306802 125024
rect 306760 124370 306788 125015
rect 306748 124364 306800 124370
rect 306748 124306 306800 124312
rect 306562 123856 306618 123865
rect 306562 123791 306618 123800
rect 306576 123010 306604 123791
rect 306564 123004 306616 123010
rect 306564 122946 306616 122952
rect 307036 122834 307064 131815
rect 307114 127664 307170 127673
rect 307114 127599 307170 127608
rect 307128 127158 307156 127599
rect 307116 127152 307168 127158
rect 307116 127094 307168 127100
rect 307116 124296 307168 124302
rect 307114 124264 307116 124273
rect 307168 124264 307170 124273
rect 307114 124199 307170 124208
rect 307036 122806 307156 122834
rect 306746 122496 306802 122505
rect 306746 122431 306802 122440
rect 306760 121514 306788 122431
rect 306748 121508 306800 121514
rect 306748 121450 306800 121456
rect 306746 121272 306802 121281
rect 306746 121207 306802 121216
rect 306760 120290 306788 121207
rect 306748 120284 306800 120290
rect 306748 120226 306800 120232
rect 306746 119640 306802 119649
rect 306746 119575 306802 119584
rect 306760 118726 306788 119575
rect 306748 118720 306800 118726
rect 306748 118662 306800 118668
rect 307022 116240 307078 116249
rect 307022 116175 307078 116184
rect 306562 112704 306618 112713
rect 306562 112639 306618 112648
rect 306576 111858 306604 112639
rect 306564 111852 306616 111858
rect 306564 111794 306616 111800
rect 306746 111480 306802 111489
rect 306746 111415 306802 111424
rect 306562 111072 306618 111081
rect 306562 111007 306618 111016
rect 306576 110634 306604 111007
rect 306564 110628 306616 110634
rect 306564 110570 306616 110576
rect 306760 110498 306788 111415
rect 306748 110492 306800 110498
rect 306748 110434 306800 110440
rect 306746 110256 306802 110265
rect 306746 110191 306802 110200
rect 306760 109206 306788 110191
rect 306748 109200 306800 109206
rect 306748 109142 306800 109148
rect 306746 105904 306802 105913
rect 306746 105839 306802 105848
rect 306104 105596 306156 105602
rect 306104 105538 306156 105544
rect 306760 105097 306788 105839
rect 305918 105088 305974 105097
rect 305918 105023 305974 105032
rect 306746 105088 306802 105097
rect 306746 105023 306802 105032
rect 305932 66910 305960 105023
rect 306562 103048 306618 103057
rect 306562 102983 306618 102992
rect 306576 102338 306604 102983
rect 306564 102332 306616 102338
rect 306564 102274 306616 102280
rect 306562 101688 306618 101697
rect 306562 101623 306618 101632
rect 306576 100910 306604 101623
rect 306564 100904 306616 100910
rect 306564 100846 306616 100852
rect 306746 100464 306802 100473
rect 306746 100399 306802 100408
rect 306562 100056 306618 100065
rect 306562 99991 306618 100000
rect 306576 99550 306604 99991
rect 306564 99544 306616 99550
rect 306564 99486 306616 99492
rect 306760 99482 306788 100399
rect 306748 99476 306800 99482
rect 306748 99418 306800 99424
rect 306746 99104 306802 99113
rect 306746 99039 306802 99048
rect 306760 98122 306788 99039
rect 306748 98116 306800 98122
rect 306748 98058 306800 98064
rect 306930 96248 306986 96257
rect 306930 96183 306986 96192
rect 306944 95266 306972 96183
rect 306932 95260 306984 95266
rect 306932 95202 306984 95208
rect 305920 66904 305972 66910
rect 305920 66846 305972 66852
rect 305828 58744 305880 58750
rect 305828 58686 305880 58692
rect 307036 42090 307064 116175
rect 307128 87650 307156 122806
rect 307220 116618 307248 153167
rect 307574 152280 307630 152289
rect 307574 152215 307630 152224
rect 307588 151910 307616 152215
rect 307576 151904 307628 151910
rect 307576 151846 307628 151852
rect 307666 151872 307722 151881
rect 307666 151807 307668 151816
rect 307720 151807 307722 151816
rect 307668 151778 307720 151784
rect 307482 151464 307538 151473
rect 307482 151399 307538 151408
rect 307496 150550 307524 151399
rect 307666 151056 307722 151065
rect 307666 150991 307722 151000
rect 307680 150618 307708 150991
rect 307668 150612 307720 150618
rect 307668 150554 307720 150560
rect 307484 150544 307536 150550
rect 307484 150486 307536 150492
rect 307574 150240 307630 150249
rect 307574 150175 307630 150184
rect 307588 149122 307616 150175
rect 307666 149288 307722 149297
rect 307666 149223 307722 149232
rect 307680 149190 307708 149223
rect 307668 149184 307720 149190
rect 307668 149126 307720 149132
rect 307576 149116 307628 149122
rect 307576 149058 307628 149064
rect 307574 148880 307630 148889
rect 307574 148815 307630 148824
rect 307390 148472 307446 148481
rect 307390 148407 307446 148416
rect 307298 147656 307354 147665
rect 307298 147591 307354 147600
rect 307312 145586 307340 147591
rect 307404 146946 307432 148407
rect 307588 147762 307616 148815
rect 307666 148064 307722 148073
rect 307666 147999 307722 148008
rect 307576 147756 307628 147762
rect 307576 147698 307628 147704
rect 307680 147694 307708 147999
rect 307668 147688 307720 147694
rect 307668 147630 307720 147636
rect 307482 147248 307538 147257
rect 307482 147183 307538 147192
rect 307392 146940 307444 146946
rect 307392 146882 307444 146888
rect 307496 146334 307524 147183
rect 307574 146840 307630 146849
rect 307574 146775 307630 146784
rect 307588 146402 307616 146775
rect 307668 146464 307720 146470
rect 307666 146432 307668 146441
rect 307720 146432 307722 146441
rect 307576 146396 307628 146402
rect 307666 146367 307722 146376
rect 307576 146338 307628 146344
rect 307484 146328 307536 146334
rect 307484 146270 307536 146276
rect 307482 145888 307538 145897
rect 307482 145823 307538 145832
rect 307300 145580 307352 145586
rect 307300 145522 307352 145528
rect 307496 144974 307524 145823
rect 307666 145480 307722 145489
rect 307666 145415 307722 145424
rect 307680 145042 307708 145415
rect 307668 145036 307720 145042
rect 307668 144978 307720 144984
rect 307484 144968 307536 144974
rect 307484 144910 307536 144916
rect 307574 144664 307630 144673
rect 307574 144599 307630 144608
rect 307588 143721 307616 144599
rect 307666 144256 307722 144265
rect 307666 144191 307722 144200
rect 307574 143712 307630 143721
rect 307574 143647 307630 143656
rect 307680 143614 307708 144191
rect 307668 143608 307720 143614
rect 307668 143550 307720 143556
rect 307574 143032 307630 143041
rect 307574 142967 307630 142976
rect 307588 142254 307616 142967
rect 307666 142488 307722 142497
rect 307666 142423 307722 142432
rect 307680 142322 307708 142423
rect 307668 142316 307720 142322
rect 307668 142258 307720 142264
rect 307576 142248 307628 142254
rect 307576 142190 307628 142196
rect 307298 141672 307354 141681
rect 307298 141607 307354 141616
rect 307208 116612 307260 116618
rect 307208 116554 307260 116560
rect 307312 113174 307340 141607
rect 307390 141264 307446 141273
rect 307390 141199 307446 141208
rect 307404 133906 307432 141199
rect 307482 140448 307538 140457
rect 307482 140383 307538 140392
rect 307496 139466 307524 140383
rect 307574 140040 307630 140049
rect 307574 139975 307630 139984
rect 307588 139534 307616 139975
rect 307666 139632 307722 139641
rect 307666 139567 307668 139576
rect 307720 139567 307722 139576
rect 307668 139538 307720 139544
rect 307576 139528 307628 139534
rect 307576 139470 307628 139476
rect 307484 139460 307536 139466
rect 307484 139402 307536 139408
rect 307482 139088 307538 139097
rect 307482 139023 307538 139032
rect 307496 138038 307524 139023
rect 307574 138680 307630 138689
rect 307574 138615 307630 138624
rect 307588 138106 307616 138615
rect 307666 138272 307722 138281
rect 307666 138207 307722 138216
rect 307680 138174 307708 138207
rect 307668 138168 307720 138174
rect 307668 138110 307720 138116
rect 307576 138100 307628 138106
rect 307576 138042 307628 138048
rect 307484 138032 307536 138038
rect 307484 137974 307536 137980
rect 307574 137864 307630 137873
rect 307574 137799 307630 137808
rect 307588 136814 307616 137799
rect 307666 137048 307722 137057
rect 307666 136983 307722 136992
rect 307576 136808 307628 136814
rect 307576 136750 307628 136756
rect 307680 136678 307708 136983
rect 307668 136672 307720 136678
rect 307482 136640 307538 136649
rect 307668 136614 307720 136620
rect 307482 136575 307538 136584
rect 307496 135522 307524 136575
rect 307574 136232 307630 136241
rect 307574 136167 307630 136176
rect 307484 135516 307536 135522
rect 307484 135458 307536 135464
rect 307588 135386 307616 136167
rect 307666 135688 307722 135697
rect 307666 135623 307722 135632
rect 307680 135454 307708 135623
rect 307668 135448 307720 135454
rect 307668 135390 307720 135396
rect 307576 135380 307628 135386
rect 307576 135322 307628 135328
rect 307668 135312 307720 135318
rect 307666 135280 307668 135289
rect 307720 135280 307722 135289
rect 307666 135215 307722 135224
rect 307482 134872 307538 134881
rect 307482 134807 307538 134816
rect 307496 134026 307524 134807
rect 307666 134464 307722 134473
rect 307666 134399 307722 134408
rect 307680 134094 307708 134399
rect 307668 134088 307720 134094
rect 307574 134056 307630 134065
rect 307484 134020 307536 134026
rect 307668 134030 307720 134036
rect 307574 133991 307630 134000
rect 307484 133962 307536 133968
rect 307588 133958 307616 133991
rect 307576 133952 307628 133958
rect 307404 133878 307524 133906
rect 307576 133894 307628 133900
rect 307390 133648 307446 133657
rect 307390 133583 307446 133592
rect 307404 132530 307432 133583
rect 307392 132524 307444 132530
rect 307392 132466 307444 132472
rect 307390 129296 307446 129305
rect 307390 129231 307446 129240
rect 307404 128450 307432 129231
rect 307392 128444 307444 128450
rect 307392 128386 307444 128392
rect 307496 119406 307524 133878
rect 307574 133240 307630 133249
rect 307574 133175 307630 133184
rect 307588 132666 307616 133175
rect 307666 132696 307722 132705
rect 307576 132660 307628 132666
rect 307666 132631 307722 132640
rect 307576 132602 307628 132608
rect 307680 132598 307708 132631
rect 307668 132592 307720 132598
rect 307668 132534 307720 132540
rect 307666 132288 307722 132297
rect 307666 132223 307722 132232
rect 307680 131170 307708 132223
rect 307668 131164 307720 131170
rect 307668 131106 307720 131112
rect 307574 130248 307630 130257
rect 307574 130183 307630 130192
rect 307588 129878 307616 130183
rect 307668 129940 307720 129946
rect 307668 129882 307720 129888
rect 307576 129872 307628 129878
rect 307680 129849 307708 129882
rect 307576 129814 307628 129820
rect 307666 129840 307722 129849
rect 307666 129775 307722 129784
rect 307666 128888 307722 128897
rect 307666 128823 307722 128832
rect 307680 128518 307708 128823
rect 307668 128512 307720 128518
rect 307574 128480 307630 128489
rect 307668 128454 307720 128460
rect 307574 128415 307630 128424
rect 307588 128382 307616 128415
rect 307576 128376 307628 128382
rect 307576 128318 307628 128324
rect 307666 128072 307722 128081
rect 307666 128007 307722 128016
rect 307680 127090 307708 128007
rect 307668 127084 307720 127090
rect 307668 127026 307720 127032
rect 307666 125896 307722 125905
rect 307666 125831 307722 125840
rect 307680 125730 307708 125831
rect 307668 125724 307720 125730
rect 307668 125666 307720 125672
rect 307574 125488 307630 125497
rect 307574 125423 307630 125432
rect 307588 124234 307616 125423
rect 307666 124672 307722 124681
rect 307666 124607 307722 124616
rect 307680 124438 307708 124607
rect 307668 124432 307720 124438
rect 307668 124374 307720 124380
rect 307576 124228 307628 124234
rect 307576 124170 307628 124176
rect 307574 123448 307630 123457
rect 307574 123383 307630 123392
rect 307588 122874 307616 123383
rect 307666 123040 307722 123049
rect 307666 122975 307722 122984
rect 307680 122942 307708 122975
rect 307668 122936 307720 122942
rect 307668 122878 307720 122884
rect 307576 122868 307628 122874
rect 307576 122810 307628 122816
rect 307574 122088 307630 122097
rect 307574 122023 307630 122032
rect 307588 121650 307616 122023
rect 307666 121680 307722 121689
rect 307576 121644 307628 121650
rect 307666 121615 307722 121624
rect 307576 121586 307628 121592
rect 307680 121582 307708 121615
rect 307668 121576 307720 121582
rect 307668 121518 307720 121524
rect 307574 120864 307630 120873
rect 307574 120799 307630 120808
rect 307588 120222 307616 120799
rect 307666 120456 307722 120465
rect 307666 120391 307722 120400
rect 307576 120216 307628 120222
rect 307576 120158 307628 120164
rect 307680 120154 307708 120391
rect 307668 120148 307720 120154
rect 307668 120090 307720 120096
rect 307666 120048 307722 120057
rect 307666 119983 307722 119992
rect 307484 119400 307536 119406
rect 307484 119342 307536 119348
rect 307680 118794 307708 119983
rect 307668 118788 307720 118794
rect 307668 118730 307720 118736
rect 307482 118280 307538 118289
rect 307482 118215 307538 118224
rect 307496 117366 307524 118215
rect 307666 117872 307722 117881
rect 307666 117807 307722 117816
rect 307680 117434 307708 117807
rect 307668 117428 307720 117434
rect 307668 117370 307720 117376
rect 307484 117360 307536 117366
rect 307484 117302 307536 117308
rect 307666 117056 307722 117065
rect 307666 116991 307722 117000
rect 307482 116648 307538 116657
rect 307482 116583 307538 116592
rect 307496 116074 307524 116583
rect 307484 116068 307536 116074
rect 307484 116010 307536 116016
rect 307680 116006 307708 116991
rect 307668 116000 307720 116006
rect 307668 115942 307720 115948
rect 307482 115696 307538 115705
rect 307482 115631 307538 115640
rect 307496 114578 307524 115631
rect 307574 115288 307630 115297
rect 307574 115223 307630 115232
rect 307588 114714 307616 115223
rect 307666 114880 307722 114889
rect 307666 114815 307722 114824
rect 307576 114708 307628 114714
rect 307576 114650 307628 114656
rect 307680 114646 307708 114815
rect 307668 114640 307720 114646
rect 307668 114582 307720 114588
rect 307484 114572 307536 114578
rect 307484 114514 307536 114520
rect 307666 113656 307722 113665
rect 307666 113591 307722 113600
rect 307576 113280 307628 113286
rect 307574 113248 307576 113257
rect 307628 113248 307630 113257
rect 307680 113218 307708 113591
rect 307574 113183 307630 113192
rect 307668 113212 307720 113218
rect 307220 113146 307340 113174
rect 307668 113154 307720 113160
rect 307220 107030 307248 113146
rect 307666 112296 307722 112305
rect 307666 112231 307722 112240
rect 307300 111988 307352 111994
rect 307300 111930 307352 111936
rect 307312 111897 307340 111930
rect 307680 111926 307708 112231
rect 307668 111920 307720 111926
rect 307298 111888 307354 111897
rect 307668 111862 307720 111868
rect 307298 111823 307354 111832
rect 307298 110664 307354 110673
rect 307298 110599 307354 110608
rect 307312 110566 307340 110599
rect 307300 110560 307352 110566
rect 307300 110502 307352 110508
rect 307574 109848 307630 109857
rect 307574 109783 307630 109792
rect 307588 109070 307616 109783
rect 307666 109304 307722 109313
rect 307666 109239 307722 109248
rect 307680 109138 307708 109239
rect 307668 109132 307720 109138
rect 307668 109074 307720 109080
rect 307576 109064 307628 109070
rect 307576 109006 307628 109012
rect 307574 108896 307630 108905
rect 307574 108831 307630 108840
rect 307482 108488 307538 108497
rect 307482 108423 307538 108432
rect 307300 107772 307352 107778
rect 307300 107714 307352 107720
rect 307312 107681 307340 107714
rect 307496 107710 307524 108423
rect 307588 107817 307616 108831
rect 307666 108080 307722 108089
rect 307666 108015 307722 108024
rect 307680 107914 307708 108015
rect 307668 107908 307720 107914
rect 307668 107850 307720 107856
rect 307574 107808 307630 107817
rect 307574 107743 307630 107752
rect 307484 107704 307536 107710
rect 307298 107672 307354 107681
rect 307484 107646 307536 107652
rect 307298 107607 307354 107616
rect 307482 107264 307538 107273
rect 307482 107199 307538 107208
rect 307208 107024 307260 107030
rect 307208 106966 307260 106972
rect 307298 106856 307354 106865
rect 307298 106791 307354 106800
rect 307312 106350 307340 106791
rect 307496 106418 307524 107199
rect 307668 106480 307720 106486
rect 307666 106448 307668 106457
rect 307720 106448 307722 106457
rect 307484 106412 307536 106418
rect 307666 106383 307722 106392
rect 307484 106354 307536 106360
rect 307300 106344 307352 106350
rect 307300 106286 307352 106292
rect 307666 105496 307722 105505
rect 307666 105431 307722 105440
rect 307680 105058 307708 105431
rect 307668 105052 307720 105058
rect 307668 104994 307720 105000
rect 307482 104680 307538 104689
rect 307482 104615 307538 104624
rect 307496 103630 307524 104615
rect 307666 104272 307722 104281
rect 307666 104207 307722 104216
rect 307574 103864 307630 103873
rect 307574 103799 307630 103808
rect 307484 103624 307536 103630
rect 307484 103566 307536 103572
rect 307588 103562 307616 103799
rect 307680 103698 307708 104207
rect 307668 103692 307720 103698
rect 307668 103634 307720 103640
rect 307576 103556 307628 103562
rect 307576 103498 307628 103504
rect 307574 103456 307630 103465
rect 307574 103391 307630 103400
rect 307588 102270 307616 103391
rect 307666 102504 307722 102513
rect 307666 102439 307722 102448
rect 307576 102264 307628 102270
rect 307576 102206 307628 102212
rect 307680 102202 307708 102439
rect 307668 102196 307720 102202
rect 307668 102138 307720 102144
rect 307482 102096 307538 102105
rect 307482 102031 307538 102040
rect 307496 100881 307524 102031
rect 307666 101280 307722 101289
rect 307666 101215 307722 101224
rect 307680 100978 307708 101215
rect 307668 100972 307720 100978
rect 307668 100914 307720 100920
rect 307482 100872 307538 100881
rect 307482 100807 307538 100816
rect 307666 100872 307722 100881
rect 307666 100807 307668 100816
rect 307720 100807 307722 100816
rect 307668 100778 307720 100784
rect 307666 99648 307722 99657
rect 307666 99583 307722 99592
rect 307680 99414 307708 99583
rect 307668 99408 307720 99414
rect 307668 99350 307720 99356
rect 307206 98696 307262 98705
rect 307206 98631 307262 98640
rect 307116 87644 307168 87650
rect 307116 87586 307168 87592
rect 307220 64190 307248 98631
rect 307666 98288 307722 98297
rect 307666 98223 307722 98232
rect 307680 98054 307708 98223
rect 307668 98048 307720 98054
rect 307668 97990 307720 97996
rect 307574 97880 307630 97889
rect 307574 97815 307630 97824
rect 307298 97472 307354 97481
rect 307298 97407 307354 97416
rect 307312 79354 307340 97407
rect 307588 96762 307616 97815
rect 307666 97064 307722 97073
rect 307666 96999 307722 97008
rect 307680 96830 307708 96999
rect 307668 96824 307720 96830
rect 307668 96766 307720 96772
rect 307576 96756 307628 96762
rect 307576 96698 307628 96704
rect 307668 96688 307720 96694
rect 307666 96656 307668 96665
rect 307720 96656 307722 96665
rect 307666 96591 307722 96600
rect 307300 79348 307352 79354
rect 307300 79290 307352 79296
rect 307208 64184 307260 64190
rect 307208 64126 307260 64132
rect 307024 42084 307076 42090
rect 307024 42026 307076 42032
rect 305736 39364 305788 39370
rect 305736 39306 305788 39312
rect 305644 36644 305696 36650
rect 305644 36586 305696 36592
rect 302884 28348 302936 28354
rect 302884 28290 302936 28296
rect 301688 26988 301740 26994
rect 301688 26930 301740 26936
rect 303618 25664 303674 25673
rect 303618 25599 303674 25608
rect 303632 16574 303660 25599
rect 303632 16546 303936 16574
rect 303158 6216 303214 6225
rect 303158 6151 303214 6160
rect 301596 3528 301648 3534
rect 301596 3470 301648 3476
rect 303172 480 303200 6151
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 308416 8974 308444 357478
rect 308496 339516 308548 339522
rect 308496 339458 308548 339464
rect 308508 84862 308536 339458
rect 309796 312594 309824 590650
rect 309784 312588 309836 312594
rect 309784 312530 309836 312536
rect 309876 295384 309928 295390
rect 309876 295326 309928 295332
rect 309692 285728 309744 285734
rect 309692 285670 309744 285676
rect 308588 202496 308640 202502
rect 308588 202438 308640 202444
rect 308496 84856 308548 84862
rect 308496 84798 308548 84804
rect 308404 8968 308456 8974
rect 308404 8910 308456 8916
rect 305550 6352 305606 6361
rect 305550 6287 305606 6296
rect 305564 480 305592 6287
rect 308600 3398 308628 202438
rect 309138 114472 309194 114481
rect 309138 114407 309194 114416
rect 309152 113121 309180 114407
rect 309138 113112 309194 113121
rect 309138 113047 309194 113056
rect 309704 79354 309732 285670
rect 309784 260908 309836 260914
rect 309784 260850 309836 260856
rect 309692 79348 309744 79354
rect 309692 79290 309744 79296
rect 309796 4826 309824 260850
rect 309888 83570 309916 295326
rect 310532 238882 310560 700266
rect 315304 364540 315356 364546
rect 315304 364482 315356 364488
rect 311900 358964 311952 358970
rect 311900 358906 311952 358912
rect 311164 327140 311216 327146
rect 311164 327082 311216 327088
rect 310980 283620 311032 283626
rect 310980 283562 311032 283568
rect 310992 282946 311020 283562
rect 310612 282940 310664 282946
rect 310612 282882 310664 282888
rect 310980 282940 311032 282946
rect 310980 282882 311032 282888
rect 310520 238876 310572 238882
rect 310520 238818 310572 238824
rect 310624 235890 310652 282882
rect 311176 259418 311204 327082
rect 311164 259412 311216 259418
rect 311164 259354 311216 259360
rect 310612 235884 310664 235890
rect 310612 235826 310664 235832
rect 311912 227186 311940 358906
rect 313280 356312 313332 356318
rect 313280 356254 313332 356260
rect 313292 229809 313320 356254
rect 314660 305652 314712 305658
rect 314660 305594 314712 305600
rect 314672 305046 314700 305594
rect 314660 305040 314712 305046
rect 314660 304982 314712 304988
rect 314672 237318 314700 304982
rect 314660 237312 314712 237318
rect 314660 237254 314712 237260
rect 313278 229800 313334 229809
rect 313278 229735 313334 229744
rect 311900 227180 311952 227186
rect 311900 227122 311952 227128
rect 311164 224324 311216 224330
rect 311164 224266 311216 224272
rect 311176 177449 311204 224266
rect 313924 220176 313976 220182
rect 313924 220118 313976 220124
rect 311256 214600 311308 214606
rect 311256 214542 311308 214548
rect 311162 177440 311218 177449
rect 311162 177375 311218 177384
rect 311268 176662 311296 214542
rect 312544 196920 312596 196926
rect 312544 196862 312596 196868
rect 312556 178906 312584 196862
rect 312544 178900 312596 178906
rect 312544 178842 312596 178848
rect 313936 178809 313964 220118
rect 313922 178800 313978 178809
rect 313922 178735 313978 178744
rect 315316 177313 315344 364482
rect 317420 357604 317472 357610
rect 317420 357546 317472 357552
rect 315396 216028 315448 216034
rect 315396 215970 315448 215976
rect 315408 177410 315436 215970
rect 317432 189689 317460 357546
rect 319456 251870 319484 700266
rect 324964 698964 325016 698970
rect 324964 698906 325016 698912
rect 319444 251864 319496 251870
rect 319444 251806 319496 251812
rect 319444 249824 319496 249830
rect 319444 249766 319496 249772
rect 319456 231130 319484 249766
rect 324976 248402 325004 698906
rect 331232 376038 331260 702986
rect 348804 697610 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 348792 697604 348844 697610
rect 348792 697546 348844 697552
rect 337384 616888 337436 616894
rect 337384 616830 337436 616836
rect 331220 376032 331272 376038
rect 331220 375974 331272 375980
rect 327724 371272 327776 371278
rect 327724 371214 327776 371220
rect 324964 248396 325016 248402
rect 324964 248338 325016 248344
rect 323584 239012 323636 239018
rect 323584 238954 323636 238960
rect 319444 231124 319496 231130
rect 319444 231066 319496 231072
rect 319444 225752 319496 225758
rect 319444 225694 319496 225700
rect 318064 218952 318116 218958
rect 318064 218894 318116 218900
rect 317418 189680 317474 189689
rect 317418 189615 317474 189624
rect 318076 177546 318104 218894
rect 318156 194064 318208 194070
rect 318156 194006 318208 194012
rect 318064 177540 318116 177546
rect 318064 177482 318116 177488
rect 315396 177404 315448 177410
rect 315396 177346 315448 177352
rect 315302 177304 315358 177313
rect 315302 177239 315358 177248
rect 316038 176760 316094 176769
rect 318168 176730 318196 194006
rect 318340 180260 318392 180266
rect 318340 180202 318392 180208
rect 318352 177478 318380 180202
rect 318708 178764 318760 178770
rect 318708 178706 318760 178712
rect 318340 177472 318392 177478
rect 318340 177414 318392 177420
rect 316038 176695 316094 176704
rect 318156 176724 318208 176730
rect 311256 176656 311308 176662
rect 311256 176598 311308 176604
rect 316052 175930 316080 176695
rect 318156 176666 318208 176672
rect 316020 175902 316080 175930
rect 318720 175914 318748 178706
rect 319456 176225 319484 225694
rect 319536 217320 319588 217326
rect 319536 217262 319588 217268
rect 319442 176216 319498 176225
rect 319442 176151 319498 176160
rect 319548 175982 319576 217262
rect 322940 213240 322992 213246
rect 322940 213182 322992 213188
rect 319628 198008 319680 198014
rect 319628 197950 319680 197956
rect 319640 176050 319668 197950
rect 320824 196716 320876 196722
rect 320824 196658 320876 196664
rect 320180 186992 320232 186998
rect 320180 186934 320232 186940
rect 320192 176769 320220 186934
rect 320836 176769 320864 196658
rect 321284 187060 321336 187066
rect 321284 187002 321336 187008
rect 320178 176760 320234 176769
rect 320178 176695 320234 176704
rect 320822 176760 320878 176769
rect 320822 176695 320878 176704
rect 319628 176044 319680 176050
rect 319628 175986 319680 175992
rect 319536 175976 319588 175982
rect 319536 175918 319588 175924
rect 318708 175908 318760 175914
rect 318708 175850 318760 175856
rect 321296 172689 321324 187002
rect 321744 185768 321796 185774
rect 321744 185710 321796 185716
rect 321650 176760 321706 176769
rect 321560 176724 321612 176730
rect 321650 176695 321706 176704
rect 321560 176666 321612 176672
rect 321468 176656 321520 176662
rect 321468 176598 321520 176604
rect 321480 175817 321508 176598
rect 321466 175808 321522 175817
rect 321466 175743 321522 175752
rect 321282 172680 321338 172689
rect 321282 172615 321338 172624
rect 321466 171456 321522 171465
rect 321466 171391 321522 171400
rect 321480 169697 321508 171391
rect 321466 169688 321522 169697
rect 321466 169623 321522 169632
rect 321572 132705 321600 176666
rect 321664 150385 321692 176695
rect 321756 167521 321784 185710
rect 321836 177472 321888 177478
rect 321836 177414 321888 177420
rect 321848 175273 321876 177414
rect 321928 175908 321980 175914
rect 321928 175850 321980 175856
rect 321834 175264 321890 175273
rect 321834 175199 321890 175208
rect 321940 171193 321968 175850
rect 321926 171184 321982 171193
rect 321926 171119 321982 171128
rect 321742 167512 321798 167521
rect 321742 167447 321798 167456
rect 321650 150376 321706 150385
rect 321650 150311 321706 150320
rect 321558 132696 321614 132705
rect 321558 132631 321614 132640
rect 322952 103193 322980 213182
rect 323124 185700 323176 185706
rect 323124 185642 323176 185648
rect 323030 184240 323086 184249
rect 323030 184175 323086 184184
rect 323044 150929 323072 184175
rect 323136 165481 323164 185642
rect 323122 165472 323178 165481
rect 323122 165407 323178 165416
rect 323030 150920 323086 150929
rect 323030 150855 323086 150864
rect 323596 143546 323624 238954
rect 324596 227044 324648 227050
rect 324596 226986 324648 226992
rect 324412 221536 324464 221542
rect 324412 221478 324464 221484
rect 324424 174049 324452 221478
rect 324608 190454 324636 226986
rect 325700 214668 325752 214674
rect 325700 214610 325752 214616
rect 324608 190426 324728 190454
rect 324504 189848 324556 189854
rect 324504 189790 324556 189796
rect 324410 174040 324466 174049
rect 324410 173975 324466 173984
rect 324320 173868 324372 173874
rect 324320 173810 324372 173816
rect 324332 173233 324360 173810
rect 324318 173224 324374 173233
rect 324318 173159 324374 173168
rect 324320 169720 324372 169726
rect 324320 169662 324372 169668
rect 324332 168609 324360 169662
rect 324318 168600 324374 168609
rect 324318 168535 324374 168544
rect 324320 168360 324372 168366
rect 324320 168302 324372 168308
rect 324332 167793 324360 168302
rect 324318 167784 324374 167793
rect 324318 167719 324374 167728
rect 324320 165572 324372 165578
rect 324320 165514 324372 165520
rect 324332 164801 324360 165514
rect 324318 164792 324374 164801
rect 324318 164727 324374 164736
rect 324412 164212 324464 164218
rect 324412 164154 324464 164160
rect 324320 164144 324372 164150
rect 324320 164086 324372 164092
rect 324332 163985 324360 164086
rect 324318 163976 324374 163985
rect 324318 163911 324374 163920
rect 324424 163169 324452 164154
rect 324410 163160 324466 163169
rect 324410 163095 324466 163104
rect 324412 162852 324464 162858
rect 324412 162794 324464 162800
rect 324320 162784 324372 162790
rect 324320 162726 324372 162732
rect 324332 162489 324360 162726
rect 324318 162480 324374 162489
rect 324318 162415 324374 162424
rect 324424 161673 324452 162794
rect 324410 161664 324466 161673
rect 324410 161599 324466 161608
rect 324320 161424 324372 161430
rect 324320 161366 324372 161372
rect 324332 160857 324360 161366
rect 324412 161356 324464 161362
rect 324412 161298 324464 161304
rect 324318 160848 324374 160857
rect 324318 160783 324374 160792
rect 324424 160177 324452 161298
rect 324410 160168 324466 160177
rect 324410 160103 324466 160112
rect 324320 160064 324372 160070
rect 324320 160006 324372 160012
rect 324332 159361 324360 160006
rect 324318 159352 324374 159361
rect 324318 159287 324374 159296
rect 324412 158704 324464 158710
rect 324412 158646 324464 158652
rect 324320 158636 324372 158642
rect 324320 158578 324372 158584
rect 324332 158545 324360 158578
rect 324318 158536 324374 158545
rect 324318 158471 324374 158480
rect 324424 157865 324452 158646
rect 324410 157856 324466 157865
rect 324410 157791 324466 157800
rect 324320 157276 324372 157282
rect 324320 157218 324372 157224
rect 324332 157049 324360 157218
rect 324318 157040 324374 157049
rect 324318 156975 324374 156984
rect 324320 155916 324372 155922
rect 324320 155858 324372 155864
rect 324332 155553 324360 155858
rect 324412 155848 324464 155854
rect 324412 155790 324464 155796
rect 324318 155544 324374 155553
rect 324318 155479 324374 155488
rect 324424 154737 324452 155790
rect 324410 154728 324466 154737
rect 324410 154663 324466 154672
rect 324320 154556 324372 154562
rect 324320 154498 324372 154504
rect 324332 154057 324360 154498
rect 324318 154048 324374 154057
rect 324318 153983 324374 153992
rect 324320 153332 324372 153338
rect 324320 153274 324372 153280
rect 324332 153241 324360 153274
rect 324318 153232 324374 153241
rect 324318 153167 324374 153176
rect 324516 152425 324544 189790
rect 324700 166297 324728 190426
rect 324686 166288 324742 166297
rect 324686 166223 324742 166232
rect 324502 152416 324558 152425
rect 324502 152351 324558 152360
rect 324320 151768 324372 151774
rect 324318 151736 324320 151745
rect 324372 151736 324374 151745
rect 324318 151671 324374 151680
rect 324320 150408 324372 150414
rect 324320 150350 324372 150356
rect 324332 149433 324360 150350
rect 324318 149424 324374 149433
rect 324318 149359 324374 149368
rect 324320 148980 324372 148986
rect 324320 148922 324372 148928
rect 324332 148617 324360 148922
rect 324412 148844 324464 148850
rect 324412 148786 324464 148792
rect 324318 148608 324374 148617
rect 324318 148543 324374 148552
rect 324424 147801 324452 148786
rect 324410 147792 324466 147801
rect 324410 147727 324466 147736
rect 324320 147620 324372 147626
rect 324320 147562 324372 147568
rect 324332 147121 324360 147562
rect 324318 147112 324374 147121
rect 324318 147047 324374 147056
rect 324320 144900 324372 144906
rect 324320 144842 324372 144848
rect 324332 143993 324360 144842
rect 324318 143984 324374 143993
rect 324318 143919 324374 143928
rect 323584 143540 323636 143546
rect 323584 143482 323636 143488
rect 324504 143540 324556 143546
rect 324504 143482 324556 143488
rect 324596 143540 324648 143546
rect 324596 143482 324648 143488
rect 324320 143472 324372 143478
rect 324320 143414 324372 143420
rect 324332 143177 324360 143414
rect 324318 143168 324374 143177
rect 324318 143103 324374 143112
rect 324320 142044 324372 142050
rect 324320 141986 324372 141992
rect 324332 141681 324360 141986
rect 324318 141672 324374 141681
rect 324318 141607 324374 141616
rect 324320 140752 324372 140758
rect 324320 140694 324372 140700
rect 324332 140185 324360 140694
rect 324318 140176 324374 140185
rect 324318 140111 324374 140120
rect 324320 139392 324372 139398
rect 324318 139360 324320 139369
rect 324372 139360 324374 139369
rect 324318 139295 324374 139304
rect 324412 137964 324464 137970
rect 324412 137906 324464 137912
rect 324320 137896 324372 137902
rect 324318 137864 324320 137873
rect 324372 137864 324374 137873
rect 324318 137799 324374 137808
rect 324424 137057 324452 137906
rect 324410 137048 324466 137057
rect 324410 136983 324466 136992
rect 324412 136604 324464 136610
rect 324412 136546 324464 136552
rect 324320 136400 324372 136406
rect 324318 136368 324320 136377
rect 324372 136368 324374 136377
rect 324318 136303 324374 136312
rect 324424 135561 324452 136546
rect 324410 135552 324466 135561
rect 324410 135487 324466 135496
rect 324516 133249 324544 143482
rect 324608 142497 324636 143482
rect 324594 142488 324650 142497
rect 324594 142423 324650 142432
rect 324596 142112 324648 142118
rect 324596 142054 324648 142060
rect 324608 140865 324636 142054
rect 324594 140856 324650 140865
rect 324594 140791 324650 140800
rect 324502 133240 324558 133249
rect 324502 133175 324558 133184
rect 324320 132456 324372 132462
rect 324320 132398 324372 132404
rect 324332 131753 324360 132398
rect 324318 131744 324374 131753
rect 324318 131679 324374 131688
rect 324320 131096 324372 131102
rect 324320 131038 324372 131044
rect 324332 130937 324360 131038
rect 324412 131028 324464 131034
rect 324412 130970 324464 130976
rect 324318 130928 324374 130937
rect 324318 130863 324374 130872
rect 324424 130121 324452 130970
rect 324410 130112 324466 130121
rect 324410 130047 324466 130056
rect 324320 129736 324372 129742
rect 324320 129678 324372 129684
rect 324332 129441 324360 129678
rect 324412 129668 324464 129674
rect 324412 129610 324464 129616
rect 324318 129432 324374 129441
rect 324318 129367 324374 129376
rect 324424 128625 324452 129610
rect 324410 128616 324466 128625
rect 324410 128551 324466 128560
rect 324320 128308 324372 128314
rect 324320 128250 324372 128256
rect 324332 127809 324360 128250
rect 324412 127968 324464 127974
rect 324412 127910 324464 127916
rect 324318 127800 324374 127809
rect 324318 127735 324374 127744
rect 324424 127129 324452 127910
rect 324410 127120 324466 127129
rect 324410 127055 324466 127064
rect 324320 125588 324372 125594
rect 324320 125530 324372 125536
rect 324332 124817 324360 125530
rect 324318 124808 324374 124817
rect 324318 124743 324374 124752
rect 324320 124160 324372 124166
rect 324320 124102 324372 124108
rect 324332 123185 324360 124102
rect 324318 123176 324374 123185
rect 324318 123111 324374 123120
rect 324320 122800 324372 122806
rect 324320 122742 324372 122748
rect 324332 122505 324360 122742
rect 324318 122496 324374 122505
rect 324318 122431 324374 122440
rect 324412 121440 324464 121446
rect 324412 121382 324464 121388
rect 324320 121372 324372 121378
rect 324320 121314 324372 121320
rect 324332 120873 324360 121314
rect 324318 120864 324374 120873
rect 324318 120799 324374 120808
rect 324424 120193 324452 121382
rect 324410 120184 324466 120193
rect 324410 120119 324466 120128
rect 324320 120080 324372 120086
rect 324320 120022 324372 120028
rect 324332 119377 324360 120022
rect 324318 119368 324374 119377
rect 324318 119303 324374 119312
rect 324320 118652 324372 118658
rect 324320 118594 324372 118600
rect 324332 118561 324360 118594
rect 324412 118584 324464 118590
rect 324318 118552 324374 118561
rect 324412 118526 324464 118532
rect 324318 118487 324374 118496
rect 324424 117881 324452 118526
rect 324410 117872 324466 117881
rect 324410 117807 324466 117816
rect 324320 117292 324372 117298
rect 324320 117234 324372 117240
rect 324332 117065 324360 117234
rect 324412 117224 324464 117230
rect 324412 117166 324464 117172
rect 324318 117056 324374 117065
rect 324318 116991 324374 117000
rect 324424 116385 324452 117166
rect 324410 116376 324466 116385
rect 324410 116311 324466 116320
rect 324320 115932 324372 115938
rect 324320 115874 324372 115880
rect 324332 115569 324360 115874
rect 324318 115560 324374 115569
rect 324318 115495 324374 115504
rect 324412 114504 324464 114510
rect 324412 114446 324464 114452
rect 324320 114436 324372 114442
rect 324320 114378 324372 114384
rect 324332 114073 324360 114378
rect 324318 114064 324374 114073
rect 324318 113999 324374 114008
rect 324424 113257 324452 114446
rect 324410 113248 324466 113257
rect 324410 113183 324466 113192
rect 324320 113144 324372 113150
rect 324320 113086 324372 113092
rect 324332 112441 324360 113086
rect 324318 112432 324374 112441
rect 324318 112367 324374 112376
rect 324320 111784 324372 111790
rect 324318 111752 324320 111761
rect 324372 111752 324374 111761
rect 324318 111687 324374 111696
rect 324320 110424 324372 110430
rect 324320 110366 324372 110372
rect 324332 109449 324360 110366
rect 324318 109440 324374 109449
rect 324318 109375 324374 109384
rect 324320 108928 324372 108934
rect 324320 108870 324372 108876
rect 324332 108633 324360 108870
rect 324318 108624 324374 108633
rect 324318 108559 324374 108568
rect 325606 107808 325662 107817
rect 325712 107794 325740 214610
rect 325884 213308 325936 213314
rect 325884 213250 325936 213256
rect 325792 203720 325844 203726
rect 325792 203662 325844 203668
rect 325804 125497 325832 203662
rect 325896 156369 325924 213250
rect 327080 209092 327132 209098
rect 327080 209034 327132 209040
rect 325976 184272 326028 184278
rect 325976 184214 326028 184220
rect 325882 156360 325938 156369
rect 325882 156295 325938 156304
rect 325988 148850 326016 184214
rect 326068 176044 326120 176050
rect 326068 175986 326120 175992
rect 326080 173874 326108 175986
rect 326068 173868 326120 173874
rect 326068 173810 326120 173816
rect 325976 148844 326028 148850
rect 325976 148786 326028 148792
rect 325790 125488 325846 125497
rect 325790 125423 325846 125432
rect 325662 107766 325740 107794
rect 325606 107743 325662 107752
rect 323030 107128 323086 107137
rect 323030 107063 323086 107072
rect 322938 103184 322994 103193
rect 322938 103119 322994 103128
rect 321558 101144 321614 101153
rect 321558 101079 321614 101088
rect 321466 97336 321522 97345
rect 321466 97271 321522 97280
rect 321480 95198 321508 97271
rect 321468 95192 321520 95198
rect 321468 95134 321520 95140
rect 310520 86284 310572 86290
rect 310520 86226 310572 86232
rect 309876 83564 309928 83570
rect 309876 83506 309928 83512
rect 309784 4820 309836 4826
rect 309784 4762 309836 4768
rect 309046 4040 309102 4049
rect 309046 3975 309102 3984
rect 308588 3392 308640 3398
rect 307942 3360 307998 3369
rect 308588 3334 308640 3340
rect 307942 3295 307998 3304
rect 306748 2168 306800 2174
rect 306748 2110 306800 2116
rect 306760 480 306788 2110
rect 307956 480 307984 3295
rect 309060 480 309088 3975
rect 310532 3482 310560 86226
rect 317420 84856 317472 84862
rect 317420 84798 317472 84804
rect 315304 76628 315356 76634
rect 315304 76570 315356 76576
rect 311900 29776 311952 29782
rect 311900 29718 311952 29724
rect 311912 16574 311940 29718
rect 313278 18728 313334 18737
rect 313278 18663 313334 18672
rect 313292 16574 313320 18663
rect 311912 16546 312216 16574
rect 313292 16546 313872 16574
rect 311440 6316 311492 6322
rect 311440 6258 311492 6264
rect 310256 3454 310560 3482
rect 310256 480 310284 3454
rect 311452 480 311480 6258
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 354 312216 16546
rect 313844 480 313872 16546
rect 315316 4146 315344 76570
rect 317432 16574 317460 84798
rect 319444 83496 319496 83502
rect 319444 83438 319496 83444
rect 317432 16546 318104 16574
rect 317328 8968 317380 8974
rect 317328 8910 317380 8916
rect 315304 4140 315356 4146
rect 315304 4082 315356 4088
rect 316224 4140 316276 4146
rect 316224 4082 316276 4088
rect 315028 3392 315080 3398
rect 315028 3334 315080 3340
rect 315040 480 315068 3334
rect 316236 480 316264 4082
rect 317340 480 317368 8910
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 319456 3602 319484 83438
rect 321572 82822 321600 101079
rect 321650 98832 321706 98841
rect 321650 98767 321706 98776
rect 321664 93838 321692 98767
rect 321652 93832 321704 93838
rect 321652 93774 321704 93780
rect 323044 88330 323072 107063
rect 324320 106276 324372 106282
rect 324320 106218 324372 106224
rect 324332 105505 324360 106218
rect 324318 105496 324374 105505
rect 324318 105431 324374 105440
rect 324320 104848 324372 104854
rect 324318 104816 324320 104825
rect 324372 104816 324374 104825
rect 324318 104751 324374 104760
rect 327092 104718 327120 209034
rect 327172 206304 327224 206310
rect 327172 206246 327224 206252
rect 327184 127974 327212 206246
rect 327736 204921 327764 371214
rect 337396 276690 337424 616830
rect 347044 524476 347096 524482
rect 347044 524418 347096 524424
rect 347056 305658 347084 524418
rect 349160 358896 349212 358902
rect 349160 358838 349212 358844
rect 347044 305652 347096 305658
rect 347044 305594 347096 305600
rect 337384 276684 337436 276690
rect 337384 276626 337436 276632
rect 345664 269136 345716 269142
rect 345664 269078 345716 269084
rect 331864 264988 331916 264994
rect 331864 264930 331916 264936
rect 328552 232552 328604 232558
rect 328552 232494 328604 232500
rect 328460 228472 328512 228478
rect 328460 228414 328512 228420
rect 327722 204912 327778 204921
rect 327722 204847 327778 204856
rect 327264 203584 327316 203590
rect 327264 203526 327316 203532
rect 327276 136406 327304 203526
rect 327356 188352 327408 188358
rect 327356 188294 327408 188300
rect 327368 153338 327396 188294
rect 327356 153332 327408 153338
rect 327356 153274 327408 153280
rect 327264 136400 327316 136406
rect 327264 136342 327316 136348
rect 328472 128314 328500 228414
rect 328564 155854 328592 232494
rect 328644 204944 328696 204950
rect 328644 204886 328696 204892
rect 328552 155848 328604 155854
rect 328552 155790 328604 155796
rect 328656 129674 328684 204886
rect 328736 195288 328788 195294
rect 328736 195230 328788 195236
rect 328748 131034 328776 195230
rect 329932 194200 329984 194206
rect 329932 194142 329984 194148
rect 329944 164150 329972 194142
rect 331312 193996 331364 194002
rect 331312 193938 331364 193944
rect 331220 193860 331272 193866
rect 331220 193802 331272 193808
rect 330116 182844 330168 182850
rect 330116 182786 330168 182792
rect 330024 177336 330076 177342
rect 330024 177278 330076 177284
rect 329932 164144 329984 164150
rect 329932 164086 329984 164092
rect 330036 150414 330064 177278
rect 330024 150408 330076 150414
rect 330024 150350 330076 150356
rect 328736 131028 328788 131034
rect 328736 130970 328788 130976
rect 328644 129668 328696 129674
rect 328644 129610 328696 129616
rect 328460 128308 328512 128314
rect 328460 128250 328512 128256
rect 327172 127968 327224 127974
rect 327172 127910 327224 127916
rect 330128 121378 330156 182786
rect 330116 121372 330168 121378
rect 330116 121314 330168 121320
rect 331232 114442 331260 193802
rect 331324 160070 331352 193938
rect 331404 177404 331456 177410
rect 331404 177346 331456 177352
rect 331416 164218 331444 177346
rect 331404 164212 331456 164218
rect 331404 164154 331456 164160
rect 331312 160064 331364 160070
rect 331312 160006 331364 160012
rect 331220 114436 331272 114442
rect 331220 114378 331272 114384
rect 324320 104712 324372 104718
rect 324320 104654 324372 104660
rect 327080 104712 327132 104718
rect 327080 104654 327132 104660
rect 324332 104009 324360 104654
rect 324318 104000 324374 104009
rect 324318 103935 324374 103944
rect 324502 100872 324558 100881
rect 324502 100807 324558 100816
rect 324410 100192 324466 100201
rect 324410 100127 324466 100136
rect 324424 92449 324452 100127
rect 324410 92440 324466 92449
rect 324410 92375 324466 92384
rect 324516 91089 324544 100807
rect 324594 97064 324650 97073
rect 324594 96999 324650 97008
rect 324608 92478 324636 96999
rect 324596 92472 324648 92478
rect 324596 92414 324648 92420
rect 324502 91080 324558 91089
rect 324502 91015 324558 91024
rect 323032 88324 323084 88330
rect 323032 88266 323084 88272
rect 324320 83564 324372 83570
rect 324320 83506 324372 83512
rect 321560 82816 321612 82822
rect 321560 82758 321612 82764
rect 322940 80708 322992 80714
rect 322940 80650 322992 80656
rect 321558 73808 321614 73817
rect 321558 73743 321614 73752
rect 321572 16574 321600 73743
rect 321572 16546 322152 16574
rect 320916 4820 320968 4826
rect 320916 4762 320968 4768
rect 319444 3596 319496 3602
rect 319444 3538 319496 3544
rect 319720 3528 319772 3534
rect 319720 3470 319772 3476
rect 319732 480 319760 3470
rect 320928 480 320956 4762
rect 322124 480 322152 16546
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 322952 354 322980 80650
rect 324332 3482 324360 83506
rect 328460 79348 328512 79354
rect 328460 79290 328512 79296
rect 324412 24268 324464 24274
rect 324412 24210 324464 24216
rect 324424 3602 324452 24210
rect 328472 16574 328500 79290
rect 328472 16546 328776 16574
rect 328000 14612 328052 14618
rect 328000 14554 328052 14560
rect 324412 3596 324464 3602
rect 324412 3538 324464 3544
rect 325608 3596 325660 3602
rect 325608 3538 325660 3544
rect 324332 3454 324452 3482
rect 324424 480 324452 3454
rect 325620 480 325648 3538
rect 326804 3460 326856 3466
rect 326804 3402 326856 3408
rect 326816 480 326844 3402
rect 328012 480 328040 14554
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 328748 354 328776 16546
rect 331218 13016 331274 13025
rect 331218 12951 331274 12960
rect 330392 3460 330444 3466
rect 330392 3402 330444 3408
rect 330404 480 330432 3402
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331232 354 331260 12951
rect 331876 8294 331904 264930
rect 340880 257372 340932 257378
rect 340880 257314 340932 257320
rect 335360 253972 335412 253978
rect 335360 253914 335412 253920
rect 333980 231124 334032 231130
rect 333980 231066 334032 231072
rect 332600 211812 332652 211818
rect 332600 211754 332652 211760
rect 332612 110430 332640 211754
rect 332784 181620 332836 181626
rect 332784 181562 332836 181568
rect 332690 181384 332746 181393
rect 332690 181319 332746 181328
rect 332704 114510 332732 181319
rect 332796 161362 332824 181562
rect 332876 177472 332928 177478
rect 332876 177414 332928 177420
rect 332888 162790 332916 177414
rect 332876 162784 332928 162790
rect 332876 162726 332928 162732
rect 332784 161356 332836 161362
rect 332784 161298 332836 161304
rect 332692 114504 332744 114510
rect 332692 114446 332744 114452
rect 332600 110424 332652 110430
rect 332600 110366 332652 110372
rect 332600 51808 332652 51814
rect 332600 51750 332652 51756
rect 332612 16574 332640 51750
rect 333992 16574 334020 231066
rect 334164 196648 334216 196654
rect 334164 196590 334216 196596
rect 334072 182980 334124 182986
rect 334072 182922 334124 182928
rect 334084 118590 334112 182922
rect 334176 168366 334204 196590
rect 334256 184408 334308 184414
rect 334256 184350 334308 184356
rect 334164 168360 334216 168366
rect 334164 168302 334216 168308
rect 334268 158642 334296 184350
rect 334256 158636 334308 158642
rect 334256 158578 334308 158584
rect 334072 118584 334124 118590
rect 334072 118526 334124 118532
rect 335372 16574 335400 253914
rect 336740 225684 336792 225690
rect 336740 225626 336792 225632
rect 335452 180192 335504 180198
rect 335452 180134 335504 180140
rect 335464 117230 335492 180134
rect 335544 178832 335596 178838
rect 335544 178774 335596 178780
rect 335556 137902 335584 178774
rect 335636 175976 335688 175982
rect 335636 175918 335688 175924
rect 335648 165578 335676 175918
rect 335636 165572 335688 165578
rect 335636 165514 335688 165520
rect 336752 142050 336780 225626
rect 338120 215960 338172 215966
rect 338120 215902 338172 215908
rect 336832 195356 336884 195362
rect 336832 195298 336884 195304
rect 336740 142044 336792 142050
rect 336740 141986 336792 141992
rect 335544 137896 335596 137902
rect 335544 137838 335596 137844
rect 336844 118658 336872 195298
rect 337016 185632 337068 185638
rect 337016 185574 337068 185580
rect 336922 178664 336978 178673
rect 336922 178599 336978 178608
rect 336936 143478 336964 178599
rect 337028 169726 337056 185574
rect 337016 169720 337068 169726
rect 337016 169662 337068 169668
rect 336924 143472 336976 143478
rect 336924 143414 336976 143420
rect 336832 118652 336884 118658
rect 336832 118594 336884 118600
rect 335452 117224 335504 117230
rect 335452 117166 335504 117172
rect 338132 113150 338160 215902
rect 339684 207732 339736 207738
rect 339684 207674 339736 207680
rect 339500 205148 339552 205154
rect 339500 205090 339552 205096
rect 338212 191276 338264 191282
rect 338212 191218 338264 191224
rect 338224 120086 338252 191218
rect 338304 182912 338356 182918
rect 338304 182854 338356 182860
rect 338316 140758 338344 182854
rect 338394 175944 338450 175953
rect 338394 175879 338450 175888
rect 338408 155922 338436 175879
rect 338396 155916 338448 155922
rect 338396 155858 338448 155864
rect 338304 140752 338356 140758
rect 338304 140694 338356 140700
rect 338212 120080 338264 120086
rect 338212 120022 338264 120028
rect 338120 113144 338172 113150
rect 338120 113086 338172 113092
rect 339512 111790 339540 205090
rect 339592 178900 339644 178906
rect 339592 178842 339644 178848
rect 339500 111784 339552 111790
rect 339500 111726 339552 111732
rect 339604 108934 339632 178842
rect 339696 139398 339724 207674
rect 339776 188556 339828 188562
rect 339776 188498 339828 188504
rect 339788 157282 339816 188498
rect 339776 157276 339828 157282
rect 339776 157218 339828 157224
rect 339684 139392 339736 139398
rect 339684 139334 339736 139340
rect 339592 108928 339644 108934
rect 339592 108870 339644 108876
rect 336738 53136 336794 53145
rect 336738 53071 336794 53080
rect 336752 16574 336780 53071
rect 339498 22672 339554 22681
rect 339498 22607 339554 22616
rect 332612 16546 332732 16574
rect 333992 16546 334664 16574
rect 335372 16546 336320 16574
rect 336752 16546 337056 16574
rect 331864 8288 331916 8294
rect 331864 8230 331916 8236
rect 332704 480 332732 16546
rect 333888 8288 333940 8294
rect 333888 8230 333940 8236
rect 333900 480 333928 8230
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 16546
rect 336292 480 336320 16546
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337028 354 337056 16546
rect 338672 3596 338724 3602
rect 338672 3538 338724 3544
rect 338684 480 338712 3538
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339512 354 339540 22607
rect 340892 16574 340920 257314
rect 345020 222896 345072 222902
rect 345020 222838 345072 222844
rect 343640 218816 343692 218822
rect 343640 218758 343692 218764
rect 342260 207664 342312 207670
rect 342260 207606 342312 207612
rect 341064 192500 341116 192506
rect 341064 192442 341116 192448
rect 340972 189780 341024 189786
rect 340972 189722 341024 189728
rect 340984 124166 341012 189722
rect 341076 136610 341104 192442
rect 341156 181552 341208 181558
rect 341156 181494 341208 181500
rect 341168 158710 341196 181494
rect 341156 158704 341208 158710
rect 341156 158646 341208 158652
rect 341064 136604 341116 136610
rect 341064 136546 341116 136552
rect 340972 124160 341024 124166
rect 340972 124102 341024 124108
rect 342272 16574 342300 207606
rect 342444 203788 342496 203794
rect 342444 203730 342496 203736
rect 342352 199504 342404 199510
rect 342352 199446 342404 199452
rect 342364 125594 342392 199446
rect 342456 144906 342484 203730
rect 342536 181484 342588 181490
rect 342536 181426 342588 181432
rect 342548 162858 342576 181426
rect 342536 162852 342588 162858
rect 342536 162794 342588 162800
rect 342444 144900 342496 144906
rect 342444 144842 342496 144848
rect 342352 125588 342404 125594
rect 342352 125530 342404 125536
rect 343652 117298 343680 218758
rect 343732 202224 343784 202230
rect 343732 202166 343784 202172
rect 343744 143546 343772 202166
rect 343824 191140 343876 191146
rect 343824 191082 343876 191088
rect 343836 147626 343864 191082
rect 343916 178696 343968 178702
rect 343916 178638 343968 178644
rect 343824 147620 343876 147626
rect 343824 147562 343876 147568
rect 343732 143540 343784 143546
rect 343732 143482 343784 143488
rect 343928 137970 343956 178638
rect 343916 137964 343968 137970
rect 343916 137906 343968 137912
rect 345032 121446 345060 222838
rect 345112 216096 345164 216102
rect 345112 216038 345164 216044
rect 345020 121440 345072 121446
rect 345020 121382 345072 121388
rect 343640 117292 343692 117298
rect 343640 117234 343692 117240
rect 345124 115938 345152 216038
rect 345204 180124 345256 180130
rect 345204 180066 345256 180072
rect 345216 142118 345244 180066
rect 345204 142112 345256 142118
rect 345204 142054 345256 142060
rect 345112 115932 345164 115938
rect 345112 115874 345164 115880
rect 343640 33924 343692 33930
rect 343640 33866 343692 33872
rect 343652 16574 343680 33866
rect 340892 16546 341012 16574
rect 342272 16546 342944 16574
rect 343652 16546 344600 16574
rect 340984 480 341012 16546
rect 342166 3496 342222 3505
rect 342166 3431 342222 3440
rect 342180 480 342208 3431
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 16546
rect 344572 480 344600 16546
rect 345676 4214 345704 269078
rect 346492 220244 346544 220250
rect 346492 220186 346544 220192
rect 346400 191208 346452 191214
rect 346400 191150 346452 191156
rect 346412 16574 346440 191150
rect 346504 161430 346532 220186
rect 347780 206372 347832 206378
rect 347780 206314 347832 206320
rect 346584 185836 346636 185842
rect 346584 185778 346636 185784
rect 346492 161424 346544 161430
rect 346492 161366 346544 161372
rect 346596 151774 346624 185778
rect 346676 184204 346728 184210
rect 346676 184146 346728 184152
rect 346688 154562 346716 184146
rect 346676 154556 346728 154562
rect 346676 154498 346728 154504
rect 346584 151768 346636 151774
rect 346584 151710 346636 151716
rect 347792 106282 347820 206314
rect 347872 195424 347924 195430
rect 347872 195366 347924 195372
rect 347884 132462 347912 195366
rect 347872 132456 347924 132462
rect 347872 132398 347924 132404
rect 347780 106276 347832 106282
rect 347780 106218 347832 106224
rect 346412 16546 346992 16574
rect 345664 4208 345716 4214
rect 345664 4150 345716 4156
rect 345756 3528 345808 3534
rect 345756 3470 345808 3476
rect 345768 480 345796 3470
rect 346964 480 346992 16546
rect 348056 4004 348108 4010
rect 348056 3946 348108 3952
rect 348068 480 348096 3946
rect 349172 3602 349200 358838
rect 349252 357876 349304 357882
rect 349252 357818 349304 357824
rect 349264 6914 349292 357818
rect 355324 324352 355376 324358
rect 355324 324294 355376 324300
rect 350540 318844 350592 318850
rect 350540 318786 350592 318792
rect 349344 196784 349396 196790
rect 349344 196726 349396 196732
rect 349356 122806 349384 196726
rect 349436 188420 349488 188426
rect 349436 188362 349488 188368
rect 349448 148986 349476 188362
rect 349436 148980 349488 148986
rect 349436 148922 349488 148928
rect 349344 122800 349396 122806
rect 349344 122742 349396 122748
rect 349344 21548 349396 21554
rect 349344 21490 349396 21496
rect 349356 16574 349384 21490
rect 350552 16574 350580 318786
rect 355336 283626 355364 324294
rect 355324 283620 355376 283626
rect 355324 283562 355376 283568
rect 353944 281580 353996 281586
rect 353944 281522 353996 281528
rect 351920 221468 351972 221474
rect 351920 221410 351972 221416
rect 350632 184476 350684 184482
rect 350632 184418 350684 184424
rect 350644 131102 350672 184418
rect 350632 131096 350684 131102
rect 350632 131038 350684 131044
rect 351932 129742 351960 221410
rect 351920 129736 351972 129742
rect 351920 129678 351972 129684
rect 353956 60722 353984 281522
rect 364352 237250 364380 702406
rect 397472 698970 397500 703520
rect 397460 698964 397512 698970
rect 397460 698906 397512 698912
rect 400864 510672 400916 510678
rect 400864 510614 400916 510620
rect 373264 360256 373316 360262
rect 373264 360198 373316 360204
rect 364340 237244 364392 237250
rect 364340 237186 364392 237192
rect 356060 217388 356112 217394
rect 356060 217330 356112 217336
rect 354680 202292 354732 202298
rect 354680 202234 354732 202240
rect 353944 60716 353996 60722
rect 353944 60658 353996 60664
rect 349356 16546 349476 16574
rect 350552 16546 351224 16574
rect 349264 6886 349384 6914
rect 349356 3602 349384 6886
rect 349160 3596 349212 3602
rect 349160 3538 349212 3544
rect 349344 3596 349396 3602
rect 349344 3538 349396 3544
rect 349448 3482 349476 16546
rect 350448 4208 350500 4214
rect 350448 4150 350500 4156
rect 349264 3454 349476 3482
rect 349264 480 349292 3454
rect 350460 480 350488 4150
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 354692 4010 354720 202234
rect 356072 104854 356100 217330
rect 373276 179382 373304 360198
rect 374644 330540 374696 330546
rect 374644 330482 374696 330488
rect 374656 303618 374684 330482
rect 374644 303612 374696 303618
rect 374644 303554 374696 303560
rect 400876 290494 400904 510614
rect 412652 330546 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 429856 700330 429884 703520
rect 462332 702642 462360 703520
rect 462320 702636 462372 702642
rect 462320 702578 462372 702584
rect 478524 702574 478552 703520
rect 494808 702710 494836 703520
rect 494796 702704 494848 702710
rect 494796 702646 494848 702652
rect 478512 702568 478564 702574
rect 478512 702510 478564 702516
rect 429844 700324 429896 700330
rect 429844 700266 429896 700272
rect 527192 699718 527220 703520
rect 543476 702545 543504 703520
rect 543462 702536 543518 702545
rect 559668 702506 559696 703520
rect 580354 702672 580410 702681
rect 580354 702607 580410 702616
rect 543462 702471 543518 702480
rect 559656 702500 559708 702506
rect 559656 702442 559708 702448
rect 525064 699712 525116 699718
rect 525064 699654 525116 699660
rect 527180 699712 527232 699718
rect 527180 699654 527232 699660
rect 449164 354748 449216 354754
rect 449164 354690 449216 354696
rect 412640 330540 412692 330546
rect 412640 330482 412692 330488
rect 418804 313948 418856 313954
rect 418804 313890 418856 313896
rect 400864 290488 400916 290494
rect 400864 290430 400916 290436
rect 395344 242956 395396 242962
rect 395344 242898 395396 242904
rect 395356 233102 395384 242898
rect 395344 233096 395396 233102
rect 395344 233038 395396 233044
rect 373264 179376 373316 179382
rect 373264 179318 373316 179324
rect 356060 104848 356112 104854
rect 356060 104790 356112 104796
rect 378784 89004 378836 89010
rect 378784 88946 378836 88952
rect 356702 61432 356758 61441
rect 356702 61367 356758 61376
rect 354680 4004 354732 4010
rect 354680 3946 354732 3952
rect 356716 3466 356744 61367
rect 378796 20670 378824 88946
rect 418816 73166 418844 313890
rect 449176 126954 449204 354690
rect 472624 345092 472676 345098
rect 472624 345034 472676 345040
rect 468484 316736 468536 316742
rect 468484 316678 468536 316684
rect 467104 245676 467156 245682
rect 467104 245618 467156 245624
rect 449164 126948 449216 126954
rect 449164 126890 449216 126896
rect 467116 100706 467144 245618
rect 468496 113150 468524 316678
rect 471244 309800 471296 309806
rect 471244 309742 471296 309748
rect 471256 219434 471284 309742
rect 471244 219428 471296 219434
rect 471244 219370 471296 219376
rect 472636 139398 472664 345034
rect 525076 238814 525104 699654
rect 580368 697241 580396 702607
rect 580354 697232 580410 697241
rect 580354 697167 580410 697176
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580262 670712 580318 670721
rect 580262 670647 580318 670656
rect 579986 630864 580042 630873
rect 579986 630799 580042 630808
rect 580000 630698 580028 630799
rect 579988 630692 580040 630698
rect 579988 630634 580040 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580184 590714 580212 590951
rect 580172 590708 580224 590714
rect 580172 590650 580224 590656
rect 579894 564360 579950 564369
rect 579894 564295 579950 564304
rect 579908 563106 579936 564295
rect 579896 563100 579948 563106
rect 579896 563042 579948 563048
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 580184 470626 580212 471407
rect 580172 470620 580224 470626
rect 580172 470562 580224 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 579986 404968 580042 404977
rect 579986 404903 580042 404912
rect 580000 404394 580028 404903
rect 579988 404388 580040 404394
rect 579988 404330 580040 404336
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 580276 374678 580304 670647
rect 582378 644056 582434 644065
rect 582378 643991 582434 644000
rect 580354 577688 580410 577697
rect 580354 577623 580410 577632
rect 580264 374672 580316 374678
rect 580264 374614 580316 374620
rect 580368 370530 580396 577623
rect 580356 370524 580408 370530
rect 580356 370466 580408 370472
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580184 364410 580212 365055
rect 580172 364404 580224 364410
rect 580172 364346 580224 364352
rect 580264 362976 580316 362982
rect 580264 362918 580316 362924
rect 580276 351937 580304 362918
rect 580356 354000 580408 354006
rect 580356 353942 580408 353948
rect 580262 351928 580318 351937
rect 580262 351863 580318 351872
rect 580264 351212 580316 351218
rect 580264 351154 580316 351160
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 324358 580212 325207
rect 580172 324352 580224 324358
rect 580172 324294 580224 324300
rect 579620 299464 579672 299470
rect 579620 299406 579672 299412
rect 579632 298761 579660 299406
rect 579618 298752 579674 298761
rect 579618 298687 579674 298696
rect 579620 259412 579672 259418
rect 579620 259354 579672 259360
rect 579632 258913 579660 259354
rect 579618 258904 579674 258913
rect 579618 258839 579674 258848
rect 579894 245576 579950 245585
rect 579894 245511 579950 245520
rect 579908 244322 579936 245511
rect 574744 244316 574796 244322
rect 574744 244258 574796 244264
rect 579896 244316 579948 244322
rect 579896 244258 579948 244264
rect 525064 238808 525116 238814
rect 525064 238750 525116 238756
rect 574756 223582 574784 244258
rect 579620 233096 579672 233102
rect 579620 233038 579672 233044
rect 579632 232393 579660 233038
rect 579618 232384 579674 232393
rect 579618 232319 579674 232328
rect 574744 223576 574796 223582
rect 574744 223518 574796 223524
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580276 165889 580304 351154
rect 580368 312089 580396 353942
rect 580354 312080 580410 312089
rect 580354 312015 580410 312024
rect 580354 272232 580410 272241
rect 580354 272167 580410 272176
rect 580368 237386 580396 272167
rect 580356 237380 580408 237386
rect 580356 237322 580408 237328
rect 582392 233170 582420 643991
rect 582470 537840 582526 537849
rect 582470 537775 582526 537784
rect 582484 238678 582512 537775
rect 582562 431624 582618 431633
rect 582562 431559 582618 431568
rect 582576 238746 582604 431559
rect 582654 418296 582710 418305
rect 582654 418231 582710 418240
rect 582564 238740 582616 238746
rect 582564 238682 582616 238688
rect 582472 238672 582524 238678
rect 582472 238614 582524 238620
rect 582668 233238 582696 418231
rect 582656 233232 582708 233238
rect 582656 233174 582708 233180
rect 582380 233164 582432 233170
rect 582380 233106 582432 233112
rect 582380 228404 582432 228410
rect 582380 228346 582432 228352
rect 580356 224256 580408 224262
rect 580356 224198 580408 224204
rect 580262 165880 580318 165889
rect 580262 165815 580318 165824
rect 580368 152697 580396 224198
rect 580448 220108 580500 220114
rect 580448 220050 580500 220056
rect 580460 192545 580488 220050
rect 582392 205737 582420 228346
rect 582472 218748 582524 218754
rect 582472 218690 582524 218696
rect 582378 205728 582434 205737
rect 582378 205663 582434 205672
rect 582380 199436 582432 199442
rect 582380 199378 582432 199384
rect 580446 192536 580502 192545
rect 580446 192471 580502 192480
rect 580354 152688 580410 152697
rect 580354 152623 580410 152632
rect 472624 139392 472676 139398
rect 580172 139392 580224 139398
rect 472624 139334 472676 139340
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 468484 113144 468536 113150
rect 468484 113086 468536 113092
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 467104 100700 467156 100706
rect 467104 100642 467156 100648
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 418804 73160 418856 73166
rect 418804 73102 418856 73108
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580170 47560 580226 47569
rect 580170 47495 580226 47504
rect 580184 46345 580212 47495
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 378784 20664 378836 20670
rect 378784 20606 378836 20612
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 582392 6633 582420 199378
rect 582484 33153 582512 218690
rect 582470 33144 582526 33153
rect 582470 33079 582526 33088
rect 582378 6624 582434 6633
rect 582378 6559 582434 6568
rect 356704 3460 356756 3466
rect 356704 3402 356756 3408
rect 579804 3460 579856 3466
rect 579804 3402 579856 3408
rect 579816 480 579844 3402
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 2778 658144 2834 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3422 606076 3478 606112
rect 3422 606056 3424 606076
rect 3424 606056 3476 606076
rect 3476 606056 3478 606076
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3422 553832 3478 553888
rect 3422 527856 3478 527912
rect 3422 501744 3478 501800
rect 3054 475632 3110 475688
rect 3146 449520 3202 449576
rect 2870 410488 2926 410544
rect 3054 358400 3110 358456
rect 3330 345344 3386 345400
rect 3514 462576 3570 462632
rect 3514 423544 3570 423600
rect 3514 397468 3516 397488
rect 3516 397468 3568 397488
rect 3568 397468 3570 397488
rect 3514 397432 3570 397468
rect 3514 371320 3570 371376
rect 3422 319232 3478 319288
rect 3238 306176 3294 306232
rect 3330 293120 3386 293176
rect 3054 267144 3110 267200
rect 2778 254108 2834 254144
rect 2778 254088 2780 254108
rect 2780 254088 2832 254108
rect 2832 254088 2834 254108
rect 3330 241032 3386 241088
rect 3330 214920 3386 214976
rect 3146 188808 3202 188864
rect 3146 110608 3202 110664
rect 2778 97552 2834 97608
rect 3146 84632 3202 84688
rect 3606 201864 3662 201920
rect 3514 162832 3570 162888
rect 3514 149776 3570 149832
rect 3514 136720 3570 136776
rect 3422 71576 3478 71632
rect 3054 58520 3110 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3514 32408 3570 32464
rect 3422 19352 3478 19408
rect 21362 266328 21418 266384
rect 9678 46144 9734 46200
rect 3422 6432 3478 6488
rect 12438 18536 12494 18592
rect 22098 17176 22154 17232
rect 35806 293936 35862 293992
rect 53562 211792 53618 211848
rect 52366 210432 52422 210488
rect 57886 298696 57942 298752
rect 54942 213152 54998 213208
rect 53746 179968 53802 180024
rect 57794 190984 57850 191040
rect 62302 271904 62358 271960
rect 60646 189624 60702 189680
rect 64602 225528 64658 225584
rect 67270 261840 67326 261896
rect 68742 296792 68798 296848
rect 67730 291080 67786 291136
rect 67638 290400 67694 290456
rect 67638 289040 67694 289096
rect 68374 288360 68430 288416
rect 67638 287680 67694 287736
rect 67730 287000 67786 287056
rect 67546 286320 67602 286376
rect 67638 285676 67640 285696
rect 67640 285676 67692 285696
rect 67692 285676 67694 285696
rect 67638 285640 67694 285676
rect 68282 284280 68338 284336
rect 67638 282920 67694 282976
rect 67638 281560 67694 281616
rect 67730 280880 67786 280936
rect 67638 280236 67640 280256
rect 67640 280236 67692 280256
rect 67692 280236 67694 280256
rect 67638 280200 67694 280236
rect 67914 279520 67970 279576
rect 67730 278160 67786 278216
rect 67638 277500 67694 277536
rect 67638 277480 67640 277500
rect 67640 277480 67692 277500
rect 67692 277480 67694 277500
rect 67730 276800 67786 276856
rect 67638 276140 67694 276176
rect 67638 276120 67640 276140
rect 67640 276120 67692 276140
rect 67692 276120 67694 276140
rect 67638 274760 67694 274816
rect 67730 274080 67786 274136
rect 67638 273400 67694 273456
rect 67730 272720 67786 272776
rect 67638 272040 67694 272096
rect 67638 271360 67694 271416
rect 67730 270680 67786 270736
rect 67638 270000 67694 270056
rect 68190 269320 68246 269376
rect 68190 268640 68246 268696
rect 67638 267960 67694 268016
rect 67638 266600 67694 266656
rect 67638 265920 67694 265976
rect 67730 265240 67786 265296
rect 67730 264560 67786 264616
rect 67638 263880 67694 263936
rect 67730 263200 67786 263256
rect 67638 262520 67694 262576
rect 67638 260480 67694 260536
rect 68098 259800 68154 259856
rect 67730 259120 67786 259176
rect 67638 258440 67694 258496
rect 67638 257080 67694 257136
rect 67638 256400 67694 256456
rect 67730 255040 67786 255096
rect 67638 254360 67694 254416
rect 67638 253680 67694 253736
rect 67638 253000 67694 253056
rect 67638 252320 67694 252376
rect 67546 251640 67602 251696
rect 55126 178608 55182 178664
rect 66074 129240 66130 129296
rect 66166 126248 66222 126304
rect 65522 125160 65578 125216
rect 66074 123528 66130 123584
rect 66074 122576 66130 122632
rect 63314 90888 63370 90944
rect 66074 102312 66130 102368
rect 67454 120808 67510 120864
rect 66166 94832 66222 94888
rect 68558 284960 68614 285016
rect 68466 283600 68522 283656
rect 68834 279520 68890 279576
rect 68926 275440 68982 275496
rect 68374 261160 68430 261216
rect 68282 257216 68338 257272
rect 68834 255720 68890 255776
rect 68742 250960 68798 251016
rect 67638 250280 67694 250336
rect 67822 248920 67878 248976
rect 67730 248240 67786 248296
rect 67638 247560 67694 247616
rect 68650 246200 68706 246256
rect 67638 245520 67694 245576
rect 67730 242120 67786 242176
rect 67638 241460 67694 241496
rect 67638 241440 67640 241460
rect 67640 241440 67692 241460
rect 67692 241440 67694 241460
rect 68742 233824 68798 233880
rect 69018 257760 69074 257816
rect 69110 244840 69166 244896
rect 68926 244160 68982 244216
rect 68834 214512 68890 214568
rect 71686 292304 71742 292360
rect 73894 292848 73950 292904
rect 76102 300872 76158 300928
rect 77758 292712 77814 292768
rect 78402 292576 78458 292632
rect 84382 299512 84438 299568
rect 89350 298152 89406 298208
rect 95146 295976 95202 296032
rect 96434 294072 96490 294128
rect 95790 293936 95846 293992
rect 104898 297336 104954 297392
rect 104898 295976 104954 296032
rect 106094 295296 106150 295352
rect 108026 294208 108082 294264
rect 114558 358808 114614 358864
rect 114466 294072 114522 294128
rect 117778 291896 117834 291952
rect 120170 286320 120226 286376
rect 120078 268640 120134 268696
rect 69202 243480 69258 243536
rect 120170 250960 120226 251016
rect 120630 250960 120686 251016
rect 119802 242528 119858 242584
rect 69846 240760 69902 240816
rect 74538 197920 74594 197976
rect 73158 184184 73214 184240
rect 77298 215872 77354 215928
rect 75182 181328 75238 181384
rect 82910 238720 82966 238776
rect 80058 186904 80114 186960
rect 84382 210296 84438 210352
rect 95698 237224 95754 237280
rect 96526 237224 96582 237280
rect 105450 238040 105506 238096
rect 106738 237088 106794 237144
rect 100758 188264 100814 188320
rect 98642 182824 98698 182880
rect 110418 206216 110474 206272
rect 117042 239808 117098 239864
rect 117962 236544 118018 236600
rect 120078 241440 120134 241496
rect 117962 200640 118018 200696
rect 100666 177520 100722 177576
rect 102046 177520 102102 177576
rect 106186 177520 106242 177576
rect 107566 177520 107622 177576
rect 97814 176840 97870 176896
rect 112994 177520 113050 177576
rect 114466 177520 114522 177576
rect 116950 177520 117006 177576
rect 118606 177520 118662 177576
rect 110694 177112 110750 177168
rect 113914 177112 113970 177168
rect 121550 291760 121606 291816
rect 121642 291080 121698 291136
rect 121550 290400 121606 290456
rect 121550 289756 121552 289776
rect 121552 289756 121604 289776
rect 121604 289756 121606 289776
rect 121550 289720 121606 289756
rect 121550 289040 121606 289096
rect 121734 288360 121790 288416
rect 121642 287680 121698 287736
rect 121458 285640 121514 285696
rect 121458 284960 121514 285016
rect 121550 284280 121606 284336
rect 121458 283600 121514 283656
rect 121550 282240 121606 282296
rect 121458 281580 121514 281616
rect 121458 281560 121460 281580
rect 121460 281560 121512 281580
rect 121512 281560 121514 281580
rect 121550 280880 121606 280936
rect 121458 280220 121514 280256
rect 121458 280200 121460 280220
rect 121460 280200 121512 280220
rect 121512 280200 121514 280220
rect 121458 278840 121514 278896
rect 121458 277480 121514 277536
rect 121550 276800 121606 276856
rect 121458 276120 121514 276176
rect 121550 275440 121606 275496
rect 121458 274780 121514 274816
rect 121458 274760 121460 274780
rect 121460 274760 121512 274780
rect 121512 274760 121514 274780
rect 121458 274080 121514 274136
rect 121458 273400 121514 273456
rect 122746 287000 122802 287056
rect 121734 282920 121790 282976
rect 122286 279520 122342 279576
rect 122194 278160 122250 278216
rect 121642 272720 121698 272776
rect 122102 272720 122158 272776
rect 121458 272040 121514 272096
rect 121458 271360 121514 271416
rect 121550 270000 121606 270056
rect 121458 269320 121514 269376
rect 121458 267960 121514 268016
rect 121550 267280 121606 267336
rect 121458 266600 121514 266656
rect 121550 265920 121606 265976
rect 121458 265240 121514 265296
rect 121550 263880 121606 263936
rect 121458 263200 121514 263256
rect 121458 262520 121514 262576
rect 121642 261840 121698 261896
rect 121550 261160 121606 261216
rect 121458 260480 121514 260536
rect 121458 259800 121514 259856
rect 121458 259120 121514 259176
rect 121550 257760 121606 257816
rect 121458 257080 121514 257136
rect 120998 255856 121054 255912
rect 120998 255312 121054 255368
rect 122102 255040 122158 255096
rect 121458 254360 121514 254416
rect 121550 253680 121606 253736
rect 121458 253000 121514 253056
rect 121458 251640 121514 251696
rect 121458 250280 121514 250336
rect 121550 249600 121606 249656
rect 121458 248920 121514 248976
rect 121458 248240 121514 248296
rect 121550 247968 121606 248024
rect 121550 246880 121606 246936
rect 121458 246200 121514 246256
rect 121550 245520 121606 245576
rect 121458 244840 121514 244896
rect 121550 244160 121606 244216
rect 121458 243480 121514 243536
rect 121458 242820 121514 242856
rect 121458 242800 121460 242820
rect 121460 242800 121512 242820
rect 121512 242800 121514 242820
rect 121550 242120 121606 242176
rect 121458 240760 121514 240816
rect 121550 240080 121606 240136
rect 122194 237904 122250 237960
rect 125138 292712 125194 292768
rect 125138 284144 125194 284200
rect 127806 177520 127862 177576
rect 131854 298152 131910 298208
rect 134706 199280 134762 199336
rect 130474 181464 130530 181520
rect 138018 235864 138074 235920
rect 137374 192480 137430 192536
rect 141514 294072 141570 294128
rect 150346 357856 150402 357912
rect 144366 241168 144422 241224
rect 145746 206352 145802 206408
rect 155406 300872 155462 300928
rect 152554 289176 152610 289232
rect 154026 299512 154082 299568
rect 154026 240760 154082 240816
rect 154118 192616 154174 192672
rect 129462 177520 129518 177576
rect 133786 177520 133842 177576
rect 108118 176704 108174 176760
rect 109866 176704 109922 176760
rect 119710 176704 119766 176760
rect 122010 176704 122066 176760
rect 123022 176704 123078 176760
rect 124954 176704 125010 176760
rect 125874 176704 125930 176760
rect 128266 176704 128322 176760
rect 132038 176704 132094 176760
rect 134430 176724 134486 176760
rect 134430 176704 134432 176724
rect 134432 176704 134484 176724
rect 134484 176704 134486 176724
rect 135718 176704 135774 176760
rect 148230 176704 148286 176760
rect 104622 175480 104678 175536
rect 157338 297336 157394 297392
rect 160742 356088 160798 356144
rect 162122 354864 162178 354920
rect 160834 291896 160890 291952
rect 158534 196560 158590 196616
rect 161386 184320 161442 184376
rect 163594 221448 163650 221504
rect 158994 176740 158996 176760
rect 158996 176740 159048 176760
rect 159048 176740 159050 176760
rect 158994 176704 159050 176740
rect 166446 298696 166502 298752
rect 166262 211928 166318 211984
rect 155222 175888 155278 175944
rect 120814 175480 120870 175536
rect 130750 175480 130806 175536
rect 115754 174936 115810 174992
rect 67638 128016 67694 128072
rect 67730 100680 67786 100736
rect 67638 93744 67694 93800
rect 67546 91024 67602 91080
rect 165526 174528 165582 174584
rect 169114 176976 169170 177032
rect 168010 171536 168066 171592
rect 170494 175344 170550 175400
rect 102046 94696 102102 94752
rect 113730 94696 113786 94752
rect 115478 94696 115534 94752
rect 133142 94696 133198 94752
rect 134430 93608 134486 93664
rect 151726 93608 151782 93664
rect 110142 93472 110198 93528
rect 118054 93472 118110 93528
rect 119526 93472 119582 93528
rect 128174 93200 128230 93256
rect 74814 92384 74870 92440
rect 85762 92384 85818 92440
rect 88062 92384 88118 92440
rect 88982 92420 88984 92440
rect 88984 92420 89036 92440
rect 89036 92420 89038 92440
rect 88982 92384 89038 92420
rect 100574 92384 100630 92440
rect 109222 92384 109278 92440
rect 112166 92384 112222 92440
rect 115478 92384 115534 92440
rect 116766 92384 116822 92440
rect 119710 92384 119766 92440
rect 125874 92384 125930 92440
rect 126518 92384 126574 92440
rect 85486 91160 85542 91216
rect 49698 62736 49754 62792
rect 56598 55800 56654 55856
rect 62118 44784 62174 44840
rect 66258 25472 66314 25528
rect 52550 4800 52606 4856
rect 99194 91432 99250 91488
rect 95054 91296 95110 91352
rect 97262 91296 97318 91352
rect 99102 91296 99158 91352
rect 86866 91160 86922 91216
rect 91006 91160 91062 91216
rect 92386 91160 92442 91216
rect 93766 91160 93822 91216
rect 95146 91160 95202 91216
rect 96158 91160 96214 91216
rect 96158 86808 96214 86864
rect 97906 91160 97962 91216
rect 99286 91160 99342 91216
rect 100482 91160 100538 91216
rect 101862 91568 101918 91624
rect 99286 78376 99342 78432
rect 107014 91296 107070 91352
rect 102046 91160 102102 91216
rect 103426 91160 103482 91216
rect 104346 91160 104402 91216
rect 104622 91160 104678 91216
rect 105726 91160 105782 91216
rect 106186 91160 106242 91216
rect 107566 91160 107622 91216
rect 107842 91160 107898 91216
rect 108946 91160 109002 91216
rect 107014 86672 107070 86728
rect 106186 84088 106242 84144
rect 110326 91160 110382 91216
rect 110970 91160 111026 91216
rect 110970 88168 111026 88224
rect 111430 91160 111486 91216
rect 113086 91160 113142 91216
rect 114466 91160 114522 91216
rect 122838 91432 122894 91488
rect 122102 91296 122158 91352
rect 115846 91160 115902 91216
rect 117226 91160 117282 91216
rect 118238 91160 118294 91216
rect 120446 91160 120502 91216
rect 121366 91160 121422 91216
rect 122746 91160 122802 91216
rect 124034 91296 124090 91352
rect 125414 91296 125470 91352
rect 124126 91160 124182 91216
rect 125506 91160 125562 91216
rect 126794 91160 126850 91216
rect 130750 92404 130806 92440
rect 130750 92384 130752 92404
rect 130752 92384 130804 92404
rect 130804 92384 130806 92404
rect 151542 92384 151598 92440
rect 152922 92384 152978 92440
rect 151358 91976 151414 92032
rect 132222 91568 132278 91624
rect 129646 91160 129702 91216
rect 136454 91160 136510 91216
rect 167550 110064 167606 110120
rect 173162 293936 173218 293992
rect 167734 111732 167736 111752
rect 167736 111732 167788 111752
rect 167788 111732 167790 111752
rect 167734 111696 167790 111732
rect 167734 108704 167790 108760
rect 169298 92248 169354 92304
rect 173898 175888 173954 175944
rect 174634 92112 174690 92168
rect 176658 354320 176714 354376
rect 176566 352144 176622 352200
rect 176474 336504 176530 336560
rect 176014 292576 176070 292632
rect 176382 263744 176438 263800
rect 176658 348064 176714 348120
rect 176658 343304 176714 343360
rect 176658 341264 176714 341320
rect 176658 332596 176660 332616
rect 176660 332596 176712 332616
rect 176712 332596 176714 332616
rect 176658 332560 176714 332596
rect 176658 321580 176660 321600
rect 176660 321580 176712 321600
rect 176712 321580 176714 321600
rect 176658 321544 176714 321580
rect 177762 318824 177818 318880
rect 176658 314744 176714 314800
rect 176658 309984 176714 310040
rect 176658 307944 176714 308000
rect 176658 305904 176714 305960
rect 177670 301144 177726 301200
rect 176658 299240 176714 299296
rect 176658 297200 176714 297256
rect 176658 295024 176714 295080
rect 176658 292304 176714 292360
rect 176658 290264 176714 290320
rect 176658 281560 176714 281616
rect 176750 279520 176806 279576
rect 176658 277480 176714 277536
rect 176658 274760 176714 274816
rect 176658 272720 176714 272776
rect 176658 268504 176714 268560
rect 176658 265920 176714 265976
rect 176658 261840 176714 261896
rect 176658 259664 176714 259720
rect 176842 254904 176898 254960
rect 176842 254088 176898 254144
rect 176658 250824 176714 250880
rect 176842 242120 176898 242176
rect 177946 334620 178002 334656
rect 177946 334600 177948 334620
rect 177948 334600 178000 334620
rect 178000 334600 178002 334620
rect 178958 312704 179014 312760
rect 177946 303864 178002 303920
rect 177854 286340 177910 286376
rect 177854 286320 177856 286340
rect 177856 286320 177908 286340
rect 177908 286320 177910 286340
rect 177854 270544 177910 270600
rect 179050 279520 179106 279576
rect 179234 288224 179290 288280
rect 179602 355000 179658 355056
rect 189998 363024 190054 363080
rect 182914 357720 182970 357776
rect 206282 356088 206338 356144
rect 233790 361664 233846 361720
rect 218334 357584 218390 357640
rect 231214 357856 231270 357912
rect 227350 357448 227406 357504
rect 228822 356088 228878 356144
rect 209870 354864 209926 354920
rect 240046 356224 240102 356280
rect 250534 357584 250590 357640
rect 262218 354728 262274 354784
rect 291750 354592 291806 354648
rect 179510 351872 179566 351928
rect 293958 352280 294014 352336
rect 293038 330384 293094 330440
rect 179510 325712 179566 325748
rect 179510 325692 179512 325712
rect 179512 325692 179564 325712
rect 179564 325692 179566 325712
rect 179510 316852 179566 316908
rect 179418 256944 179474 257000
rect 179326 254904 179382 254960
rect 179418 252864 179474 252920
rect 179234 248104 179290 248160
rect 179142 245928 179198 245984
rect 179326 244024 179382 244080
rect 293130 301280 293186 301336
rect 293038 287408 293094 287464
rect 179510 242936 179566 242992
rect 188342 240624 188398 240680
rect 186962 175888 187018 175944
rect 189998 238992 190054 239048
rect 192482 184320 192538 184376
rect 198002 196560 198058 196616
rect 196622 193840 196678 193896
rect 196898 94832 196954 94888
rect 204902 238448 204958 238504
rect 202326 90888 202382 90944
rect 214562 184320 214618 184376
rect 213918 175616 213974 175672
rect 213918 174936 213974 174992
rect 213918 173576 213974 173632
rect 214654 174256 214710 174312
rect 214010 172896 214066 172952
rect 213918 172216 213974 172272
rect 214746 171536 214802 171592
rect 213918 171012 213974 171048
rect 213918 170992 213920 171012
rect 213920 170992 213972 171012
rect 213972 170992 213974 171012
rect 214010 170312 214066 170368
rect 213918 168292 213974 168328
rect 213918 168272 213920 168292
rect 213920 168272 213972 168292
rect 213972 168272 213974 168292
rect 214010 167592 214066 167648
rect 213918 166368 213974 166424
rect 214102 166912 214158 166968
rect 214010 165688 214066 165744
rect 213918 165008 213974 165064
rect 214010 164328 214066 164384
rect 213918 163648 213974 163704
rect 214010 162968 214066 163024
rect 213918 162288 213974 162344
rect 214010 161744 214066 161800
rect 214930 169632 214986 169688
rect 214562 161064 214618 161120
rect 214102 160656 214158 160712
rect 213918 160384 213974 160440
rect 213918 159704 213974 159760
rect 214010 159024 214066 159080
rect 213918 157664 213974 157720
rect 214654 158344 214710 158400
rect 214102 157120 214158 157176
rect 213918 156440 213974 156496
rect 213918 155796 213920 155816
rect 213920 155796 213972 155816
rect 213972 155796 213974 155816
rect 213918 155760 213974 155796
rect 214010 155080 214066 155136
rect 214010 154400 214066 154456
rect 213918 153720 213974 153776
rect 213918 153040 213974 153096
rect 214010 152496 214066 152552
rect 214378 151816 214434 151872
rect 214010 151136 214066 151192
rect 213918 150476 213974 150512
rect 213918 150456 213920 150476
rect 213920 150456 213972 150476
rect 213972 150456 213974 150476
rect 214010 149776 214066 149832
rect 213918 149096 213974 149152
rect 213918 148416 213974 148472
rect 213918 147872 213974 147928
rect 214010 147192 214066 147248
rect 213918 146512 213974 146568
rect 214010 145832 214066 145888
rect 213918 145152 213974 145208
rect 214010 144472 214066 144528
rect 213918 143792 213974 143848
rect 213918 143248 213974 143304
rect 214746 142568 214802 142624
rect 213918 141888 213974 141944
rect 214010 141208 214066 141264
rect 213918 140528 213974 140584
rect 213182 139848 213238 139904
rect 214010 139168 214066 139224
rect 213918 138624 213974 138680
rect 214654 137944 214710 138000
rect 213918 137264 213974 137320
rect 214562 136584 214618 136640
rect 214010 135904 214066 135960
rect 213918 135260 213920 135280
rect 213920 135260 213972 135280
rect 213972 135260 213974 135280
rect 213918 135224 213974 135260
rect 213918 133900 213920 133920
rect 213920 133900 213972 133920
rect 213972 133900 213974 133920
rect 213918 133864 213974 133900
rect 213918 133320 213974 133376
rect 213918 131280 213974 131336
rect 213918 129920 213974 129976
rect 213918 129240 213974 129296
rect 214010 128016 214066 128072
rect 213918 127336 213974 127392
rect 213918 126656 213974 126712
rect 214470 125976 214526 126032
rect 214010 125296 214066 125352
rect 213918 124616 213974 124672
rect 214010 124072 214066 124128
rect 213918 123392 213974 123448
rect 214010 122712 214066 122768
rect 213918 122032 213974 122088
rect 214010 121352 214066 121408
rect 213918 120672 213974 120728
rect 214102 119992 214158 120048
rect 214010 119448 214066 119504
rect 213918 118804 213920 118824
rect 213920 118804 213972 118824
rect 213972 118804 213974 118824
rect 213918 118768 213974 118804
rect 214010 118088 214066 118144
rect 213918 117408 213974 117464
rect 214010 116728 214066 116784
rect 213918 116048 213974 116104
rect 214010 115368 214066 115424
rect 213918 114824 213974 114880
rect 214010 114144 214066 114200
rect 213918 113464 213974 113520
rect 213918 112784 213974 112840
rect 214010 111424 214066 111480
rect 213918 110744 213974 110800
rect 213918 110200 213974 110256
rect 214010 108840 214066 108896
rect 213918 108160 213974 108216
rect 213918 107480 213974 107536
rect 214470 106800 214526 106856
rect 214010 106120 214066 106176
rect 213918 105576 213974 105632
rect 214010 104216 214066 104272
rect 213918 103572 213920 103592
rect 213920 103572 213972 103592
rect 213972 103572 213974 103592
rect 213918 103536 213974 103572
rect 214010 102856 214066 102912
rect 213918 102196 213974 102232
rect 213918 102176 213920 102196
rect 213920 102176 213972 102196
rect 213972 102176 213974 102196
rect 213918 100952 213974 101008
rect 214102 100272 214158 100328
rect 213918 99592 213974 99648
rect 214010 98912 214066 98968
rect 213918 98232 213974 98288
rect 213918 97552 213974 97608
rect 214930 130600 214986 130656
rect 214746 112104 214802 112160
rect 214654 96872 214710 96928
rect 214562 96328 214618 96384
rect 214838 101496 214894 101552
rect 232502 185544 232558 185600
rect 239494 180104 239550 180160
rect 242254 210568 242310 210624
rect 239402 177248 239458 177304
rect 244922 176024 244978 176080
rect 250810 238040 250866 238096
rect 247774 177656 247830 177712
rect 248050 175788 248052 175808
rect 248052 175788 248104 175808
rect 248104 175788 248106 175808
rect 248050 175752 248106 175788
rect 249154 174664 249210 174720
rect 249338 173304 249394 173360
rect 249246 172352 249302 172408
rect 250074 175208 250130 175264
rect 250074 159160 250130 159216
rect 251362 170040 251418 170096
rect 252098 172760 252154 172816
rect 252466 171808 252522 171864
rect 252558 171400 252614 171456
rect 251730 170892 251732 170912
rect 251732 170892 251784 170912
rect 251784 170892 251786 170912
rect 251362 160112 251418 160168
rect 251270 159568 251326 159624
rect 251178 158752 251234 158808
rect 251730 170856 251786 170892
rect 251822 170448 251878 170504
rect 252466 169496 252522 169552
rect 252282 169088 252338 169144
rect 252466 168136 252522 168192
rect 252466 167592 252522 167648
rect 251914 167184 251970 167240
rect 252098 166640 252154 166696
rect 252374 166368 252430 166424
rect 252466 165688 252522 165744
rect 251730 164736 251786 164792
rect 252466 165280 252522 165336
rect 252098 164328 252154 164384
rect 252190 162968 252246 163024
rect 252466 162424 252522 162480
rect 253202 163920 253258 163976
rect 253202 162968 253258 163024
rect 252466 160520 252522 160576
rect 251914 157800 251970 157856
rect 252466 157292 252468 157312
rect 252468 157292 252520 157312
rect 252520 157292 252522 157312
rect 252466 157256 252522 157292
rect 251546 156848 251602 156904
rect 252374 156304 252430 156360
rect 251914 155916 251970 155952
rect 251914 155896 251916 155916
rect 251916 155896 251968 155916
rect 251968 155896 251970 155916
rect 251178 155352 251234 155408
rect 252466 154944 252522 155000
rect 251086 154400 251142 154456
rect 251638 153992 251694 154048
rect 252466 153448 252522 153504
rect 250534 152904 250590 152960
rect 249982 141344 250038 141400
rect 249798 138488 249854 138544
rect 241518 94424 241574 94480
rect 242898 3304 242954 3360
rect 249154 97008 249210 97064
rect 252466 153060 252522 153096
rect 252466 153040 252468 153060
rect 252468 153040 252520 153060
rect 252520 153040 252522 153060
rect 252374 152632 252430 152688
rect 251914 152088 251970 152144
rect 252466 151680 252522 151736
rect 252374 151136 252430 151192
rect 251914 150728 251970 150784
rect 251178 149776 251234 149832
rect 252466 150220 252468 150240
rect 252468 150220 252520 150240
rect 252520 150220 252522 150240
rect 252466 150184 252522 150220
rect 252006 149232 252062 149288
rect 251914 148860 251916 148880
rect 251916 148860 251968 148880
rect 251968 148860 251970 148880
rect 251914 148824 251970 148860
rect 251822 143112 251878 143168
rect 250534 136584 250590 136640
rect 252466 148280 252522 148336
rect 252466 147464 252522 147520
rect 252374 146512 252430 146568
rect 252466 145968 252522 146024
rect 252282 145560 252338 145616
rect 252098 145016 252154 145072
rect 252098 143656 252154 143712
rect 252466 144064 252522 144120
rect 252282 142704 252338 142760
rect 251638 134680 251694 134736
rect 251454 133320 251510 133376
rect 251546 131824 251602 131880
rect 251546 130872 251602 130928
rect 252098 140392 252154 140448
rect 252098 137536 252154 137592
rect 252098 136176 252154 136232
rect 251822 130056 251878 130112
rect 252006 132776 252062 132832
rect 251730 129104 251786 129160
rect 252466 137944 252522 138000
rect 252374 136992 252430 137048
rect 252374 135632 252430 135688
rect 252466 135224 252522 135280
rect 252466 134272 252522 134328
rect 252466 133764 252468 133784
rect 252468 133764 252520 133784
rect 252520 133764 252522 133784
rect 252466 133728 252522 133764
rect 252466 132404 252468 132424
rect 252468 132404 252520 132424
rect 252520 132404 252522 132424
rect 252466 132368 252522 132404
rect 252282 131416 252338 131472
rect 252466 130464 252522 130520
rect 251178 125332 251180 125352
rect 251180 125332 251232 125352
rect 251232 125332 251234 125352
rect 251178 125296 251234 125332
rect 251270 124752 251326 124808
rect 251730 122984 251786 123040
rect 252466 129548 252468 129568
rect 252468 129548 252520 129568
rect 252520 129548 252522 129568
rect 252466 129512 252522 129548
rect 252006 128560 252062 128616
rect 252466 128188 252468 128208
rect 252468 128188 252520 128208
rect 252520 128188 252522 128208
rect 252466 128152 252522 128188
rect 252374 127608 252430 127664
rect 252006 127200 252062 127256
rect 251914 126248 251970 126304
rect 252466 126692 252468 126712
rect 252468 126692 252520 126712
rect 252520 126692 252522 126712
rect 252466 126656 252522 126692
rect 252190 125704 252246 125760
rect 252190 124344 252246 124400
rect 252466 123936 252522 123992
rect 251914 120536 251970 120592
rect 251822 118768 251878 118824
rect 251546 118224 251602 118280
rect 251546 116900 251548 116920
rect 251548 116900 251600 116920
rect 251600 116900 251602 116920
rect 251546 116864 251602 116900
rect 251638 115368 251694 115424
rect 251730 110744 251786 110800
rect 251546 110200 251602 110256
rect 251454 109248 251510 109304
rect 252098 123392 252154 123448
rect 252098 120128 252154 120184
rect 252098 117272 252154 117328
rect 252466 122440 252522 122496
rect 252374 122032 252430 122088
rect 252466 121524 252468 121544
rect 252468 121524 252520 121544
rect 252520 121524 252522 121544
rect 252466 121488 252522 121524
rect 252466 121080 252522 121136
rect 252466 119584 252522 119640
rect 252374 119176 252430 119232
rect 252466 117816 252522 117872
rect 252374 116320 252430 116376
rect 252282 115912 252338 115968
rect 252374 114960 252430 115016
rect 252466 114452 252468 114472
rect 252468 114452 252520 114472
rect 252520 114452 252522 114472
rect 252466 114416 252522 114452
rect 252466 114008 252522 114064
rect 252006 113464 252062 113520
rect 251914 112648 251970 112704
rect 251178 108876 251180 108896
rect 251180 108876 251232 108896
rect 251232 108876 251234 108896
rect 251178 108840 251234 108876
rect 251546 106528 251602 106584
rect 251178 105984 251234 106040
rect 251822 108296 251878 108352
rect 251914 107888 251970 107944
rect 251730 104624 251786 104680
rect 252190 113076 252246 113112
rect 252190 113056 252192 113076
rect 252192 113056 252244 113076
rect 252244 113056 252246 113076
rect 252098 112104 252154 112160
rect 252374 111732 252376 111752
rect 252376 111732 252428 111752
rect 252428 111732 252430 111752
rect 252374 111696 252430 111732
rect 252006 103672 252062 103728
rect 252466 109792 252522 109848
rect 252466 107516 252468 107536
rect 252468 107516 252520 107536
rect 252520 107516 252522 107536
rect 252466 107480 252522 107516
rect 252374 106936 252430 106992
rect 252374 105576 252430 105632
rect 252282 105032 252338 105088
rect 252466 104080 252522 104136
rect 252282 102720 252338 102776
rect 252466 103128 252522 103184
rect 252374 102176 252430 102232
rect 252190 101360 252246 101416
rect 252466 100816 252522 100872
rect 252006 100408 252062 100464
rect 252466 99864 252522 99920
rect 252098 99456 252154 99512
rect 252466 98912 252522 98968
rect 252374 98504 252430 98560
rect 251638 97960 251694 98016
rect 252466 97552 252522 97608
rect 251178 96600 251234 96656
rect 251270 96192 251326 96248
rect 256698 138624 256754 138680
rect 255870 3440 255926 3496
rect 257526 148280 257582 148336
rect 258998 144064 259054 144120
rect 264978 233144 265034 233200
rect 262218 162016 262274 162072
rect 264150 3304 264206 3360
rect 269762 238448 269818 238504
rect 273718 238856 273774 238912
rect 269762 231648 269818 231704
rect 276662 227568 276718 227624
rect 287058 231784 287114 231840
rect 287702 166232 287758 166288
rect 285770 80688 285826 80744
rect 293222 259120 293278 259176
rect 293314 241848 293370 241904
rect 293314 241032 293370 241088
rect 294142 338680 294198 338736
rect 294050 327800 294106 327856
rect 294050 325760 294106 325816
rect 294142 323040 294198 323096
rect 295338 343440 295394 343496
rect 295338 340720 295394 340776
rect 295430 334600 295486 334656
rect 295338 331880 295394 331936
rect 294418 327800 294474 327856
rect 294234 303320 294290 303376
rect 295614 354320 295670 354376
rect 296166 345480 296222 345536
rect 295614 336640 295670 336696
rect 295522 321000 295578 321056
rect 295522 318960 295578 319016
rect 295614 316920 295670 316976
rect 295522 314200 295578 314256
rect 295522 312160 295578 312216
rect 295522 310120 295578 310176
rect 295522 308080 295578 308136
rect 295430 305360 295486 305416
rect 295430 296520 295486 296576
rect 295338 294480 295394 294536
rect 294234 267960 294290 268016
rect 296626 299240 296682 299296
rect 295614 292440 295670 292496
rect 295338 243480 295394 243536
rect 295338 241440 295394 241496
rect 295522 290400 295578 290456
rect 295522 285676 295524 285696
rect 295524 285676 295576 285696
rect 295576 285676 295578 285696
rect 295522 285640 295578 285676
rect 295522 283600 295578 283656
rect 295522 281580 295578 281616
rect 295522 281560 295524 281580
rect 295524 281560 295576 281580
rect 295576 281560 295578 281580
rect 295522 278840 295578 278896
rect 295614 276800 295670 276856
rect 295706 274760 295762 274816
rect 295614 272720 295670 272776
rect 295614 270000 295670 270056
rect 295614 265920 295670 265976
rect 295614 263880 295670 263936
rect 295614 261160 295670 261216
rect 295706 257100 295762 257136
rect 295706 257080 295708 257100
rect 295708 257080 295760 257100
rect 295760 257080 295762 257100
rect 295706 255040 295762 255096
rect 296442 252320 296498 252376
rect 295798 250280 295854 250336
rect 296626 248240 296682 248296
rect 296902 246200 296958 246256
rect 298742 357448 298798 357504
rect 298098 354592 298154 354648
rect 297362 238856 297418 238912
rect 298098 228248 298154 228304
rect 299478 355000 299534 355056
rect 293682 3440 293738 3496
rect 296074 3440 296130 3496
rect 299662 247016 299718 247072
rect 299754 241848 299810 241904
rect 300950 241168 301006 241224
rect 300766 149640 300822 149696
rect 302330 238584 302386 238640
rect 305182 237224 305238 237280
rect 307574 175616 307630 175672
rect 307114 175208 307170 175264
rect 306746 174800 306802 174856
rect 306562 173576 306618 173632
rect 306930 173168 306986 173224
rect 306930 172216 306986 172272
rect 306746 170584 306802 170640
rect 306930 169768 306986 169824
rect 307022 165008 307078 165064
rect 306746 163784 306802 163840
rect 306470 161608 306526 161664
rect 306562 160384 306618 160440
rect 306930 159976 306986 160032
rect 306930 158616 306986 158672
rect 306654 152632 306710 152688
rect 306746 150592 306802 150648
rect 306746 149776 306802 149832
rect 306654 143792 306710 143848
rect 305734 143656 305790 143712
rect 305642 131688 305698 131744
rect 305642 104896 305698 104952
rect 306562 143384 306618 143440
rect 306010 142296 306066 142352
rect 306562 142296 306618 142352
rect 305826 107752 305882 107808
rect 305734 100816 305790 100872
rect 306930 142024 306986 142080
rect 306562 141344 306618 141400
rect 307666 174392 307722 174448
rect 307574 173984 307630 174040
rect 307298 172644 307354 172680
rect 307298 172624 307300 172644
rect 307300 172624 307352 172644
rect 307352 172624 307354 172644
rect 307574 171808 307630 171864
rect 307666 171400 307722 171456
rect 307206 170992 307262 171048
rect 307666 170176 307722 170232
rect 307482 169224 307538 169280
rect 307574 168816 307630 168872
rect 307666 168408 307722 168464
rect 307482 168000 307538 168056
rect 307298 167204 307354 167240
rect 307298 167184 307300 167204
rect 307300 167184 307352 167204
rect 307352 167184 307354 167204
rect 307666 167592 307722 167648
rect 307574 166776 307630 166832
rect 307482 166368 307538 166424
rect 307390 165416 307446 165472
rect 307298 164228 307300 164248
rect 307300 164228 307352 164248
rect 307352 164228 307354 164248
rect 307298 164192 307354 164228
rect 307298 163004 307300 163024
rect 307300 163004 307352 163024
rect 307352 163004 307354 163024
rect 307298 162968 307354 163004
rect 307114 159568 307170 159624
rect 307666 165824 307722 165880
rect 307666 164600 307722 164656
rect 307666 163376 307722 163432
rect 307482 162424 307538 162480
rect 307666 162016 307722 162072
rect 307574 161200 307630 161256
rect 307666 160792 307722 160848
rect 307666 159024 307722 159080
rect 307482 158208 307538 158264
rect 307666 157800 307722 157856
rect 307482 156984 307538 157040
rect 307574 156576 307630 156632
rect 307666 156168 307722 156224
rect 307666 155624 307722 155680
rect 307482 155216 307538 155272
rect 307574 154400 307630 154456
rect 307482 153992 307538 154048
rect 307666 153584 307722 153640
rect 307206 153176 307262 153232
rect 307114 145016 307170 145072
rect 306102 140800 306158 140856
rect 306562 137400 306618 137456
rect 307022 131824 307078 131880
rect 306746 131008 306802 131064
rect 306746 127200 306802 127256
rect 306746 126792 306802 126848
rect 306746 125024 306802 125080
rect 306562 123800 306618 123856
rect 307114 127608 307170 127664
rect 307114 124244 307116 124264
rect 307116 124244 307168 124264
rect 307168 124244 307170 124264
rect 307114 124208 307170 124244
rect 306746 122440 306802 122496
rect 306746 121216 306802 121272
rect 306746 119584 306802 119640
rect 307022 116184 307078 116240
rect 306562 112648 306618 112704
rect 306746 111424 306802 111480
rect 306562 111016 306618 111072
rect 306746 110200 306802 110256
rect 306746 105848 306802 105904
rect 305918 105032 305974 105088
rect 306746 105032 306802 105088
rect 306562 102992 306618 103048
rect 306562 101632 306618 101688
rect 306746 100408 306802 100464
rect 306562 100000 306618 100056
rect 306746 99048 306802 99104
rect 306930 96192 306986 96248
rect 307574 152224 307630 152280
rect 307666 151836 307722 151872
rect 307666 151816 307668 151836
rect 307668 151816 307720 151836
rect 307720 151816 307722 151836
rect 307482 151408 307538 151464
rect 307666 151000 307722 151056
rect 307574 150184 307630 150240
rect 307666 149232 307722 149288
rect 307574 148824 307630 148880
rect 307390 148416 307446 148472
rect 307298 147600 307354 147656
rect 307666 148008 307722 148064
rect 307482 147192 307538 147248
rect 307574 146784 307630 146840
rect 307666 146412 307668 146432
rect 307668 146412 307720 146432
rect 307720 146412 307722 146432
rect 307666 146376 307722 146412
rect 307482 145832 307538 145888
rect 307666 145424 307722 145480
rect 307574 144608 307630 144664
rect 307666 144200 307722 144256
rect 307574 143656 307630 143712
rect 307574 142976 307630 143032
rect 307666 142432 307722 142488
rect 307298 141616 307354 141672
rect 307390 141208 307446 141264
rect 307482 140392 307538 140448
rect 307574 139984 307630 140040
rect 307666 139596 307722 139632
rect 307666 139576 307668 139596
rect 307668 139576 307720 139596
rect 307720 139576 307722 139596
rect 307482 139032 307538 139088
rect 307574 138624 307630 138680
rect 307666 138216 307722 138272
rect 307574 137808 307630 137864
rect 307666 136992 307722 137048
rect 307482 136584 307538 136640
rect 307574 136176 307630 136232
rect 307666 135632 307722 135688
rect 307666 135260 307668 135280
rect 307668 135260 307720 135280
rect 307720 135260 307722 135280
rect 307666 135224 307722 135260
rect 307482 134816 307538 134872
rect 307666 134408 307722 134464
rect 307574 134000 307630 134056
rect 307390 133592 307446 133648
rect 307390 129240 307446 129296
rect 307574 133184 307630 133240
rect 307666 132640 307722 132696
rect 307666 132232 307722 132288
rect 307574 130192 307630 130248
rect 307666 129784 307722 129840
rect 307666 128832 307722 128888
rect 307574 128424 307630 128480
rect 307666 128016 307722 128072
rect 307666 125840 307722 125896
rect 307574 125432 307630 125488
rect 307666 124616 307722 124672
rect 307574 123392 307630 123448
rect 307666 122984 307722 123040
rect 307574 122032 307630 122088
rect 307666 121624 307722 121680
rect 307574 120808 307630 120864
rect 307666 120400 307722 120456
rect 307666 119992 307722 120048
rect 307482 118224 307538 118280
rect 307666 117816 307722 117872
rect 307666 117000 307722 117056
rect 307482 116592 307538 116648
rect 307482 115640 307538 115696
rect 307574 115232 307630 115288
rect 307666 114824 307722 114880
rect 307666 113600 307722 113656
rect 307574 113228 307576 113248
rect 307576 113228 307628 113248
rect 307628 113228 307630 113248
rect 307574 113192 307630 113228
rect 307666 112240 307722 112296
rect 307298 111832 307354 111888
rect 307298 110608 307354 110664
rect 307574 109792 307630 109848
rect 307666 109248 307722 109304
rect 307574 108840 307630 108896
rect 307482 108432 307538 108488
rect 307666 108024 307722 108080
rect 307574 107752 307630 107808
rect 307298 107616 307354 107672
rect 307482 107208 307538 107264
rect 307298 106800 307354 106856
rect 307666 106428 307668 106448
rect 307668 106428 307720 106448
rect 307720 106428 307722 106448
rect 307666 106392 307722 106428
rect 307666 105440 307722 105496
rect 307482 104624 307538 104680
rect 307666 104216 307722 104272
rect 307574 103808 307630 103864
rect 307574 103400 307630 103456
rect 307666 102448 307722 102504
rect 307482 102040 307538 102096
rect 307666 101224 307722 101280
rect 307482 100816 307538 100872
rect 307666 100836 307722 100872
rect 307666 100816 307668 100836
rect 307668 100816 307720 100836
rect 307720 100816 307722 100836
rect 307666 99592 307722 99648
rect 307206 98640 307262 98696
rect 307666 98232 307722 98288
rect 307574 97824 307630 97880
rect 307298 97416 307354 97472
rect 307666 97008 307722 97064
rect 307666 96636 307668 96656
rect 307668 96636 307720 96656
rect 307720 96636 307722 96656
rect 307666 96600 307722 96636
rect 303618 25608 303674 25664
rect 303158 6160 303214 6216
rect 305550 6296 305606 6352
rect 309138 114416 309194 114472
rect 309138 113056 309194 113112
rect 313278 229744 313334 229800
rect 311162 177384 311218 177440
rect 313922 178744 313978 178800
rect 317418 189624 317474 189680
rect 315302 177248 315358 177304
rect 316038 176704 316094 176760
rect 319442 176160 319498 176216
rect 320178 176704 320234 176760
rect 320822 176704 320878 176760
rect 321650 176704 321706 176760
rect 321466 175752 321522 175808
rect 321282 172624 321338 172680
rect 321466 171400 321522 171456
rect 321466 169632 321522 169688
rect 321834 175208 321890 175264
rect 321926 171128 321982 171184
rect 321742 167456 321798 167512
rect 321650 150320 321706 150376
rect 321558 132640 321614 132696
rect 323030 184184 323086 184240
rect 323122 165416 323178 165472
rect 323030 150864 323086 150920
rect 324410 173984 324466 174040
rect 324318 173168 324374 173224
rect 324318 168544 324374 168600
rect 324318 167728 324374 167784
rect 324318 164736 324374 164792
rect 324318 163920 324374 163976
rect 324410 163104 324466 163160
rect 324318 162424 324374 162480
rect 324410 161608 324466 161664
rect 324318 160792 324374 160848
rect 324410 160112 324466 160168
rect 324318 159296 324374 159352
rect 324318 158480 324374 158536
rect 324410 157800 324466 157856
rect 324318 156984 324374 157040
rect 324318 155488 324374 155544
rect 324410 154672 324466 154728
rect 324318 153992 324374 154048
rect 324318 153176 324374 153232
rect 324686 166232 324742 166288
rect 324502 152360 324558 152416
rect 324318 151716 324320 151736
rect 324320 151716 324372 151736
rect 324372 151716 324374 151736
rect 324318 151680 324374 151716
rect 324318 149368 324374 149424
rect 324318 148552 324374 148608
rect 324410 147736 324466 147792
rect 324318 147056 324374 147112
rect 324318 143928 324374 143984
rect 324318 143112 324374 143168
rect 324318 141616 324374 141672
rect 324318 140120 324374 140176
rect 324318 139340 324320 139360
rect 324320 139340 324372 139360
rect 324372 139340 324374 139360
rect 324318 139304 324374 139340
rect 324318 137844 324320 137864
rect 324320 137844 324372 137864
rect 324372 137844 324374 137864
rect 324318 137808 324374 137844
rect 324410 136992 324466 137048
rect 324318 136348 324320 136368
rect 324320 136348 324372 136368
rect 324372 136348 324374 136368
rect 324318 136312 324374 136348
rect 324410 135496 324466 135552
rect 324594 142432 324650 142488
rect 324594 140800 324650 140856
rect 324502 133184 324558 133240
rect 324318 131688 324374 131744
rect 324318 130872 324374 130928
rect 324410 130056 324466 130112
rect 324318 129376 324374 129432
rect 324410 128560 324466 128616
rect 324318 127744 324374 127800
rect 324410 127064 324466 127120
rect 324318 124752 324374 124808
rect 324318 123120 324374 123176
rect 324318 122440 324374 122496
rect 324318 120808 324374 120864
rect 324410 120128 324466 120184
rect 324318 119312 324374 119368
rect 324318 118496 324374 118552
rect 324410 117816 324466 117872
rect 324318 117000 324374 117056
rect 324410 116320 324466 116376
rect 324318 115504 324374 115560
rect 324318 114008 324374 114064
rect 324410 113192 324466 113248
rect 324318 112376 324374 112432
rect 324318 111732 324320 111752
rect 324320 111732 324372 111752
rect 324372 111732 324374 111752
rect 324318 111696 324374 111732
rect 324318 109384 324374 109440
rect 324318 108568 324374 108624
rect 325606 107752 325662 107808
rect 325882 156304 325938 156360
rect 325790 125432 325846 125488
rect 323030 107072 323086 107128
rect 322938 103128 322994 103184
rect 321558 101088 321614 101144
rect 321466 97280 321522 97336
rect 309046 3984 309102 4040
rect 307942 3304 307998 3360
rect 313278 18672 313334 18728
rect 321650 98776 321706 98832
rect 324318 105440 324374 105496
rect 324318 104796 324320 104816
rect 324320 104796 324372 104816
rect 324372 104796 324374 104816
rect 324318 104760 324374 104796
rect 327722 204856 327778 204912
rect 324318 103944 324374 104000
rect 324502 100816 324558 100872
rect 324410 100136 324466 100192
rect 324410 92384 324466 92440
rect 324594 97008 324650 97064
rect 324502 91024 324558 91080
rect 321558 73752 321614 73808
rect 331218 12960 331274 13016
rect 332690 181328 332746 181384
rect 336922 178608 336978 178664
rect 338394 175888 338450 175944
rect 336738 53080 336794 53136
rect 339498 22616 339554 22672
rect 342166 3440 342222 3496
rect 543462 702480 543518 702536
rect 580354 702616 580410 702672
rect 356702 61376 356758 61432
rect 580354 697176 580410 697232
rect 580170 683848 580226 683904
rect 580262 670656 580318 670712
rect 579986 630808 580042 630864
rect 580170 617480 580226 617536
rect 580170 590960 580226 591016
rect 579894 564304 579950 564360
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 471416 580226 471472
rect 580170 458088 580226 458144
rect 579986 404912 580042 404968
rect 580170 378392 580226 378448
rect 582378 644000 582434 644056
rect 580354 577632 580410 577688
rect 580170 365064 580226 365120
rect 580262 351872 580318 351928
rect 580170 325216 580226 325272
rect 579618 298696 579674 298752
rect 579618 258848 579674 258904
rect 579894 245520 579950 245576
rect 579618 232328 579674 232384
rect 580170 219000 580226 219056
rect 580170 179152 580226 179208
rect 580354 312024 580410 312080
rect 580354 272176 580410 272232
rect 582470 537784 582526 537840
rect 582562 431568 582618 431624
rect 582654 418240 582710 418296
rect 580262 165824 580318 165880
rect 582378 205672 582434 205728
rect 580446 192480 580502 192536
rect 580354 152632 580410 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 579802 112784 579858 112840
rect 580170 99456 580226 99512
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 47504 580226 47560
rect 580170 46280 580226 46336
rect 579986 19760 580042 19816
rect 582470 33088 582526 33144
rect 582378 6568 582434 6624
<< obsm2 >>
rect 68800 95100 164756 174600
<< metal3 >>
rect 179270 702612 179276 702676
rect 179340 702674 179346 702676
rect 580349 702674 580415 702677
rect 179340 702672 580415 702674
rect 179340 702616 580354 702672
rect 580410 702616 580415 702672
rect 179340 702614 580415 702616
rect 179340 702612 179346 702614
rect 580349 702611 580415 702614
rect 180558 702476 180564 702540
rect 180628 702538 180634 702540
rect 543457 702538 543523 702541
rect 180628 702536 543523 702538
rect 180628 702480 543462 702536
rect 543518 702480 543523 702536
rect 180628 702478 543523 702480
rect 180628 702476 180634 702478
rect 543457 702475 543523 702478
rect -960 697220 480 697460
rect 580349 697234 580415 697237
rect 583520 697234 584960 697324
rect 580349 697232 584960 697234
rect 580349 697176 580354 697232
rect 580410 697176 584960 697232
rect 580349 697174 584960 697176
rect 580349 697171 580415 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580257 670714 580323 670717
rect 583520 670714 584960 670804
rect 580257 670712 584960 670714
rect 580257 670656 580262 670712
rect 580318 670656 584960 670712
rect 580257 670654 584960 670656
rect 580257 670651 580323 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 2773 658202 2839 658205
rect -960 658200 2839 658202
rect -960 658144 2778 658200
rect 2834 658144 2839 658200
rect -960 658142 2839 658144
rect -960 658052 480 658142
rect 2773 658139 2839 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 582373 644058 582439 644061
rect 583520 644058 584960 644148
rect 582373 644056 584960 644058
rect 582373 644000 582378 644056
rect 582434 644000 584960 644056
rect 582373 643998 584960 644000
rect 582373 643995 582439 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 579981 630866 580047 630869
rect 583520 630866 584960 630956
rect 579981 630864 584960 630866
rect 579981 630808 579986 630864
rect 580042 630808 584960 630864
rect 579981 630806 584960 630808
rect 579981 630803 580047 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3417 606114 3483 606117
rect -960 606112 3483 606114
rect -960 606056 3422 606112
rect 3478 606056 3483 606112
rect -960 606054 3483 606056
rect -960 605964 480 606054
rect 3417 606051 3483 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580349 577690 580415 577693
rect 583520 577690 584960 577780
rect 580349 577688 584960 577690
rect 580349 577632 580354 577688
rect 580410 577632 584960 577688
rect 580349 577630 584960 577632
rect 580349 577627 580415 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 579889 564362 579955 564365
rect 583520 564362 584960 564452
rect 579889 564360 584960 564362
rect 579889 564304 579894 564360
rect 579950 564304 584960 564360
rect 579889 564302 584960 564304
rect 579889 564299 579955 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 582465 537842 582531 537845
rect 583520 537842 584960 537932
rect 582465 537840 584960 537842
rect 582465 537784 582470 537840
rect 582526 537784 584960 537840
rect 582465 537782 584960 537784
rect 582465 537779 582531 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 120022 514858 120028 514860
rect -960 514798 120028 514858
rect -960 514708 480 514798
rect 120022 514796 120028 514798
rect 120092 514796 120098 514860
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3417 501802 3483 501805
rect -960 501800 3483 501802
rect -960 501744 3422 501800
rect 3478 501744 3483 501800
rect -960 501742 3483 501744
rect -960 501652 480 501742
rect 3417 501739 3483 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484666 584960 484756
rect 567150 484606 584960 484666
rect 299974 484468 299980 484532
rect 300044 484530 300050 484532
rect 567150 484530 567210 484606
rect 300044 484470 567210 484530
rect 583520 484516 584960 484606
rect 300044 484468 300050 484470
rect -960 475690 480 475780
rect 3049 475690 3115 475693
rect -960 475688 3115 475690
rect -960 475632 3054 475688
rect 3110 475632 3115 475688
rect -960 475630 3115 475632
rect -960 475540 480 475630
rect 3049 475627 3115 475630
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 582557 431626 582623 431629
rect 583520 431626 584960 431716
rect 582557 431624 584960 431626
rect 582557 431568 582562 431624
rect 582618 431568 584960 431624
rect 582557 431566 584960 431568
rect 582557 431563 582623 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3509 423602 3575 423605
rect -960 423600 3575 423602
rect -960 423544 3514 423600
rect 3570 423544 3575 423600
rect -960 423542 3575 423544
rect -960 423452 480 423542
rect 3509 423539 3575 423542
rect 582649 418298 582715 418301
rect 583520 418298 584960 418388
rect 582649 418296 584960 418298
rect 582649 418240 582654 418296
rect 582710 418240 584960 418296
rect 582649 418238 584960 418240
rect 582649 418235 582715 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 2865 410546 2931 410549
rect -960 410544 2931 410546
rect -960 410488 2870 410544
rect 2926 410488 2931 410544
rect -960 410486 2931 410488
rect -960 410396 480 410486
rect 2865 410483 2931 410486
rect 579981 404970 580047 404973
rect 583520 404970 584960 405060
rect 579981 404968 584960 404970
rect 579981 404912 579986 404968
rect 580042 404912 584960 404968
rect 579981 404910 584960 404912
rect 579981 404907 580047 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3509 397490 3575 397493
rect -960 397488 3575 397490
rect -960 397432 3514 397488
rect 3570 397432 3575 397488
rect -960 397430 3575 397432
rect -960 397340 480 397430
rect 3509 397427 3575 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3509 371378 3575 371381
rect -960 371376 3575 371378
rect -960 371320 3514 371376
rect 3570 371320 3575 371376
rect -960 371318 3575 371320
rect -960 371228 480 371318
rect 3509 371315 3575 371318
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect 189993 363082 190059 363085
rect 342294 363082 342300 363084
rect 189993 363080 342300 363082
rect 189993 363024 189998 363080
rect 190054 363024 342300 363080
rect 189993 363022 342300 363024
rect 189993 363019 190059 363022
rect 342294 363020 342300 363022
rect 342364 363020 342370 363084
rect 233785 361722 233851 361725
rect 332542 361722 332548 361724
rect 233785 361720 332548 361722
rect 233785 361664 233790 361720
rect 233846 361664 332548 361720
rect 233785 361662 332548 361664
rect 233785 361659 233851 361662
rect 332542 361660 332548 361662
rect 332612 361660 332618 361724
rect 114553 358866 114619 358869
rect 293902 358866 293908 358868
rect 114553 358864 293908 358866
rect 114553 358808 114558 358864
rect 114614 358808 293908 358864
rect 114553 358806 293908 358808
rect 114553 358803 114619 358806
rect 293902 358804 293908 358806
rect 293972 358804 293978 358868
rect -960 358458 480 358548
rect 3049 358458 3115 358461
rect -960 358456 3115 358458
rect -960 358400 3054 358456
rect 3110 358400 3115 358456
rect -960 358398 3115 358400
rect -960 358308 480 358398
rect 3049 358395 3115 358398
rect 150341 357914 150407 357917
rect 231209 357914 231275 357917
rect 150341 357912 231275 357914
rect 150341 357856 150346 357912
rect 150402 357856 231214 357912
rect 231270 357856 231275 357912
rect 150341 357854 231275 357856
rect 150341 357851 150407 357854
rect 231209 357851 231275 357854
rect 152958 357716 152964 357780
rect 153028 357778 153034 357780
rect 182909 357778 182975 357781
rect 153028 357776 182975 357778
rect 153028 357720 182914 357776
rect 182970 357720 182975 357776
rect 153028 357718 182975 357720
rect 153028 357716 153034 357718
rect 182909 357715 182975 357718
rect 170990 357580 170996 357644
rect 171060 357642 171066 357644
rect 218329 357642 218395 357645
rect 171060 357640 218395 357642
rect 171060 357584 218334 357640
rect 218390 357584 218395 357640
rect 171060 357582 218395 357584
rect 171060 357580 171066 357582
rect 218329 357579 218395 357582
rect 250529 357642 250595 357645
rect 297214 357642 297220 357644
rect 250529 357640 297220 357642
rect 250529 357584 250534 357640
rect 250590 357584 297220 357640
rect 250529 357582 297220 357584
rect 250529 357579 250595 357582
rect 297214 357580 297220 357582
rect 297284 357580 297290 357644
rect 227345 357506 227411 357509
rect 298737 357506 298803 357509
rect 227345 357504 298803 357506
rect 227345 357448 227350 357504
rect 227406 357448 298742 357504
rect 298798 357448 298803 357504
rect 227345 357446 298803 357448
rect 227345 357443 227411 357446
rect 298737 357443 298803 357446
rect 240041 356282 240107 356285
rect 292798 356282 292804 356284
rect 240041 356280 292804 356282
rect 240041 356224 240046 356280
rect 240102 356224 292804 356280
rect 240041 356222 292804 356224
rect 240041 356219 240107 356222
rect 292798 356220 292804 356222
rect 292868 356220 292874 356284
rect 160737 356146 160803 356149
rect 206277 356146 206343 356149
rect 160737 356144 206343 356146
rect 160737 356088 160742 356144
rect 160798 356088 206282 356144
rect 206338 356088 206343 356144
rect 160737 356086 206343 356088
rect 160737 356083 160803 356086
rect 206277 356083 206343 356086
rect 228817 356146 228883 356149
rect 301446 356146 301452 356148
rect 228817 356144 301452 356146
rect 228817 356088 228822 356144
rect 228878 356088 301452 356144
rect 228817 356086 301452 356088
rect 228817 356083 228883 356086
rect 301446 356084 301452 356086
rect 301516 356084 301522 356148
rect 179597 355058 179663 355061
rect 299473 355058 299539 355061
rect 179597 355056 299539 355058
rect 179597 355000 179602 355056
rect 179658 355000 299478 355056
rect 299534 355000 299539 355056
rect 179597 354998 299539 355000
rect 179597 354995 179663 354998
rect 299473 354995 299539 354998
rect 162117 354922 162183 354925
rect 209865 354922 209931 354925
rect 162117 354920 209931 354922
rect 162117 354864 162122 354920
rect 162178 354864 209870 354920
rect 209926 354864 209931 354920
rect 162117 354862 209931 354864
rect 162117 354859 162183 354862
rect 209865 354859 209931 354862
rect 70894 354724 70900 354788
rect 70964 354786 70970 354788
rect 262213 354786 262279 354789
rect 70964 354784 262279 354786
rect 70964 354728 262218 354784
rect 262274 354728 262279 354784
rect 70964 354726 262279 354728
rect 70964 354724 70970 354726
rect 262213 354723 262279 354726
rect 291745 354650 291811 354653
rect 298093 354650 298159 354653
rect 291745 354648 298159 354650
rect 291745 354592 291750 354648
rect 291806 354592 298098 354648
rect 298154 354592 298159 354648
rect 291745 354590 298159 354592
rect 291745 354587 291811 354590
rect 298093 354587 298159 354590
rect 176653 354378 176719 354381
rect 295609 354378 295675 354381
rect 176653 354376 180044 354378
rect 176653 354320 176658 354376
rect 176714 354320 180044 354376
rect 176653 354318 180044 354320
rect 292836 354376 295675 354378
rect 292836 354320 295614 354376
rect 295670 354320 295675 354376
rect 292836 354318 295675 354320
rect 176653 354315 176719 354318
rect 295609 354315 295675 354318
rect 293953 352338 294019 352341
rect 292836 352336 294019 352338
rect 292836 352280 293958 352336
rect 294014 352280 294019 352336
rect 292836 352278 294019 352280
rect 293953 352275 294019 352278
rect 179462 352210 180044 352270
rect 176561 352202 176627 352205
rect 179462 352202 179522 352210
rect 176561 352200 179522 352202
rect 176561 352144 176566 352200
rect 176622 352144 179522 352200
rect 176561 352142 179522 352144
rect 176561 352139 176627 352142
rect 179505 351930 179571 351933
rect 179822 351930 179828 351932
rect 179505 351928 179828 351930
rect 179505 351872 179510 351928
rect 179566 351872 179828 351928
rect 179505 351870 179828 351872
rect 179505 351867 179571 351870
rect 179822 351868 179828 351870
rect 179892 351868 179898 351932
rect 580257 351930 580323 351933
rect 583520 351930 584960 352020
rect 580257 351928 584960 351930
rect 580257 351872 580262 351928
rect 580318 351872 584960 351928
rect 580257 351870 584960 351872
rect 580257 351867 580323 351870
rect 583520 351780 584960 351870
rect 179462 350170 180044 350230
rect 175038 350100 175044 350164
rect 175108 350162 175114 350164
rect 179462 350162 179522 350170
rect 175108 350102 179522 350162
rect 175108 350100 175114 350102
rect 295374 349618 295380 349620
rect 292836 349558 295380 349618
rect 295374 349556 295380 349558
rect 295444 349556 295450 349620
rect 179462 348130 180044 348190
rect 176653 348122 176719 348125
rect 179462 348122 179522 348130
rect 176653 348120 179522 348122
rect 176653 348064 176658 348120
rect 176714 348064 179522 348120
rect 176653 348062 179522 348064
rect 176653 348059 176719 348062
rect 292622 347036 292682 347548
rect 292614 346972 292620 347036
rect 292684 346972 292690 347036
rect 293902 345538 293908 345540
rect -960 345402 480 345492
rect 292836 345478 293908 345538
rect 293902 345476 293908 345478
rect 293972 345538 293978 345540
rect 296161 345538 296227 345541
rect 293972 345536 296227 345538
rect 293972 345480 296166 345536
rect 296222 345480 296227 345536
rect 293972 345478 296227 345480
rect 293972 345476 293978 345478
rect 296161 345475 296227 345478
rect 179462 345410 180044 345470
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 156454 345068 156460 345132
rect 156524 345130 156530 345132
rect 179462 345130 179522 345410
rect 156524 345070 179522 345130
rect 156524 345068 156530 345070
rect 295333 343498 295399 343501
rect 292836 343496 295399 343498
rect 292836 343440 295338 343496
rect 295394 343440 295399 343496
rect 292836 343438 295399 343440
rect 295333 343435 295399 343438
rect 179462 343370 180044 343430
rect 176653 343362 176719 343365
rect 179462 343362 179522 343370
rect 176653 343360 179522 343362
rect 176653 343304 176658 343360
rect 176714 343304 179522 343360
rect 176653 343302 179522 343304
rect 176653 343299 176719 343302
rect 179462 341330 180044 341390
rect 176653 341322 176719 341325
rect 179462 341322 179522 341330
rect 176653 341320 179522 341322
rect 176653 341264 176658 341320
rect 176714 341264 179522 341320
rect 176653 341262 179522 341264
rect 176653 341259 176719 341262
rect 295333 340778 295399 340781
rect 292836 340776 295399 340778
rect 292836 340720 295338 340776
rect 295394 340720 295399 340776
rect 292836 340718 295399 340720
rect 295333 340715 295399 340718
rect 179462 339290 180044 339350
rect 177062 339220 177068 339284
rect 177132 339282 177138 339284
rect 179462 339282 179522 339290
rect 177132 339222 179522 339282
rect 177132 339220 177138 339222
rect 294137 338738 294203 338741
rect 292836 338736 294203 338738
rect 292836 338680 294142 338736
rect 294198 338680 294203 338736
rect 292836 338678 294203 338680
rect 294137 338675 294203 338678
rect 583520 338452 584960 338692
rect 295609 336698 295675 336701
rect 292836 336696 295675 336698
rect 292836 336640 295614 336696
rect 295670 336640 295675 336696
rect 292836 336638 295675 336640
rect 295609 336635 295675 336638
rect 179462 336570 180044 336630
rect 176469 336562 176535 336565
rect 179462 336562 179522 336570
rect 176469 336560 179522 336562
rect 176469 336504 176474 336560
rect 176530 336504 179522 336560
rect 176469 336502 179522 336504
rect 176469 336499 176535 336502
rect 177941 334658 178007 334661
rect 295425 334658 295491 334661
rect 177941 334656 179890 334658
rect 177941 334600 177946 334656
rect 178002 334600 179890 334656
rect 177941 334598 179890 334600
rect 292836 334656 295491 334658
rect 292836 334600 295430 334656
rect 295486 334600 295491 334656
rect 292836 334598 295491 334600
rect 177941 334595 178007 334598
rect 179830 334590 179890 334598
rect 295425 334595 295491 334598
rect 179830 334530 180044 334590
rect 176653 332618 176719 332621
rect 176653 332616 179890 332618
rect 176653 332560 176658 332616
rect 176714 332560 179890 332616
rect 176653 332558 179890 332560
rect 176653 332555 176719 332558
rect 179830 332550 179890 332558
rect 179830 332490 180044 332550
rect -960 332196 480 332436
rect 295333 331938 295399 331941
rect 292836 331936 295399 331938
rect 292836 331880 295338 331936
rect 295394 331880 295399 331936
rect 292836 331878 295399 331880
rect 295333 331875 295399 331878
rect 179462 330450 180044 330510
rect 174854 330380 174860 330444
rect 174924 330442 174930 330444
rect 179462 330442 179522 330450
rect 293033 330442 293099 330445
rect 174924 330382 179522 330442
rect 292806 330440 293099 330442
rect 292806 330384 293038 330440
rect 293094 330384 293099 330440
rect 292806 330382 293099 330384
rect 174924 330380 174930 330382
rect 292806 329868 292866 330382
rect 293033 330379 293099 330382
rect 294045 327858 294111 327861
rect 294413 327858 294479 327861
rect 292836 327856 294479 327858
rect 292836 327800 294050 327856
rect 294106 327800 294418 327856
rect 294474 327800 294479 327856
rect 292836 327798 294479 327800
rect 294045 327795 294111 327798
rect 294413 327795 294479 327798
rect 179462 327730 180044 327790
rect 176510 327660 176516 327724
rect 176580 327722 176586 327724
rect 179462 327722 179522 327730
rect 176580 327662 179522 327722
rect 176580 327660 176586 327662
rect 294045 325818 294111 325821
rect 292836 325816 294111 325818
rect 292836 325760 294050 325816
rect 294106 325760 294111 325816
rect 292836 325758 294111 325760
rect 294045 325755 294111 325758
rect 179505 325750 179571 325753
rect 179505 325748 180044 325750
rect 179505 325692 179510 325748
rect 179566 325692 180044 325748
rect 179505 325690 180044 325692
rect 179505 325687 179571 325690
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 179462 323650 180044 323710
rect 176326 323580 176332 323644
rect 176396 323642 176402 323644
rect 179462 323642 179522 323650
rect 176396 323582 179522 323642
rect 176396 323580 176402 323582
rect 294137 323098 294203 323101
rect 292836 323096 294203 323098
rect 292836 323040 294142 323096
rect 294198 323040 294203 323096
rect 292836 323038 294203 323040
rect 294137 323035 294203 323038
rect 179462 321610 180044 321670
rect 176653 321602 176719 321605
rect 179462 321602 179522 321610
rect 176653 321600 179522 321602
rect 176653 321544 176658 321600
rect 176714 321544 179522 321600
rect 176653 321542 179522 321544
rect 176653 321539 176719 321542
rect 295517 321058 295583 321061
rect 292836 321056 295583 321058
rect 292836 321000 295522 321056
rect 295578 321000 295583 321056
rect 292836 320998 295583 321000
rect 295517 320995 295583 320998
rect -960 319290 480 319380
rect 3417 319290 3483 319293
rect -960 319288 3483 319290
rect -960 319232 3422 319288
rect 3478 319232 3483 319288
rect -960 319230 3483 319232
rect -960 319140 480 319230
rect 3417 319227 3483 319230
rect 295517 319018 295583 319021
rect 292836 319016 295583 319018
rect 292836 318960 295522 319016
rect 295578 318960 295583 319016
rect 292836 318958 295583 318960
rect 295517 318955 295583 318958
rect 179462 318890 180044 318950
rect 177757 318882 177823 318885
rect 179462 318882 179522 318890
rect 177757 318880 179522 318882
rect 177757 318824 177762 318880
rect 177818 318824 179522 318880
rect 177757 318822 179522 318824
rect 177757 318819 177823 318822
rect 295609 316978 295675 316981
rect 292836 316976 295675 316978
rect 292836 316920 295614 316976
rect 295670 316920 295675 316976
rect 292836 316918 295675 316920
rect 295609 316915 295675 316918
rect 179505 316910 179571 316913
rect 179505 316908 180044 316910
rect 179505 316852 179510 316908
rect 179566 316852 180044 316908
rect 179505 316850 180044 316852
rect 179505 316847 179571 316850
rect 179462 314810 180044 314870
rect 176653 314802 176719 314805
rect 179462 314802 179522 314810
rect 176653 314800 179522 314802
rect 176653 314744 176658 314800
rect 176714 314744 179522 314800
rect 176653 314742 179522 314744
rect 176653 314739 176719 314742
rect 295517 314258 295583 314261
rect 292836 314256 295583 314258
rect 292836 314200 295522 314256
rect 295578 314200 295583 314256
rect 292836 314198 295583 314200
rect 295517 314195 295583 314198
rect 179830 312770 180044 312830
rect 178953 312762 179019 312765
rect 179830 312762 179890 312770
rect 178953 312760 179890 312762
rect 178953 312704 178958 312760
rect 179014 312704 179890 312760
rect 178953 312702 179890 312704
rect 178953 312699 179019 312702
rect 295517 312218 295583 312221
rect 292836 312216 295583 312218
rect 292836 312160 295522 312216
rect 295578 312160 295583 312216
rect 292836 312158 295583 312160
rect 295517 312155 295583 312158
rect 580349 312082 580415 312085
rect 583520 312082 584960 312172
rect 580349 312080 584960 312082
rect 580349 312024 580354 312080
rect 580410 312024 584960 312080
rect 580349 312022 584960 312024
rect 580349 312019 580415 312022
rect 583520 311932 584960 312022
rect 295517 310178 295583 310181
rect 292836 310176 295583 310178
rect 292836 310120 295522 310176
rect 295578 310120 295583 310176
rect 292836 310118 295583 310120
rect 295517 310115 295583 310118
rect 179462 310050 180044 310110
rect 176653 310042 176719 310045
rect 179462 310042 179522 310050
rect 176653 310040 179522 310042
rect 176653 309984 176658 310040
rect 176714 309984 179522 310040
rect 176653 309982 179522 309984
rect 176653 309979 176719 309982
rect 295517 308138 295583 308141
rect 292836 308136 295583 308138
rect 292836 308080 295522 308136
rect 295578 308080 295583 308136
rect 292836 308078 295583 308080
rect 295517 308075 295583 308078
rect 179462 308010 180044 308070
rect 176653 308002 176719 308005
rect 179462 308002 179522 308010
rect 176653 308000 179522 308002
rect 176653 307944 176658 308000
rect 176714 307944 179522 308000
rect 176653 307942 179522 307944
rect 176653 307939 176719 307942
rect -960 306234 480 306324
rect 3233 306234 3299 306237
rect -960 306232 3299 306234
rect -960 306176 3238 306232
rect 3294 306176 3299 306232
rect -960 306174 3299 306176
rect -960 306084 480 306174
rect 3233 306171 3299 306174
rect 179462 305970 180044 306030
rect 176653 305962 176719 305965
rect 179462 305962 179522 305970
rect 176653 305960 179522 305962
rect 176653 305904 176658 305960
rect 176714 305904 179522 305960
rect 176653 305902 179522 305904
rect 176653 305899 176719 305902
rect 295425 305418 295491 305421
rect 292836 305416 295491 305418
rect 292836 305360 295430 305416
rect 295486 305360 295491 305416
rect 292836 305358 295491 305360
rect 295425 305355 295491 305358
rect 179462 303930 180044 303990
rect 177941 303922 178007 303925
rect 179462 303922 179522 303930
rect 177941 303920 179522 303922
rect 177941 303864 177946 303920
rect 178002 303864 179522 303920
rect 177941 303862 179522 303864
rect 177941 303859 178007 303862
rect 294229 303378 294295 303381
rect 292836 303376 294295 303378
rect 292836 303320 294234 303376
rect 294290 303320 294295 303376
rect 292836 303318 294295 303320
rect 294229 303315 294295 303318
rect 293125 301338 293191 301341
rect 292836 301336 293191 301338
rect 292836 301280 293130 301336
rect 293186 301280 293191 301336
rect 292836 301278 293191 301280
rect 293125 301275 293191 301278
rect 179462 301210 180044 301270
rect 177665 301202 177731 301205
rect 179462 301202 179522 301210
rect 177665 301200 179522 301202
rect 177665 301144 177670 301200
rect 177726 301144 179522 301200
rect 177665 301142 179522 301144
rect 177665 301139 177731 301142
rect 76097 300930 76163 300933
rect 155401 300930 155467 300933
rect 76097 300928 155467 300930
rect 76097 300872 76102 300928
rect 76158 300872 155406 300928
rect 155462 300872 155467 300928
rect 76097 300870 155467 300872
rect 76097 300867 76163 300870
rect 155401 300867 155467 300870
rect 84377 299570 84443 299573
rect 154021 299570 154087 299573
rect 84377 299568 154087 299570
rect 84377 299512 84382 299568
rect 84438 299512 154026 299568
rect 154082 299512 154087 299568
rect 84377 299510 154087 299512
rect 84377 299507 84443 299510
rect 154021 299507 154087 299510
rect 176653 299298 176719 299301
rect 296621 299298 296687 299301
rect 176653 299296 179522 299298
rect 176653 299240 176658 299296
rect 176714 299240 179522 299296
rect 176653 299238 179522 299240
rect 292836 299296 296687 299298
rect 292836 299240 296626 299296
rect 296682 299240 296687 299296
rect 292836 299238 296687 299240
rect 176653 299235 176719 299238
rect 179462 299230 179522 299238
rect 296621 299235 296687 299238
rect 179462 299170 180044 299230
rect 57881 298754 57947 298757
rect 166441 298754 166507 298757
rect 57881 298752 166507 298754
rect 57881 298696 57886 298752
rect 57942 298696 166446 298752
rect 166502 298696 166507 298752
rect 57881 298694 166507 298696
rect 57881 298691 57947 298694
rect 166441 298691 166507 298694
rect 579613 298754 579679 298757
rect 583520 298754 584960 298844
rect 579613 298752 584960 298754
rect 579613 298696 579618 298752
rect 579674 298696 584960 298752
rect 579613 298694 584960 298696
rect 579613 298691 579679 298694
rect 583520 298604 584960 298694
rect 89345 298210 89411 298213
rect 131849 298210 131915 298213
rect 89345 298208 131915 298210
rect 89345 298152 89350 298208
rect 89406 298152 131854 298208
rect 131910 298152 131915 298208
rect 89345 298150 131915 298152
rect 89345 298147 89411 298150
rect 131849 298147 131915 298150
rect 104893 297394 104959 297397
rect 157333 297394 157399 297397
rect 104893 297392 157399 297394
rect 104893 297336 104898 297392
rect 104954 297336 157338 297392
rect 157394 297336 157399 297392
rect 104893 297334 157399 297336
rect 104893 297331 104959 297334
rect 157333 297331 157399 297334
rect 176653 297258 176719 297261
rect 176653 297256 179522 297258
rect 176653 297200 176658 297256
rect 176714 297200 179522 297256
rect 176653 297198 179522 297200
rect 176653 297195 176719 297198
rect 179462 297190 179522 297198
rect 179462 297130 180044 297190
rect 68737 296850 68803 296853
rect 170254 296850 170260 296852
rect 68737 296848 170260 296850
rect 68737 296792 68742 296848
rect 68798 296792 170260 296848
rect 68737 296790 170260 296792
rect 68737 296787 68803 296790
rect 170254 296788 170260 296790
rect 170324 296788 170330 296852
rect 295425 296578 295491 296581
rect 292836 296576 295491 296578
rect 292836 296520 295430 296576
rect 295486 296520 295491 296576
rect 292836 296518 295491 296520
rect 295425 296515 295491 296518
rect 95141 296034 95207 296037
rect 104893 296034 104959 296037
rect 95141 296032 104959 296034
rect 95141 295976 95146 296032
rect 95202 295976 104898 296032
rect 104954 295976 104959 296032
rect 95141 295974 104959 295976
rect 95141 295971 95207 295974
rect 104893 295971 104959 295974
rect 106089 295354 106155 295357
rect 171910 295354 171916 295356
rect 106089 295352 171916 295354
rect 106089 295296 106094 295352
rect 106150 295296 171916 295352
rect 106089 295294 171916 295296
rect 106089 295291 106155 295294
rect 171910 295292 171916 295294
rect 171980 295292 171986 295356
rect 179462 295090 180044 295150
rect 176653 295082 176719 295085
rect 179462 295082 179522 295090
rect 176653 295080 179522 295082
rect 176653 295024 176658 295080
rect 176714 295024 179522 295080
rect 176653 295022 179522 295024
rect 176653 295019 176719 295022
rect 295333 294538 295399 294541
rect 292836 294536 295399 294538
rect 292836 294480 295338 294536
rect 295394 294480 295399 294536
rect 292836 294478 295399 294480
rect 295333 294475 295399 294478
rect 108021 294266 108087 294269
rect 119654 294266 119660 294268
rect 108021 294264 119660 294266
rect 108021 294208 108026 294264
rect 108082 294208 119660 294264
rect 108021 294206 119660 294208
rect 108021 294203 108087 294206
rect 119654 294204 119660 294206
rect 119724 294204 119730 294268
rect 96429 294130 96495 294133
rect 84150 294128 96495 294130
rect 84150 294072 96434 294128
rect 96490 294072 96495 294128
rect 84150 294070 96495 294072
rect 35801 293994 35867 293997
rect 84150 293994 84210 294070
rect 96429 294067 96495 294070
rect 114461 294130 114527 294133
rect 141509 294130 141575 294133
rect 114461 294128 141575 294130
rect 114461 294072 114466 294128
rect 114522 294072 141514 294128
rect 141570 294072 141575 294128
rect 114461 294070 141575 294072
rect 114461 294067 114527 294070
rect 141509 294067 141575 294070
rect 35801 293992 84210 293994
rect 35801 293936 35806 293992
rect 35862 293936 84210 293992
rect 35801 293934 84210 293936
rect 95785 293994 95851 293997
rect 173157 293994 173223 293997
rect 95785 293992 173223 293994
rect 95785 293936 95790 293992
rect 95846 293936 173162 293992
rect 173218 293936 173223 293992
rect 95785 293934 173223 293936
rect 35801 293931 35867 293934
rect 95785 293931 95851 293934
rect 173157 293931 173223 293934
rect -960 293178 480 293268
rect 3325 293178 3391 293181
rect -960 293176 3391 293178
rect -960 293120 3330 293176
rect 3386 293120 3391 293176
rect -960 293118 3391 293120
rect -960 293028 480 293118
rect 3325 293115 3391 293118
rect 73889 292906 73955 292909
rect 119286 292906 119292 292908
rect 73889 292904 119292 292906
rect 73889 292848 73894 292904
rect 73950 292848 119292 292904
rect 73889 292846 119292 292848
rect 73889 292843 73955 292846
rect 119286 292844 119292 292846
rect 119356 292844 119362 292908
rect 77753 292770 77819 292773
rect 125133 292770 125199 292773
rect 77753 292768 125199 292770
rect 77753 292712 77758 292768
rect 77814 292712 125138 292768
rect 125194 292712 125199 292768
rect 77753 292710 125199 292712
rect 77753 292707 77819 292710
rect 125133 292707 125199 292710
rect 78397 292634 78463 292637
rect 176009 292634 176075 292637
rect 78397 292632 176075 292634
rect 78397 292576 78402 292632
rect 78458 292576 176014 292632
rect 176070 292576 176075 292632
rect 78397 292574 176075 292576
rect 78397 292571 78463 292574
rect 176009 292571 176075 292574
rect 295609 292498 295675 292501
rect 292836 292496 295675 292498
rect 292836 292440 295614 292496
rect 295670 292440 295675 292496
rect 292836 292438 295675 292440
rect 295609 292435 295675 292438
rect 179462 292370 180044 292430
rect 71681 292362 71747 292365
rect 70718 292360 71747 292362
rect 70718 292304 71686 292360
rect 71742 292304 71747 292360
rect 70718 292302 71747 292304
rect 70718 291788 70778 292302
rect 71681 292299 71747 292302
rect 176653 292362 176719 292365
rect 179462 292362 179522 292370
rect 176653 292360 179522 292362
rect 176653 292304 176658 292360
rect 176714 292304 179522 292360
rect 176653 292302 179522 292304
rect 176653 292299 176719 292302
rect 117773 291954 117839 291957
rect 160829 291954 160895 291957
rect 117773 291952 160895 291954
rect 117773 291896 117778 291952
rect 117834 291896 160834 291952
rect 160890 291896 160895 291952
rect 117773 291894 160895 291896
rect 117773 291891 117839 291894
rect 160829 291891 160895 291894
rect 121545 291818 121611 291821
rect 119876 291816 121611 291818
rect 119876 291760 121550 291816
rect 121606 291760 121611 291816
rect 119876 291758 121611 291760
rect 121545 291755 121611 291758
rect 67725 291138 67791 291141
rect 121637 291138 121703 291141
rect 67725 291136 70196 291138
rect 67725 291080 67730 291136
rect 67786 291080 70196 291136
rect 67725 291078 70196 291080
rect 119876 291136 121703 291138
rect 119876 291080 121642 291136
rect 121698 291080 121703 291136
rect 119876 291078 121703 291080
rect 67725 291075 67791 291078
rect 121637 291075 121703 291078
rect 67633 290458 67699 290461
rect 121545 290458 121611 290461
rect 295517 290458 295583 290461
rect 67633 290456 70196 290458
rect 67633 290400 67638 290456
rect 67694 290400 70196 290456
rect 67633 290398 70196 290400
rect 119876 290456 121611 290458
rect 119876 290400 121550 290456
rect 121606 290400 121611 290456
rect 119876 290398 121611 290400
rect 292836 290456 295583 290458
rect 292836 290400 295522 290456
rect 295578 290400 295583 290456
rect 292836 290398 295583 290400
rect 67633 290395 67699 290398
rect 121545 290395 121611 290398
rect 295517 290395 295583 290398
rect 179462 290330 180044 290390
rect 176653 290322 176719 290325
rect 179462 290322 179522 290330
rect 176653 290320 179522 290322
rect 176653 290264 176658 290320
rect 176714 290264 179522 290320
rect 176653 290262 179522 290264
rect 176653 290259 176719 290262
rect 121545 289778 121611 289781
rect 119876 289776 121611 289778
rect 70166 289234 70226 289748
rect 119876 289720 121550 289776
rect 121606 289720 121611 289776
rect 119876 289718 121611 289720
rect 121545 289715 121611 289718
rect 64830 289174 70226 289234
rect 64638 288628 64644 288692
rect 64708 288690 64714 288692
rect 64830 288690 64890 289174
rect 119654 289172 119660 289236
rect 119724 289234 119730 289236
rect 152549 289234 152615 289237
rect 119724 289232 152615 289234
rect 119724 289176 152554 289232
rect 152610 289176 152615 289232
rect 119724 289174 152615 289176
rect 119724 289172 119730 289174
rect 152549 289171 152615 289174
rect 67633 289098 67699 289101
rect 121545 289098 121611 289101
rect 67633 289096 70196 289098
rect 67633 289040 67638 289096
rect 67694 289040 70196 289096
rect 67633 289038 70196 289040
rect 119876 289096 121611 289098
rect 119876 289040 121550 289096
rect 121606 289040 121611 289096
rect 119876 289038 121611 289040
rect 67633 289035 67699 289038
rect 121545 289035 121611 289038
rect 64708 288630 64890 288690
rect 64708 288628 64714 288630
rect 68369 288418 68435 288421
rect 121729 288418 121795 288421
rect 68369 288416 70196 288418
rect 68369 288360 68374 288416
rect 68430 288360 70196 288416
rect 68369 288358 70196 288360
rect 119876 288416 121795 288418
rect 119876 288360 121734 288416
rect 121790 288360 121795 288416
rect 119876 288358 121795 288360
rect 68369 288355 68435 288358
rect 121729 288355 121795 288358
rect 179462 288290 180044 288350
rect 179229 288282 179295 288285
rect 179462 288282 179522 288290
rect 161430 288280 179522 288282
rect 161430 288224 179234 288280
rect 179290 288224 179522 288280
rect 161430 288222 179522 288224
rect 119286 288084 119292 288148
rect 119356 288146 119362 288148
rect 161430 288146 161490 288222
rect 179229 288219 179295 288222
rect 119356 288086 161490 288146
rect 119356 288084 119362 288086
rect 67633 287738 67699 287741
rect 121637 287738 121703 287741
rect 67633 287736 70196 287738
rect 67633 287680 67638 287736
rect 67694 287680 70196 287736
rect 67633 287678 70196 287680
rect 119876 287736 121703 287738
rect 119876 287680 121642 287736
rect 121698 287680 121703 287736
rect 119876 287678 121703 287680
rect 67633 287675 67699 287678
rect 121637 287675 121703 287678
rect 292806 287466 292866 287708
rect 293033 287466 293099 287469
rect 292806 287464 293099 287466
rect 292806 287408 293038 287464
rect 293094 287408 293099 287464
rect 292806 287406 293099 287408
rect 293033 287403 293099 287406
rect 67725 287058 67791 287061
rect 122741 287058 122807 287061
rect 67725 287056 70196 287058
rect 67725 287000 67730 287056
rect 67786 287000 70196 287056
rect 67725 286998 70196 287000
rect 119876 287056 122807 287058
rect 119876 287000 122746 287056
rect 122802 287000 122807 287056
rect 119876 286998 122807 287000
rect 67725 286995 67791 286998
rect 122741 286995 122807 286998
rect 67541 286378 67607 286381
rect 120165 286378 120231 286381
rect 67541 286376 70196 286378
rect 67541 286320 67546 286376
rect 67602 286320 70196 286376
rect 67541 286318 70196 286320
rect 119876 286376 120231 286378
rect 119876 286320 120170 286376
rect 120226 286320 120231 286376
rect 119876 286318 120231 286320
rect 67541 286315 67607 286318
rect 120165 286315 120231 286318
rect 177849 286378 177915 286381
rect 177849 286376 179890 286378
rect 177849 286320 177854 286376
rect 177910 286320 179890 286376
rect 177849 286318 179890 286320
rect 177849 286315 177915 286318
rect 179830 286310 179890 286318
rect 179830 286250 180044 286310
rect 67633 285698 67699 285701
rect 121453 285698 121519 285701
rect 295517 285698 295583 285701
rect 67633 285696 70196 285698
rect 67633 285640 67638 285696
rect 67694 285640 70196 285696
rect 67633 285638 70196 285640
rect 119876 285696 121519 285698
rect 119876 285640 121458 285696
rect 121514 285640 121519 285696
rect 119876 285638 121519 285640
rect 292836 285696 295583 285698
rect 292836 285640 295522 285696
rect 295578 285640 295583 285696
rect 292836 285638 295583 285640
rect 67633 285635 67699 285638
rect 121453 285635 121519 285638
rect 295517 285635 295583 285638
rect 583520 285276 584960 285516
rect 68553 285018 68619 285021
rect 121453 285018 121519 285021
rect 68553 285016 70196 285018
rect 68553 284960 68558 285016
rect 68614 284960 70196 285016
rect 68553 284958 70196 284960
rect 119876 285016 121519 285018
rect 119876 284960 121458 285016
rect 121514 284960 121519 285016
rect 119876 284958 121519 284960
rect 68553 284955 68619 284958
rect 121453 284955 121519 284958
rect 68277 284338 68343 284341
rect 121545 284338 121611 284341
rect 68277 284336 70196 284338
rect 68277 284280 68282 284336
rect 68338 284280 70196 284336
rect 68277 284278 70196 284280
rect 119876 284336 121611 284338
rect 119876 284280 121550 284336
rect 121606 284280 121611 284336
rect 119876 284278 121611 284280
rect 68277 284275 68343 284278
rect 121545 284275 121611 284278
rect 125133 284202 125199 284205
rect 125133 284200 161490 284202
rect 125133 284144 125138 284200
rect 125194 284144 161490 284200
rect 125133 284142 161490 284144
rect 125133 284139 125199 284142
rect 68461 283658 68527 283661
rect 121453 283658 121519 283661
rect 68461 283656 70196 283658
rect 68461 283600 68466 283656
rect 68522 283600 70196 283656
rect 68461 283598 70196 283600
rect 119876 283656 121519 283658
rect 119876 283600 121458 283656
rect 121514 283600 121519 283656
rect 119876 283598 121519 283600
rect 161430 283658 161490 284142
rect 179270 283658 179276 283660
rect 161430 283598 179276 283658
rect 68461 283595 68527 283598
rect 121453 283595 121519 283598
rect 179270 283596 179276 283598
rect 179340 283658 179346 283660
rect 295517 283658 295583 283661
rect 179340 283598 179522 283658
rect 292836 283656 295583 283658
rect 292836 283600 295522 283656
rect 295578 283600 295583 283656
rect 292836 283598 295583 283600
rect 179340 283596 179346 283598
rect 179462 283590 179522 283598
rect 295517 283595 295583 283598
rect 179462 283530 180044 283590
rect 67633 282978 67699 282981
rect 121729 282978 121795 282981
rect 67633 282976 70196 282978
rect 67633 282920 67638 282976
rect 67694 282920 70196 282976
rect 67633 282918 70196 282920
rect 119876 282976 121795 282978
rect 119876 282920 121734 282976
rect 121790 282920 121795 282976
rect 119876 282918 121795 282920
rect 67633 282915 67699 282918
rect 121729 282915 121795 282918
rect 121545 282298 121611 282301
rect 119876 282296 121611 282298
rect 119876 282240 121550 282296
rect 121606 282240 121611 282296
rect 119876 282238 121611 282240
rect 121545 282235 121611 282238
rect 67633 281618 67699 281621
rect 121453 281618 121519 281621
rect 67633 281616 70196 281618
rect 67633 281560 67638 281616
rect 67694 281560 70196 281616
rect 67633 281558 70196 281560
rect 119876 281616 121519 281618
rect 119876 281560 121458 281616
rect 121514 281560 121519 281616
rect 119876 281558 121519 281560
rect 67633 281555 67699 281558
rect 121453 281555 121519 281558
rect 176653 281618 176719 281621
rect 293902 281618 293908 281620
rect 176653 281616 179522 281618
rect 176653 281560 176658 281616
rect 176714 281560 179522 281616
rect 176653 281558 179522 281560
rect 292836 281558 293908 281618
rect 176653 281555 176719 281558
rect 179462 281550 179522 281558
rect 293902 281556 293908 281558
rect 293972 281618 293978 281620
rect 295517 281618 295583 281621
rect 293972 281616 295583 281618
rect 293972 281560 295522 281616
rect 295578 281560 295583 281616
rect 293972 281558 295583 281560
rect 293972 281556 293978 281558
rect 295517 281555 295583 281558
rect 179462 281490 180044 281550
rect 67725 280938 67791 280941
rect 121545 280938 121611 280941
rect 67725 280936 70196 280938
rect 67725 280880 67730 280936
rect 67786 280880 70196 280936
rect 67725 280878 70196 280880
rect 119876 280936 121611 280938
rect 119876 280880 121550 280936
rect 121606 280880 121611 280936
rect 119876 280878 121611 280880
rect 67725 280875 67791 280878
rect 121545 280875 121611 280878
rect 67633 280258 67699 280261
rect 121453 280258 121519 280261
rect 67633 280256 70196 280258
rect -960 279972 480 280212
rect 67633 280200 67638 280256
rect 67694 280200 70196 280256
rect 67633 280198 70196 280200
rect 119876 280256 121519 280258
rect 119876 280200 121458 280256
rect 121514 280200 121519 280256
rect 119876 280198 121519 280200
rect 67633 280195 67699 280198
rect 121453 280195 121519 280198
rect 67909 279578 67975 279581
rect 68829 279578 68895 279581
rect 122281 279578 122347 279581
rect 67909 279576 70196 279578
rect 67909 279520 67914 279576
rect 67970 279520 68834 279576
rect 68890 279520 70196 279576
rect 67909 279518 70196 279520
rect 119876 279576 122347 279578
rect 119876 279520 122286 279576
rect 122342 279520 122347 279576
rect 119876 279518 122347 279520
rect 67909 279515 67975 279518
rect 68829 279515 68895 279518
rect 122281 279515 122347 279518
rect 176745 279578 176811 279581
rect 179045 279578 179111 279581
rect 176745 279576 179890 279578
rect 176745 279520 176750 279576
rect 176806 279520 179050 279576
rect 179106 279520 179890 279576
rect 176745 279518 179890 279520
rect 176745 279515 176811 279518
rect 179045 279515 179111 279518
rect 179830 279510 179890 279518
rect 179830 279450 180044 279510
rect 57830 278836 57836 278900
rect 57900 278898 57906 278900
rect 121453 278898 121519 278901
rect 295517 278898 295583 278901
rect 57900 278838 70196 278898
rect 119876 278896 121519 278898
rect 119876 278840 121458 278896
rect 121514 278840 121519 278896
rect 119876 278838 121519 278840
rect 292836 278896 295583 278898
rect 292836 278840 295522 278896
rect 295578 278840 295583 278896
rect 292836 278838 295583 278840
rect 57900 278836 57906 278838
rect 121453 278835 121519 278838
rect 295517 278835 295583 278838
rect 67725 278218 67791 278221
rect 122189 278218 122255 278221
rect 67725 278216 70196 278218
rect 67725 278160 67730 278216
rect 67786 278160 70196 278216
rect 67725 278158 70196 278160
rect 119876 278216 122255 278218
rect 119876 278160 122194 278216
rect 122250 278160 122255 278216
rect 119876 278158 122255 278160
rect 67725 278155 67791 278158
rect 122189 278155 122255 278158
rect 67633 277538 67699 277541
rect 121453 277538 121519 277541
rect 67633 277536 70196 277538
rect 67633 277480 67638 277536
rect 67694 277480 70196 277536
rect 67633 277478 70196 277480
rect 119876 277536 121519 277538
rect 119876 277480 121458 277536
rect 121514 277480 121519 277536
rect 119876 277478 121519 277480
rect 67633 277475 67699 277478
rect 121453 277475 121519 277478
rect 176653 277538 176719 277541
rect 176653 277536 179522 277538
rect 176653 277480 176658 277536
rect 176714 277480 179522 277536
rect 176653 277478 179522 277480
rect 176653 277475 176719 277478
rect 179462 277470 179522 277478
rect 179462 277410 180044 277470
rect 67725 276858 67791 276861
rect 121545 276858 121611 276861
rect 295609 276858 295675 276861
rect 67725 276856 70196 276858
rect 67725 276800 67730 276856
rect 67786 276800 70196 276856
rect 67725 276798 70196 276800
rect 119876 276856 121611 276858
rect 119876 276800 121550 276856
rect 121606 276800 121611 276856
rect 119876 276798 121611 276800
rect 292836 276856 295675 276858
rect 292836 276800 295614 276856
rect 295670 276800 295675 276856
rect 292836 276798 295675 276800
rect 67725 276795 67791 276798
rect 121545 276795 121611 276798
rect 295609 276795 295675 276798
rect 67633 276178 67699 276181
rect 121453 276178 121519 276181
rect 67633 276176 70196 276178
rect 67633 276120 67638 276176
rect 67694 276120 70196 276176
rect 67633 276118 70196 276120
rect 119876 276176 121519 276178
rect 119876 276120 121458 276176
rect 121514 276120 121519 276176
rect 119876 276118 121519 276120
rect 67633 276115 67699 276118
rect 121453 276115 121519 276118
rect 68921 275498 68987 275501
rect 121545 275498 121611 275501
rect 68921 275496 70196 275498
rect 68921 275440 68926 275496
rect 68982 275440 70196 275496
rect 68921 275438 70196 275440
rect 119876 275496 121611 275498
rect 119876 275440 121550 275496
rect 121606 275440 121611 275496
rect 119876 275438 121611 275440
rect 68921 275435 68987 275438
rect 121545 275435 121611 275438
rect 67633 274818 67699 274821
rect 121453 274818 121519 274821
rect 67633 274816 70196 274818
rect 67633 274760 67638 274816
rect 67694 274760 70196 274816
rect 67633 274758 70196 274760
rect 119876 274816 121519 274818
rect 119876 274760 121458 274816
rect 121514 274760 121519 274816
rect 119876 274758 121519 274760
rect 67633 274755 67699 274758
rect 121453 274755 121519 274758
rect 176653 274818 176719 274821
rect 295701 274818 295767 274821
rect 176653 274816 179522 274818
rect 176653 274760 176658 274816
rect 176714 274760 179522 274816
rect 176653 274758 179522 274760
rect 292836 274816 295767 274818
rect 292836 274760 295706 274816
rect 295762 274760 295767 274816
rect 292836 274758 295767 274760
rect 176653 274755 176719 274758
rect 179462 274750 179522 274758
rect 295701 274755 295767 274758
rect 179462 274690 180044 274750
rect 67725 274138 67791 274141
rect 121453 274138 121519 274141
rect 67725 274136 70196 274138
rect 67725 274080 67730 274136
rect 67786 274080 70196 274136
rect 67725 274078 70196 274080
rect 119876 274136 121519 274138
rect 119876 274080 121458 274136
rect 121514 274080 121519 274136
rect 119876 274078 121519 274080
rect 67725 274075 67791 274078
rect 121453 274075 121519 274078
rect 67633 273458 67699 273461
rect 121453 273458 121519 273461
rect 67633 273456 70196 273458
rect 67633 273400 67638 273456
rect 67694 273400 70196 273456
rect 67633 273398 70196 273400
rect 119876 273456 121519 273458
rect 119876 273400 121458 273456
rect 121514 273400 121519 273456
rect 119876 273398 121519 273400
rect 67633 273395 67699 273398
rect 121453 273395 121519 273398
rect 67725 272778 67791 272781
rect 121637 272778 121703 272781
rect 122097 272778 122163 272781
rect 67725 272776 70196 272778
rect 67725 272720 67730 272776
rect 67786 272720 70196 272776
rect 67725 272718 70196 272720
rect 119876 272776 122163 272778
rect 119876 272720 121642 272776
rect 121698 272720 122102 272776
rect 122158 272720 122163 272776
rect 119876 272718 122163 272720
rect 67725 272715 67791 272718
rect 121637 272715 121703 272718
rect 122097 272715 122163 272718
rect 176653 272778 176719 272781
rect 295609 272778 295675 272781
rect 176653 272776 179522 272778
rect 176653 272720 176658 272776
rect 176714 272720 179522 272776
rect 176653 272718 179522 272720
rect 292836 272776 295675 272778
rect 292836 272720 295614 272776
rect 295670 272720 295675 272776
rect 292836 272718 295675 272720
rect 176653 272715 176719 272718
rect 179462 272710 179522 272718
rect 295609 272715 295675 272718
rect 179462 272650 180044 272710
rect 580349 272234 580415 272237
rect 583520 272234 584960 272324
rect 580349 272232 584960 272234
rect 580349 272176 580354 272232
rect 580410 272176 584960 272232
rect 580349 272174 584960 272176
rect 580349 272171 580415 272174
rect 67633 272098 67699 272101
rect 121453 272098 121519 272101
rect 67633 272096 70196 272098
rect 67633 272040 67638 272096
rect 67694 272040 70196 272096
rect 67633 272038 70196 272040
rect 119876 272096 121519 272098
rect 119876 272040 121458 272096
rect 121514 272040 121519 272096
rect 583520 272084 584960 272174
rect 119876 272038 121519 272040
rect 67633 272035 67699 272038
rect 121453 272035 121519 272038
rect 59118 271900 59124 271964
rect 59188 271962 59194 271964
rect 62297 271962 62363 271965
rect 59188 271960 62363 271962
rect 59188 271904 62302 271960
rect 62358 271904 62363 271960
rect 59188 271902 62363 271904
rect 59188 271900 59194 271902
rect 62297 271899 62363 271902
rect 67633 271418 67699 271421
rect 121453 271418 121519 271421
rect 67633 271416 70196 271418
rect 67633 271360 67638 271416
rect 67694 271360 70196 271416
rect 67633 271358 70196 271360
rect 119876 271416 121519 271418
rect 119876 271360 121458 271416
rect 121514 271360 121519 271416
rect 119876 271358 121519 271360
rect 67633 271355 67699 271358
rect 121453 271355 121519 271358
rect 67725 270738 67791 270741
rect 67725 270736 70196 270738
rect 67725 270680 67730 270736
rect 67786 270680 70196 270736
rect 67725 270678 70196 270680
rect 67725 270675 67791 270678
rect 179462 270610 180044 270670
rect 177849 270602 177915 270605
rect 179462 270602 179522 270610
rect 177849 270600 179522 270602
rect 177849 270544 177854 270600
rect 177910 270544 179522 270600
rect 177849 270542 179522 270544
rect 177849 270539 177915 270542
rect 67633 270058 67699 270061
rect 121545 270058 121611 270061
rect 295609 270058 295675 270061
rect 67633 270056 70196 270058
rect 67633 270000 67638 270056
rect 67694 270000 70196 270056
rect 67633 269998 70196 270000
rect 119876 270056 121611 270058
rect 119876 270000 121550 270056
rect 121606 270000 121611 270056
rect 119876 269998 121611 270000
rect 292836 270056 295675 270058
rect 292836 270000 295614 270056
rect 295670 270000 295675 270056
rect 292836 269998 295675 270000
rect 67633 269995 67699 269998
rect 121545 269995 121611 269998
rect 295609 269995 295675 269998
rect 68185 269378 68251 269381
rect 121453 269378 121519 269381
rect 68185 269376 70196 269378
rect 68185 269320 68190 269376
rect 68246 269320 70196 269376
rect 68185 269318 70196 269320
rect 119876 269376 121519 269378
rect 119876 269320 121458 269376
rect 121514 269320 121519 269376
rect 119876 269318 121519 269320
rect 68185 269315 68251 269318
rect 121453 269315 121519 269318
rect 68185 268698 68251 268701
rect 120073 268698 120139 268701
rect 68185 268696 70196 268698
rect 68185 268640 68190 268696
rect 68246 268640 70196 268696
rect 68185 268638 70196 268640
rect 119876 268696 120139 268698
rect 119876 268640 120078 268696
rect 120134 268640 120139 268696
rect 119876 268638 120139 268640
rect 68185 268635 68251 268638
rect 120073 268635 120139 268638
rect 179462 268570 180044 268630
rect 176653 268562 176719 268565
rect 179462 268562 179522 268570
rect 176653 268560 179522 268562
rect 176653 268504 176658 268560
rect 176714 268504 179522 268560
rect 176653 268502 179522 268504
rect 176653 268499 176719 268502
rect 67633 268018 67699 268021
rect 121453 268018 121519 268021
rect 294229 268018 294295 268021
rect 67633 268016 70196 268018
rect 67633 267960 67638 268016
rect 67694 267960 70196 268016
rect 67633 267958 70196 267960
rect 119876 268016 121519 268018
rect 119876 267960 121458 268016
rect 121514 267960 121519 268016
rect 119876 267958 121519 267960
rect 292836 268016 294295 268018
rect 292836 267960 294234 268016
rect 294290 267960 294295 268016
rect 292836 267958 294295 267960
rect 67633 267955 67699 267958
rect 121453 267955 121519 267958
rect 294229 267955 294295 267958
rect 70526 267474 70532 267476
rect 70350 267414 70532 267474
rect 70350 267338 70410 267414
rect 70526 267412 70532 267414
rect 70596 267412 70602 267476
rect 121545 267338 121611 267341
rect 70196 267308 70410 267338
rect 119876 267336 121611 267338
rect -960 267202 480 267292
rect 70166 267278 70380 267308
rect 119876 267280 121550 267336
rect 121606 267280 121611 267336
rect 119876 267278 121611 267280
rect 3049 267202 3115 267205
rect -960 267200 3115 267202
rect -960 267144 3054 267200
rect 3110 267144 3115 267200
rect -960 267142 3115 267144
rect -960 267052 480 267142
rect 3049 267139 3115 267142
rect 70166 266794 70226 267278
rect 121545 267275 121611 267278
rect 64830 266734 70226 266794
rect 21357 266386 21423 266389
rect 64830 266386 64890 266734
rect 67633 266658 67699 266661
rect 121453 266658 121519 266661
rect 67633 266656 70196 266658
rect 67633 266600 67638 266656
rect 67694 266600 70196 266656
rect 67633 266598 70196 266600
rect 119876 266656 121519 266658
rect 119876 266600 121458 266656
rect 121514 266600 121519 266656
rect 119876 266598 121519 266600
rect 67633 266595 67699 266598
rect 121453 266595 121519 266598
rect 21357 266384 64890 266386
rect 21357 266328 21362 266384
rect 21418 266328 64890 266384
rect 21357 266326 64890 266328
rect 21357 266323 21423 266326
rect 67633 265978 67699 265981
rect 121545 265978 121611 265981
rect 67633 265976 70196 265978
rect 67633 265920 67638 265976
rect 67694 265920 70196 265976
rect 67633 265918 70196 265920
rect 119876 265976 121611 265978
rect 119876 265920 121550 265976
rect 121606 265920 121611 265976
rect 119876 265918 121611 265920
rect 67633 265915 67699 265918
rect 121545 265915 121611 265918
rect 176653 265978 176719 265981
rect 295609 265978 295675 265981
rect 176653 265976 179522 265978
rect 176653 265920 176658 265976
rect 176714 265920 179522 265976
rect 176653 265918 179522 265920
rect 292836 265976 295675 265978
rect 292836 265920 295614 265976
rect 295670 265920 295675 265976
rect 292836 265918 295675 265920
rect 176653 265915 176719 265918
rect 179462 265910 179522 265918
rect 295609 265915 295675 265918
rect 179462 265850 180044 265910
rect 67725 265298 67791 265301
rect 121453 265298 121519 265301
rect 67725 265296 70196 265298
rect 67725 265240 67730 265296
rect 67786 265240 70196 265296
rect 67725 265238 70196 265240
rect 119876 265296 121519 265298
rect 119876 265240 121458 265296
rect 121514 265240 121519 265296
rect 119876 265238 121519 265240
rect 67725 265235 67791 265238
rect 121453 265235 121519 265238
rect 67725 264618 67791 264621
rect 67725 264616 70196 264618
rect 67725 264560 67730 264616
rect 67786 264560 70196 264616
rect 67725 264558 70196 264560
rect 67725 264555 67791 264558
rect 119846 264074 119906 264588
rect 119846 264014 122850 264074
rect 67633 263938 67699 263941
rect 121545 263938 121611 263941
rect 67633 263936 70196 263938
rect 67633 263880 67638 263936
rect 67694 263880 70196 263936
rect 67633 263878 70196 263880
rect 119876 263936 121611 263938
rect 119876 263880 121550 263936
rect 121606 263880 121611 263936
rect 119876 263878 121611 263880
rect 67633 263875 67699 263878
rect 121545 263875 121611 263878
rect 122790 263666 122850 264014
rect 295609 263938 295675 263941
rect 292836 263936 295675 263938
rect 292836 263880 295614 263936
rect 295670 263880 295675 263936
rect 292836 263878 295675 263880
rect 295609 263875 295675 263878
rect 179462 263810 180044 263870
rect 176377 263802 176443 263805
rect 179462 263802 179522 263810
rect 176377 263800 179522 263802
rect 176377 263744 176382 263800
rect 176438 263744 179522 263800
rect 176377 263742 179522 263744
rect 176377 263739 176443 263742
rect 153694 263666 153700 263668
rect 122790 263606 153700 263666
rect 153694 263604 153700 263606
rect 153764 263604 153770 263668
rect 67725 263258 67791 263261
rect 121453 263258 121519 263261
rect 67725 263256 70196 263258
rect 67725 263200 67730 263256
rect 67786 263200 70196 263256
rect 67725 263198 70196 263200
rect 119876 263256 121519 263258
rect 119876 263200 121458 263256
rect 121514 263200 121519 263256
rect 119876 263198 121519 263200
rect 67725 263195 67791 263198
rect 121453 263195 121519 263198
rect 67633 262578 67699 262581
rect 121453 262578 121519 262581
rect 67633 262576 70196 262578
rect 67633 262520 67638 262576
rect 67694 262520 70196 262576
rect 67633 262518 70196 262520
rect 119876 262576 121519 262578
rect 119876 262520 121458 262576
rect 121514 262520 121519 262576
rect 119876 262518 121519 262520
rect 67633 262515 67699 262518
rect 121453 262515 121519 262518
rect 67265 261898 67331 261901
rect 121637 261898 121703 261901
rect 67265 261896 70196 261898
rect 67265 261840 67270 261896
rect 67326 261840 70196 261896
rect 67265 261838 70196 261840
rect 119876 261896 121703 261898
rect 119876 261840 121642 261896
rect 121698 261840 121703 261896
rect 119876 261838 121703 261840
rect 67265 261835 67331 261838
rect 121637 261835 121703 261838
rect 176653 261898 176719 261901
rect 176653 261896 179522 261898
rect 176653 261840 176658 261896
rect 176714 261840 179522 261896
rect 176653 261838 179522 261840
rect 176653 261835 176719 261838
rect 179462 261830 179522 261838
rect 179462 261770 180044 261830
rect 68369 261218 68435 261221
rect 121545 261218 121611 261221
rect 295609 261218 295675 261221
rect 68369 261216 70196 261218
rect 68369 261160 68374 261216
rect 68430 261160 70196 261216
rect 68369 261158 70196 261160
rect 119876 261216 121611 261218
rect 119876 261160 121550 261216
rect 121606 261160 121611 261216
rect 119876 261158 121611 261160
rect 292836 261216 295675 261218
rect 292836 261160 295614 261216
rect 295670 261160 295675 261216
rect 292836 261158 295675 261160
rect 68369 261155 68435 261158
rect 121545 261155 121611 261158
rect 295609 261155 295675 261158
rect 67633 260538 67699 260541
rect 121453 260538 121519 260541
rect 67633 260536 70196 260538
rect 67633 260480 67638 260536
rect 67694 260480 70196 260536
rect 67633 260478 70196 260480
rect 119876 260536 121519 260538
rect 119876 260480 121458 260536
rect 121514 260480 121519 260536
rect 119876 260478 121519 260480
rect 67633 260475 67699 260478
rect 121453 260475 121519 260478
rect 68093 259858 68159 259861
rect 121453 259858 121519 259861
rect 68093 259856 70196 259858
rect 68093 259800 68098 259856
rect 68154 259800 70196 259856
rect 68093 259798 70196 259800
rect 119876 259856 121519 259858
rect 119876 259800 121458 259856
rect 121514 259800 121519 259856
rect 119876 259798 121519 259800
rect 68093 259795 68159 259798
rect 121453 259795 121519 259798
rect 179462 259730 180044 259790
rect 176653 259722 176719 259725
rect 179462 259722 179522 259730
rect 176653 259720 179522 259722
rect 176653 259664 176658 259720
rect 176714 259664 179522 259720
rect 176653 259662 179522 259664
rect 176653 259659 176719 259662
rect 67725 259178 67791 259181
rect 121453 259178 121519 259181
rect 293217 259178 293283 259181
rect 67725 259176 70196 259178
rect 67725 259120 67730 259176
rect 67786 259120 70196 259176
rect 67725 259118 70196 259120
rect 119876 259176 121519 259178
rect 119876 259120 121458 259176
rect 121514 259120 121519 259176
rect 119876 259118 121519 259120
rect 292836 259176 293283 259178
rect 292836 259120 293222 259176
rect 293278 259120 293283 259176
rect 292836 259118 293283 259120
rect 67725 259115 67791 259118
rect 121453 259115 121519 259118
rect 293217 259115 293283 259118
rect 579613 258906 579679 258909
rect 583520 258906 584960 258996
rect 579613 258904 584960 258906
rect 579613 258848 579618 258904
rect 579674 258848 584960 258904
rect 579613 258846 584960 258848
rect 579613 258843 579679 258846
rect 583520 258756 584960 258846
rect 67633 258498 67699 258501
rect 67633 258496 70196 258498
rect 67633 258440 67638 258496
rect 67694 258440 70196 258496
rect 67633 258438 70196 258440
rect 67633 258435 67699 258438
rect 119846 257954 119906 258468
rect 157926 258028 157932 258092
rect 157996 258028 158002 258092
rect 157934 257954 157994 258028
rect 119846 257894 157994 257954
rect 69013 257818 69079 257821
rect 121545 257818 121611 257821
rect 69013 257816 70196 257818
rect 69013 257760 69018 257816
rect 69074 257760 70196 257816
rect 69013 257758 70196 257760
rect 119876 257816 121611 257818
rect 119876 257760 121550 257816
rect 121606 257760 121611 257816
rect 119876 257758 121611 257760
rect 69013 257755 69079 257758
rect 121545 257755 121611 257758
rect 64454 257212 64460 257276
rect 64524 257274 64530 257276
rect 68277 257274 68343 257277
rect 64524 257272 68343 257274
rect 64524 257216 68282 257272
rect 68338 257216 68343 257272
rect 64524 257214 68343 257216
rect 64524 257212 64530 257214
rect 68277 257211 68343 257214
rect 67633 257138 67699 257141
rect 121453 257138 121519 257141
rect 295701 257138 295767 257141
rect 67633 257136 70196 257138
rect 67633 257080 67638 257136
rect 67694 257080 70196 257136
rect 67633 257078 70196 257080
rect 119876 257136 121519 257138
rect 119876 257080 121458 257136
rect 121514 257080 121519 257136
rect 119876 257078 121519 257080
rect 292836 257136 295767 257138
rect 292836 257080 295706 257136
rect 295762 257080 295767 257136
rect 292836 257078 295767 257080
rect 67633 257075 67699 257078
rect 121453 257075 121519 257078
rect 295701 257075 295767 257078
rect 179462 257010 180044 257070
rect 179462 257005 179522 257010
rect 120574 256940 120580 257004
rect 120644 257002 120650 257004
rect 179413 257002 179522 257005
rect 120644 257000 179522 257002
rect 120644 256944 179418 257000
rect 179474 256944 179522 257000
rect 120644 256942 179522 256944
rect 120644 256940 120650 256942
rect 179413 256939 179479 256942
rect 67633 256458 67699 256461
rect 67633 256456 70196 256458
rect 67633 256400 67638 256456
rect 67694 256400 70196 256456
rect 67633 256398 70196 256400
rect 67633 256395 67699 256398
rect 119846 255914 119906 256428
rect 120993 255914 121059 255917
rect 119846 255912 121059 255914
rect 119846 255856 120998 255912
rect 121054 255856 121059 255912
rect 119846 255854 121059 255856
rect 120993 255851 121059 255854
rect 68829 255778 68895 255781
rect 68829 255776 70196 255778
rect 68829 255720 68834 255776
rect 68890 255720 70196 255776
rect 68829 255718 70196 255720
rect 68829 255715 68895 255718
rect 119846 255506 119906 255748
rect 160686 255506 160692 255508
rect 119846 255446 160692 255506
rect 160686 255444 160692 255446
rect 160756 255444 160762 255508
rect 120993 255370 121059 255373
rect 178534 255370 178540 255372
rect 120993 255368 178540 255370
rect 120993 255312 120998 255368
rect 121054 255312 178540 255368
rect 120993 255310 178540 255312
rect 120993 255307 121059 255310
rect 178534 255308 178540 255310
rect 178604 255308 178610 255372
rect 67725 255098 67791 255101
rect 122097 255098 122163 255101
rect 295701 255098 295767 255101
rect 67725 255096 70196 255098
rect 67725 255040 67730 255096
rect 67786 255040 70196 255096
rect 67725 255038 70196 255040
rect 119876 255096 122163 255098
rect 119876 255040 122102 255096
rect 122158 255040 122163 255096
rect 119876 255038 122163 255040
rect 292836 255096 295767 255098
rect 292836 255040 295706 255096
rect 295762 255040 295767 255096
rect 292836 255038 295767 255040
rect 67725 255035 67791 255038
rect 122097 255035 122163 255038
rect 295701 255035 295767 255038
rect 179830 254970 180044 255030
rect 176837 254962 176903 254965
rect 179321 254962 179387 254965
rect 179830 254962 179890 254970
rect 176837 254960 179890 254962
rect 176837 254904 176842 254960
rect 176898 254904 179326 254960
rect 179382 254904 179890 254960
rect 176837 254902 179890 254904
rect 176837 254899 176903 254902
rect 179321 254899 179387 254902
rect 67633 254418 67699 254421
rect 121453 254418 121519 254421
rect 67633 254416 70196 254418
rect 67633 254360 67638 254416
rect 67694 254360 70196 254416
rect 67633 254358 70196 254360
rect 119876 254416 121519 254418
rect 119876 254360 121458 254416
rect 121514 254360 121519 254416
rect 119876 254358 121519 254360
rect 67633 254355 67699 254358
rect 121453 254355 121519 254358
rect -960 254146 480 254236
rect 2773 254146 2839 254149
rect -960 254144 2839 254146
rect -960 254088 2778 254144
rect 2834 254088 2839 254144
rect -960 254086 2839 254088
rect -960 253996 480 254086
rect 2773 254083 2839 254086
rect 119286 254084 119292 254148
rect 119356 254146 119362 254148
rect 176837 254146 176903 254149
rect 119356 254144 176903 254146
rect 119356 254088 176842 254144
rect 176898 254088 176903 254144
rect 119356 254086 176903 254088
rect 119356 254084 119362 254086
rect 176837 254083 176903 254086
rect 67633 253738 67699 253741
rect 121545 253738 121611 253741
rect 67633 253736 70196 253738
rect 67633 253680 67638 253736
rect 67694 253680 70196 253736
rect 67633 253678 70196 253680
rect 119876 253736 121611 253738
rect 119876 253680 121550 253736
rect 121606 253680 121611 253736
rect 119876 253678 121611 253680
rect 67633 253675 67699 253678
rect 121545 253675 121611 253678
rect 67633 253058 67699 253061
rect 121453 253058 121519 253061
rect 67633 253056 70196 253058
rect 67633 253000 67638 253056
rect 67694 253000 70196 253056
rect 67633 252998 70196 253000
rect 119876 253056 121519 253058
rect 119876 253000 121458 253056
rect 121514 253000 121519 253056
rect 119876 252998 121519 253000
rect 67633 252995 67699 252998
rect 121453 252995 121519 252998
rect 179462 252930 180044 252990
rect 179462 252925 179522 252930
rect 179413 252920 179522 252925
rect 179413 252864 179418 252920
rect 179474 252864 179522 252920
rect 179413 252862 179522 252864
rect 179413 252859 179479 252862
rect 67633 252378 67699 252381
rect 296437 252378 296503 252381
rect 67633 252376 70196 252378
rect 67633 252320 67638 252376
rect 67694 252320 70196 252376
rect 292836 252376 296503 252378
rect 67633 252318 70196 252320
rect 67633 252315 67699 252318
rect 119846 251834 119906 252348
rect 292836 252320 296442 252376
rect 296498 252320 296503 252376
rect 292836 252318 296503 252320
rect 296437 252315 296503 252318
rect 119846 251774 122850 251834
rect 67541 251698 67607 251701
rect 121453 251698 121519 251701
rect 67541 251696 70196 251698
rect 67541 251640 67546 251696
rect 67602 251640 70196 251696
rect 67541 251638 70196 251640
rect 119876 251696 121519 251698
rect 119876 251640 121458 251696
rect 121514 251640 121519 251696
rect 119876 251638 121519 251640
rect 67541 251635 67607 251638
rect 121453 251635 121519 251638
rect 122790 251290 122850 251774
rect 161974 251290 161980 251292
rect 122790 251230 161980 251290
rect 161974 251228 161980 251230
rect 162044 251228 162050 251292
rect 68737 251018 68803 251021
rect 120165 251018 120231 251021
rect 120625 251018 120691 251021
rect 68737 251016 70196 251018
rect 68737 250960 68742 251016
rect 68798 250960 70196 251016
rect 68737 250958 70196 250960
rect 119876 251016 120691 251018
rect 119876 250960 120170 251016
rect 120226 250960 120630 251016
rect 120686 250960 120691 251016
rect 119876 250958 120691 250960
rect 68737 250955 68803 250958
rect 120165 250955 120231 250958
rect 120625 250955 120691 250958
rect 179462 250890 180044 250950
rect 176653 250882 176719 250885
rect 179462 250882 179522 250890
rect 176653 250880 179522 250882
rect 176653 250824 176658 250880
rect 176714 250824 179522 250880
rect 176653 250822 179522 250824
rect 176653 250819 176719 250822
rect 67633 250338 67699 250341
rect 121453 250338 121519 250341
rect 295793 250338 295859 250341
rect 67633 250336 70196 250338
rect 67633 250280 67638 250336
rect 67694 250280 70196 250336
rect 67633 250278 70196 250280
rect 119876 250336 121519 250338
rect 119876 250280 121458 250336
rect 121514 250280 121519 250336
rect 119876 250278 121519 250280
rect 292836 250336 295859 250338
rect 292836 250280 295798 250336
rect 295854 250280 295859 250336
rect 292836 250278 295859 250280
rect 67633 250275 67699 250278
rect 121453 250275 121519 250278
rect 295793 250275 295859 250278
rect 121545 249658 121611 249661
rect 119876 249656 121611 249658
rect 70166 249114 70226 249628
rect 119876 249600 121550 249656
rect 121606 249600 121611 249656
rect 119876 249598 121611 249600
rect 121545 249595 121611 249598
rect 64830 249054 70226 249114
rect 61878 248508 61884 248572
rect 61948 248570 61954 248572
rect 64830 248570 64890 249054
rect 67817 248978 67883 248981
rect 121453 248978 121519 248981
rect 67817 248976 70196 248978
rect 67817 248920 67822 248976
rect 67878 248920 70196 248976
rect 67817 248918 70196 248920
rect 119876 248976 121519 248978
rect 119876 248920 121458 248976
rect 121514 248920 121519 248976
rect 119876 248918 121519 248920
rect 67817 248915 67883 248918
rect 121453 248915 121519 248918
rect 61948 248510 64890 248570
rect 61948 248508 61954 248510
rect 67725 248298 67791 248301
rect 121453 248298 121519 248301
rect 296621 248298 296687 248301
rect 67725 248296 70196 248298
rect 67725 248240 67730 248296
rect 67786 248240 70196 248296
rect 67725 248238 70196 248240
rect 119876 248296 121519 248298
rect 119876 248240 121458 248296
rect 121514 248240 121519 248296
rect 119876 248238 121519 248240
rect 292836 248296 296687 248298
rect 292836 248240 296626 248296
rect 296682 248240 296687 248296
rect 292836 248238 296687 248240
rect 67725 248235 67791 248238
rect 121453 248235 121519 248238
rect 296621 248235 296687 248238
rect 179462 248170 180044 248230
rect 179229 248162 179295 248165
rect 179462 248162 179522 248170
rect 179229 248160 179522 248162
rect 179229 248104 179234 248160
rect 179290 248104 179522 248160
rect 179229 248102 179522 248104
rect 179229 248099 179295 248102
rect 120022 248026 120028 248028
rect 119846 247966 120028 248026
rect 67633 247618 67699 247621
rect 67633 247616 70196 247618
rect 67633 247560 67638 247616
rect 67694 247560 70196 247616
rect 119846 247588 119906 247966
rect 120022 247964 120028 247966
rect 120092 248026 120098 248028
rect 121545 248026 121611 248029
rect 120092 248024 121611 248026
rect 120092 247968 121550 248024
rect 121606 247968 121611 248024
rect 120092 247966 121611 247968
rect 120092 247964 120098 247966
rect 121545 247963 121611 247966
rect 67633 247558 70196 247560
rect 67633 247555 67699 247558
rect 299657 247076 299723 247077
rect 299606 247074 299612 247076
rect 299566 247014 299612 247074
rect 299676 247072 299723 247076
rect 299718 247016 299723 247072
rect 299606 247012 299612 247014
rect 299676 247012 299723 247016
rect 299657 247011 299723 247012
rect 121545 246938 121611 246941
rect 119876 246936 121611 246938
rect 70166 246394 70226 246908
rect 119876 246880 121550 246936
rect 121606 246880 121611 246936
rect 119876 246878 121611 246880
rect 121545 246875 121611 246878
rect 64830 246334 70226 246394
rect 63350 245788 63356 245852
rect 63420 245850 63426 245852
rect 64830 245850 64890 246334
rect 68645 246258 68711 246261
rect 121453 246258 121519 246261
rect 296897 246258 296963 246261
rect 68645 246256 70196 246258
rect 68645 246200 68650 246256
rect 68706 246200 70196 246256
rect 68645 246198 70196 246200
rect 119876 246256 121519 246258
rect 119876 246200 121458 246256
rect 121514 246200 121519 246256
rect 119876 246198 121519 246200
rect 292836 246256 296963 246258
rect 292836 246200 296902 246256
rect 296958 246200 296963 246256
rect 292836 246198 296963 246200
rect 68645 246195 68711 246198
rect 121453 246195 121519 246198
rect 296897 246195 296963 246198
rect 179830 246130 180044 246190
rect 120942 245924 120948 245988
rect 121012 245986 121018 245988
rect 179137 245986 179203 245989
rect 179830 245986 179890 246130
rect 121012 245984 179890 245986
rect 121012 245928 179142 245984
rect 179198 245928 179890 245984
rect 121012 245926 179890 245928
rect 121012 245924 121018 245926
rect 179137 245923 179203 245926
rect 63420 245790 64890 245850
rect 63420 245788 63426 245790
rect 67633 245578 67699 245581
rect 121545 245578 121611 245581
rect 67633 245576 70196 245578
rect 67633 245520 67638 245576
rect 67694 245520 70196 245576
rect 67633 245518 70196 245520
rect 119876 245576 121611 245578
rect 119876 245520 121550 245576
rect 121606 245520 121611 245576
rect 119876 245518 121611 245520
rect 67633 245515 67699 245518
rect 121545 245515 121611 245518
rect 579889 245578 579955 245581
rect 583520 245578 584960 245668
rect 579889 245576 584960 245578
rect 579889 245520 579894 245576
rect 579950 245520 584960 245576
rect 579889 245518 584960 245520
rect 579889 245515 579955 245518
rect 583520 245428 584960 245518
rect 69105 244898 69171 244901
rect 121453 244898 121519 244901
rect 69105 244896 70196 244898
rect 69105 244840 69110 244896
rect 69166 244840 70196 244896
rect 69105 244838 70196 244840
rect 119876 244896 121519 244898
rect 119876 244840 121458 244896
rect 121514 244840 121519 244896
rect 119876 244838 121519 244840
rect 69105 244835 69171 244838
rect 121453 244835 121519 244838
rect 68921 244218 68987 244221
rect 121545 244218 121611 244221
rect 68921 244216 70196 244218
rect 68921 244160 68926 244216
rect 68982 244160 70196 244216
rect 68921 244158 70196 244160
rect 119876 244216 121611 244218
rect 119876 244160 121550 244216
rect 121606 244160 121611 244216
rect 119876 244158 121611 244160
rect 68921 244155 68987 244158
rect 121545 244155 121611 244158
rect 179462 244090 180044 244150
rect 179321 244082 179387 244085
rect 179462 244082 179522 244090
rect 179321 244080 179522 244082
rect 179321 244024 179326 244080
rect 179382 244024 179522 244080
rect 179321 244022 179522 244024
rect 179321 244019 179387 244022
rect 69197 243538 69263 243541
rect 121453 243538 121519 243541
rect 295333 243538 295399 243541
rect 69197 243536 70196 243538
rect 69197 243480 69202 243536
rect 69258 243480 70196 243536
rect 69197 243478 70196 243480
rect 119876 243536 121519 243538
rect 119876 243480 121458 243536
rect 121514 243480 121519 243536
rect 119876 243478 121519 243480
rect 292836 243536 295399 243538
rect 292836 243480 295338 243536
rect 295394 243480 295399 243536
rect 292836 243478 295399 243480
rect 69197 243475 69263 243478
rect 121453 243475 121519 243478
rect 295333 243475 295399 243478
rect 179505 242994 179571 242997
rect 179822 242994 179828 242996
rect 179505 242992 179828 242994
rect 179505 242936 179510 242992
rect 179566 242936 179828 242992
rect 179505 242934 179828 242936
rect 179505 242931 179571 242934
rect 179822 242932 179828 242934
rect 179892 242932 179898 242996
rect 121453 242858 121519 242861
rect 119876 242856 121519 242858
rect 70166 242314 70226 242828
rect 119876 242800 121458 242856
rect 121514 242800 121519 242856
rect 119876 242798 121519 242800
rect 121453 242795 121519 242798
rect 119797 242586 119863 242589
rect 120942 242586 120948 242588
rect 119797 242584 120948 242586
rect 119797 242528 119802 242584
rect 119858 242528 120948 242584
rect 119797 242526 120948 242528
rect 119797 242523 119863 242526
rect 120942 242524 120948 242526
rect 121012 242524 121018 242588
rect 64830 242254 70226 242314
rect 63166 241708 63172 241772
rect 63236 241770 63242 241772
rect 64830 241770 64890 242254
rect 67725 242178 67791 242181
rect 121545 242178 121611 242181
rect 67725 242176 70196 242178
rect 67725 242120 67730 242176
rect 67786 242120 70196 242176
rect 67725 242118 70196 242120
rect 119876 242176 121611 242178
rect 119876 242120 121550 242176
rect 121606 242120 121611 242176
rect 119876 242118 121611 242120
rect 67725 242115 67791 242118
rect 121545 242115 121611 242118
rect 176837 242178 176903 242181
rect 176837 242176 179522 242178
rect 176837 242120 176842 242176
rect 176898 242120 179522 242176
rect 176837 242118 179522 242120
rect 176837 242115 176903 242118
rect 179462 242110 179522 242118
rect 179462 242050 180044 242110
rect 293309 241906 293375 241909
rect 299749 241906 299815 241909
rect 293309 241904 299815 241906
rect 293309 241848 293314 241904
rect 293370 241848 299754 241904
rect 299810 241848 299815 241904
rect 293309 241846 299815 241848
rect 293309 241843 293375 241846
rect 299749 241843 299815 241846
rect 63236 241710 64890 241770
rect 63236 241708 63242 241710
rect 67633 241498 67699 241501
rect 120073 241498 120139 241501
rect 295333 241498 295399 241501
rect 67633 241496 70196 241498
rect 67633 241440 67638 241496
rect 67694 241440 70196 241496
rect 67633 241438 70196 241440
rect 119876 241496 120139 241498
rect 119876 241440 120078 241496
rect 120134 241440 120139 241496
rect 119876 241438 120139 241440
rect 292836 241496 295399 241498
rect 292836 241440 295338 241496
rect 295394 241440 295399 241496
rect 292836 241438 295399 241440
rect 67633 241435 67699 241438
rect 120073 241435 120139 241438
rect 295333 241435 295399 241438
rect 144361 241226 144427 241229
rect 300945 241226 301011 241229
rect 144361 241224 301011 241226
rect -960 241090 480 241180
rect 144361 241168 144366 241224
rect 144422 241168 300950 241224
rect 301006 241168 301011 241224
rect 144361 241166 301011 241168
rect 144361 241163 144427 241166
rect 300945 241163 301011 241166
rect 3325 241090 3391 241093
rect -960 241088 3391 241090
rect -960 241032 3330 241088
rect 3386 241032 3391 241088
rect -960 241030 3391 241032
rect -960 240940 480 241030
rect 3325 241027 3391 241030
rect 291694 241028 291700 241092
rect 291764 241090 291770 241092
rect 293309 241090 293375 241093
rect 291764 241088 293375 241090
rect 291764 241032 293314 241088
rect 293370 241032 293375 241088
rect 291764 241030 293375 241032
rect 291764 241028 291770 241030
rect 293309 241027 293375 241030
rect 69841 240818 69907 240821
rect 121453 240818 121519 240821
rect 69841 240816 70196 240818
rect 69841 240760 69846 240816
rect 69902 240760 70196 240816
rect 69841 240758 70196 240760
rect 119876 240816 121519 240818
rect 119876 240760 121458 240816
rect 121514 240760 121519 240816
rect 119876 240758 121519 240760
rect 69841 240755 69907 240758
rect 121453 240755 121519 240758
rect 154021 240818 154087 240821
rect 154021 240816 176670 240818
rect 154021 240760 154026 240816
rect 154082 240760 176670 240816
rect 154021 240758 176670 240760
rect 154021 240755 154087 240758
rect 176610 240682 176670 240758
rect 188337 240682 188403 240685
rect 176610 240680 188403 240682
rect 176610 240624 188342 240680
rect 188398 240624 188403 240680
rect 176610 240622 188403 240624
rect 188337 240619 188403 240622
rect 121545 240138 121611 240141
rect 119876 240136 121611 240138
rect 119876 240080 121550 240136
rect 121606 240080 121611 240136
rect 119876 240078 121611 240080
rect 121545 240075 121611 240078
rect 117037 239866 117103 239869
rect 119102 239866 119108 239868
rect 117037 239864 119108 239866
rect 117037 239808 117042 239864
rect 117098 239808 119108 239864
rect 117037 239806 119108 239808
rect 117037 239803 117103 239806
rect 119102 239804 119108 239806
rect 119172 239804 119178 239868
rect 178534 238988 178540 239052
rect 178604 239050 178610 239052
rect 189993 239050 190059 239053
rect 178604 239048 190059 239050
rect 178604 238992 189998 239048
rect 190054 238992 190059 239048
rect 178604 238990 190059 238992
rect 178604 238988 178610 238990
rect 189993 238987 190059 238990
rect 161974 238852 161980 238916
rect 162044 238914 162050 238916
rect 273713 238914 273779 238917
rect 297357 238914 297423 238917
rect 162044 238912 297423 238914
rect 162044 238856 273718 238912
rect 273774 238856 297362 238912
rect 297418 238856 297423 238912
rect 162044 238854 297423 238856
rect 162044 238852 162050 238854
rect 273713 238851 273779 238854
rect 297357 238851 297423 238854
rect 82905 238778 82971 238781
rect 293902 238778 293908 238780
rect 82905 238776 293908 238778
rect 82905 238720 82910 238776
rect 82966 238720 293908 238776
rect 82905 238718 293908 238720
rect 82905 238715 82971 238718
rect 293902 238716 293908 238718
rect 293972 238716 293978 238780
rect 57830 238580 57836 238644
rect 57900 238642 57906 238644
rect 302325 238642 302391 238645
rect 57900 238640 302391 238642
rect 57900 238584 302330 238640
rect 302386 238584 302391 238640
rect 57900 238582 302391 238584
rect 57900 238580 57906 238582
rect 302325 238579 302391 238582
rect 171910 238444 171916 238508
rect 171980 238506 171986 238508
rect 204897 238506 204963 238509
rect 171980 238504 204963 238506
rect 171980 238448 204902 238504
rect 204958 238448 204963 238504
rect 171980 238446 204963 238448
rect 171980 238444 171986 238446
rect 204897 238443 204963 238446
rect 269757 238506 269823 238509
rect 299974 238506 299980 238508
rect 269757 238504 299980 238506
rect 269757 238448 269762 238504
rect 269818 238448 299980 238504
rect 269757 238446 299980 238448
rect 269757 238443 269823 238446
rect 299974 238444 299980 238446
rect 300044 238444 300050 238508
rect 105445 238098 105511 238101
rect 171726 238098 171732 238100
rect 105445 238096 171732 238098
rect 105445 238040 105450 238096
rect 105506 238040 171732 238096
rect 105445 238038 171732 238040
rect 105445 238035 105511 238038
rect 171726 238036 171732 238038
rect 171796 238036 171802 238100
rect 250805 238098 250871 238101
rect 265566 238098 265572 238100
rect 250805 238096 265572 238098
rect 250805 238040 250810 238096
rect 250866 238040 265572 238096
rect 250805 238038 265572 238040
rect 250805 238035 250871 238038
rect 265566 238036 265572 238038
rect 265636 238036 265642 238100
rect 122189 237962 122255 237965
rect 328494 237962 328500 237964
rect 122189 237960 328500 237962
rect 122189 237904 122194 237960
rect 122250 237904 328500 237960
rect 122189 237902 328500 237904
rect 122189 237899 122255 237902
rect 328494 237900 328500 237902
rect 328564 237900 328570 237964
rect 95693 237282 95759 237285
rect 96521 237282 96587 237285
rect 156454 237282 156460 237284
rect 95693 237280 156460 237282
rect 95693 237224 95698 237280
rect 95754 237224 96526 237280
rect 96582 237224 156460 237280
rect 95693 237222 156460 237224
rect 95693 237219 95759 237222
rect 96521 237219 96587 237222
rect 156454 237220 156460 237222
rect 156524 237220 156530 237284
rect 160686 237220 160692 237284
rect 160756 237282 160762 237284
rect 305177 237282 305243 237285
rect 160756 237280 305243 237282
rect 160756 237224 305182 237280
rect 305238 237224 305243 237280
rect 160756 237222 305243 237224
rect 160756 237220 160762 237222
rect 305177 237219 305243 237222
rect 106733 237146 106799 237149
rect 120574 237146 120580 237148
rect 106733 237144 120580 237146
rect 106733 237088 106738 237144
rect 106794 237088 120580 237144
rect 106733 237086 120580 237088
rect 106733 237083 106799 237086
rect 120574 237084 120580 237086
rect 120644 237084 120650 237148
rect 64454 236540 64460 236604
rect 64524 236602 64530 236604
rect 117957 236602 118023 236605
rect 64524 236600 118023 236602
rect 64524 236544 117962 236600
rect 118018 236544 118023 236600
rect 64524 236542 118023 236544
rect 64524 236540 64530 236542
rect 117957 236539 118023 236542
rect 61878 235860 61884 235924
rect 61948 235922 61954 235924
rect 138013 235922 138079 235925
rect 295374 235922 295380 235924
rect 61948 235920 295380 235922
rect 61948 235864 138018 235920
rect 138074 235864 295380 235920
rect 61948 235862 295380 235864
rect 61948 235860 61954 235862
rect 138013 235859 138079 235862
rect 295374 235860 295380 235862
rect 295444 235860 295450 235924
rect 68737 233882 68803 233885
rect 322054 233882 322060 233884
rect 68737 233880 322060 233882
rect 68737 233824 68742 233880
rect 68798 233824 322060 233880
rect 68737 233822 322060 233824
rect 68737 233819 68803 233822
rect 322054 233820 322060 233822
rect 322124 233820 322130 233884
rect 63166 233140 63172 233204
rect 63236 233202 63242 233204
rect 264973 233202 265039 233205
rect 63236 233200 265039 233202
rect 63236 233144 264978 233200
rect 265034 233144 265039 233200
rect 63236 233142 265039 233144
rect 63236 233140 63242 233142
rect 264973 233139 265039 233142
rect 579613 232386 579679 232389
rect 583520 232386 584960 232476
rect 579613 232384 584960 232386
rect 579613 232328 579618 232384
rect 579674 232328 584960 232384
rect 579613 232326 584960 232328
rect 579613 232323 579679 232326
rect 583520 232236 584960 232326
rect 59118 231780 59124 231844
rect 59188 231842 59194 231844
rect 287053 231842 287119 231845
rect 59188 231840 287119 231842
rect 59188 231784 287058 231840
rect 287114 231784 287119 231840
rect 59188 231782 287119 231784
rect 59188 231780 59194 231782
rect 287053 231779 287119 231782
rect 153694 231644 153700 231708
rect 153764 231706 153770 231708
rect 269757 231706 269823 231709
rect 153764 231704 269823 231706
rect 153764 231648 269762 231704
rect 269818 231648 269823 231704
rect 153764 231646 269823 231648
rect 153764 231644 153770 231646
rect 269757 231643 269823 231646
rect 63350 230420 63356 230484
rect 63420 230482 63426 230484
rect 299606 230482 299612 230484
rect 63420 230422 299612 230482
rect 63420 230420 63426 230422
rect 299606 230420 299612 230422
rect 299676 230420 299682 230484
rect 269614 229740 269620 229804
rect 269684 229802 269690 229804
rect 313273 229802 313339 229805
rect 269684 229800 313339 229802
rect 269684 229744 313278 229800
rect 313334 229744 313339 229800
rect 269684 229742 313339 229744
rect 269684 229740 269690 229742
rect 313273 229739 313339 229742
rect 271086 228244 271092 228308
rect 271156 228306 271162 228308
rect 298093 228306 298159 228309
rect 271156 228304 298159 228306
rect 271156 228248 298098 228304
rect 298154 228248 298159 228304
rect 271156 228246 298159 228248
rect 271156 228244 271162 228246
rect 298093 228243 298159 228246
rect -960 227884 480 228124
rect 157926 227564 157932 227628
rect 157996 227626 158002 227628
rect 276657 227626 276723 227629
rect 157996 227624 276723 227626
rect 157996 227568 276662 227624
rect 276718 227568 276723 227624
rect 157996 227566 276723 227568
rect 157996 227564 158002 227566
rect 276657 227563 276723 227566
rect 273846 226884 273852 226948
rect 273916 226946 273922 226948
rect 291694 226946 291700 226948
rect 273916 226886 291700 226946
rect 273916 226884 273922 226886
rect 291694 226884 291700 226886
rect 291764 226884 291770 226948
rect 64597 225586 64663 225589
rect 251214 225586 251220 225588
rect 64597 225584 251220 225586
rect 64597 225528 64602 225584
rect 64658 225528 251220 225584
rect 64597 225526 251220 225528
rect 64597 225523 64663 225526
rect 251214 225524 251220 225526
rect 251284 225524 251290 225588
rect 163589 221506 163655 221509
rect 336958 221506 336964 221508
rect 163589 221504 336964 221506
rect 163589 221448 163594 221504
rect 163650 221448 336964 221504
rect 163589 221446 336964 221448
rect 163589 221443 163655 221446
rect 336958 221444 336964 221446
rect 337028 221444 337034 221508
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect 77293 215930 77359 215933
rect 260966 215930 260972 215932
rect 77293 215928 260972 215930
rect 77293 215872 77298 215928
rect 77354 215872 260972 215928
rect 77293 215870 260972 215872
rect 77293 215867 77359 215870
rect 260966 215868 260972 215870
rect 261036 215868 261042 215932
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 68829 214570 68895 214573
rect 327206 214570 327212 214572
rect 68829 214568 327212 214570
rect 68829 214512 68834 214568
rect 68890 214512 327212 214568
rect 68829 214510 327212 214512
rect 68829 214507 68895 214510
rect 327206 214508 327212 214510
rect 327276 214508 327282 214572
rect 54937 213210 55003 213213
rect 265014 213210 265020 213212
rect 54937 213208 265020 213210
rect 54937 213152 54942 213208
rect 54998 213152 265020 213208
rect 54937 213150 265020 213152
rect 54937 213147 55003 213150
rect 265014 213148 265020 213150
rect 265084 213148 265090 213212
rect 166257 211986 166323 211989
rect 335854 211986 335860 211988
rect 166257 211984 335860 211986
rect 166257 211928 166262 211984
rect 166318 211928 335860 211984
rect 166257 211926 335860 211928
rect 166257 211923 166323 211926
rect 335854 211924 335860 211926
rect 335924 211924 335930 211988
rect 53557 211850 53623 211853
rect 335670 211850 335676 211852
rect 53557 211848 335676 211850
rect 53557 211792 53562 211848
rect 53618 211792 335676 211848
rect 53557 211790 335676 211792
rect 53557 211787 53623 211790
rect 335670 211788 335676 211790
rect 335740 211788 335746 211852
rect 242249 210626 242315 210629
rect 346342 210626 346348 210628
rect 242249 210624 346348 210626
rect 242249 210568 242254 210624
rect 242310 210568 346348 210624
rect 242249 210566 346348 210568
rect 242249 210563 242315 210566
rect 346342 210564 346348 210566
rect 346412 210564 346418 210628
rect 52361 210490 52427 210493
rect 269062 210490 269068 210492
rect 52361 210488 269068 210490
rect 52361 210432 52366 210488
rect 52422 210432 269068 210488
rect 52361 210430 269068 210432
rect 52361 210427 52427 210430
rect 269062 210428 269068 210430
rect 269132 210428 269138 210492
rect 84377 210354 84443 210357
rect 328678 210354 328684 210356
rect 84377 210352 328684 210354
rect 84377 210296 84382 210352
rect 84438 210296 328684 210352
rect 84377 210294 328684 210296
rect 84377 210291 84443 210294
rect 328678 210292 328684 210294
rect 328748 210292 328754 210356
rect 145741 206410 145807 206413
rect 263542 206410 263548 206412
rect 145741 206408 263548 206410
rect 145741 206352 145746 206408
rect 145802 206352 263548 206408
rect 145741 206350 263548 206352
rect 145741 206347 145807 206350
rect 263542 206348 263548 206350
rect 263612 206348 263618 206412
rect 110413 206274 110479 206277
rect 255262 206274 255268 206276
rect 110413 206272 255268 206274
rect 110413 206216 110418 206272
rect 110474 206216 255268 206272
rect 110413 206214 255268 206216
rect 110413 206211 110479 206214
rect 255262 206212 255268 206214
rect 255332 206212 255338 206276
rect 582373 205730 582439 205733
rect 583520 205730 584960 205820
rect 582373 205728 584960 205730
rect 582373 205672 582378 205728
rect 582434 205672 584960 205728
rect 582373 205670 584960 205672
rect 582373 205667 582439 205670
rect 583520 205580 584960 205670
rect 327717 204914 327783 204917
rect 331254 204914 331260 204916
rect 327717 204912 331260 204914
rect 327717 204856 327722 204912
rect 327778 204856 331260 204912
rect 327717 204854 331260 204856
rect 327717 204851 327783 204854
rect 331254 204852 331260 204854
rect 331324 204852 331330 204916
rect -960 201922 480 202012
rect 3601 201922 3667 201925
rect -960 201920 3667 201922
rect -960 201864 3606 201920
rect 3662 201864 3667 201920
rect -960 201862 3667 201864
rect -960 201772 480 201862
rect 3601 201859 3667 201862
rect 117957 200698 118023 200701
rect 340822 200698 340828 200700
rect 117957 200696 340828 200698
rect 117957 200640 117962 200696
rect 118018 200640 340828 200696
rect 117957 200638 340828 200640
rect 117957 200635 118023 200638
rect 340822 200636 340828 200638
rect 340892 200636 340898 200700
rect 134701 199338 134767 199341
rect 270534 199338 270540 199340
rect 134701 199336 270540 199338
rect 134701 199280 134706 199336
rect 134762 199280 270540 199336
rect 134701 199278 270540 199280
rect 134701 199275 134767 199278
rect 270534 199276 270540 199278
rect 270604 199276 270610 199340
rect 74533 197978 74599 197981
rect 327022 197978 327028 197980
rect 74533 197976 327028 197978
rect 74533 197920 74538 197976
rect 74594 197920 327028 197976
rect 74533 197918 327028 197920
rect 74533 197915 74599 197918
rect 327022 197916 327028 197918
rect 327092 197916 327098 197980
rect 158529 196618 158595 196621
rect 197997 196618 198063 196621
rect 158529 196616 198063 196618
rect 158529 196560 158534 196616
rect 158590 196560 198002 196616
rect 198058 196560 198063 196616
rect 158529 196558 198063 196560
rect 158529 196555 158595 196558
rect 197997 196555 198063 196558
rect 152958 193836 152964 193900
rect 153028 193898 153034 193900
rect 196617 193898 196683 193901
rect 153028 193896 196683 193898
rect 153028 193840 196622 193896
rect 196678 193840 196683 193896
rect 153028 193838 196683 193840
rect 153028 193836 153034 193838
rect 196617 193835 196683 193838
rect 154113 192674 154179 192677
rect 259678 192674 259684 192676
rect 154113 192672 259684 192674
rect 154113 192616 154118 192672
rect 154174 192616 259684 192672
rect 154113 192614 259684 192616
rect 154113 192611 154179 192614
rect 259678 192612 259684 192614
rect 259748 192612 259754 192676
rect 137369 192538 137435 192541
rect 329782 192538 329788 192540
rect 137369 192536 329788 192538
rect 137369 192480 137374 192536
rect 137430 192480 329788 192536
rect 137369 192478 329788 192480
rect 137369 192475 137435 192478
rect 329782 192476 329788 192478
rect 329852 192476 329858 192540
rect 580441 192538 580507 192541
rect 583520 192538 584960 192628
rect 580441 192536 584960 192538
rect 580441 192480 580446 192536
rect 580502 192480 584960 192536
rect 580441 192478 584960 192480
rect 580441 192475 580507 192478
rect 583520 192388 584960 192478
rect 57789 191042 57855 191045
rect 259494 191042 259500 191044
rect 57789 191040 259500 191042
rect 57789 190984 57794 191040
rect 57850 190984 259500 191040
rect 57789 190982 259500 190984
rect 57789 190979 57855 190982
rect 259494 190980 259500 190982
rect 259564 190980 259570 191044
rect 60641 189682 60707 189685
rect 260966 189682 260972 189684
rect 60641 189680 260972 189682
rect 60641 189624 60646 189680
rect 60702 189624 260972 189680
rect 60641 189622 260972 189624
rect 60641 189619 60707 189622
rect 260966 189620 260972 189622
rect 261036 189620 261042 189684
rect 306230 189620 306236 189684
rect 306300 189682 306306 189684
rect 317413 189682 317479 189685
rect 306300 189680 317479 189682
rect 306300 189624 317418 189680
rect 317474 189624 317479 189680
rect 306300 189622 317479 189624
rect 306300 189620 306306 189622
rect 317413 189619 317479 189622
rect -960 188866 480 188956
rect 3141 188866 3207 188869
rect -960 188864 3207 188866
rect -960 188808 3146 188864
rect 3202 188808 3207 188864
rect -960 188806 3207 188808
rect -960 188716 480 188806
rect 3141 188803 3207 188806
rect 100753 188322 100819 188325
rect 254526 188322 254532 188324
rect 100753 188320 254532 188322
rect 100753 188264 100758 188320
rect 100814 188264 254532 188320
rect 100753 188262 254532 188264
rect 100753 188259 100819 188262
rect 254526 188260 254532 188262
rect 254596 188260 254602 188324
rect 80053 186962 80119 186965
rect 320398 186962 320404 186964
rect 80053 186960 320404 186962
rect 80053 186904 80058 186960
rect 80114 186904 320404 186960
rect 80053 186902 320404 186904
rect 80053 186899 80119 186902
rect 320398 186900 320404 186902
rect 320468 186900 320474 186964
rect 232497 185602 232563 185605
rect 256918 185602 256924 185604
rect 232497 185600 256924 185602
rect 232497 185544 232502 185600
rect 232558 185544 256924 185600
rect 232497 185542 256924 185544
rect 232497 185539 232563 185542
rect 256918 185540 256924 185542
rect 256988 185540 256994 185604
rect 161381 184378 161447 184381
rect 192477 184378 192543 184381
rect 161381 184376 192543 184378
rect 161381 184320 161386 184376
rect 161442 184320 192482 184376
rect 192538 184320 192543 184376
rect 161381 184318 192543 184320
rect 161381 184315 161447 184318
rect 192477 184315 192543 184318
rect 214557 184378 214623 184381
rect 266302 184378 266308 184380
rect 214557 184376 266308 184378
rect 214557 184320 214562 184376
rect 214618 184320 266308 184376
rect 214557 184318 266308 184320
rect 214557 184315 214623 184318
rect 266302 184316 266308 184318
rect 266372 184316 266378 184380
rect 73153 184242 73219 184245
rect 323025 184242 323091 184245
rect 73153 184240 323091 184242
rect 73153 184184 73158 184240
rect 73214 184184 323030 184240
rect 323086 184184 323091 184240
rect 73153 184182 323091 184184
rect 73153 184179 73219 184182
rect 323025 184179 323091 184182
rect 98637 182882 98703 182885
rect 332726 182882 332732 182884
rect 98637 182880 332732 182882
rect 98637 182824 98642 182880
rect 98698 182824 332732 182880
rect 98637 182822 332732 182824
rect 98637 182819 98703 182822
rect 332726 182820 332732 182822
rect 332796 182820 332802 182884
rect 130469 181522 130535 181525
rect 255446 181522 255452 181524
rect 130469 181520 255452 181522
rect 130469 181464 130474 181520
rect 130530 181464 255452 181520
rect 130469 181462 255452 181464
rect 130469 181459 130535 181462
rect 255446 181460 255452 181462
rect 255516 181460 255522 181524
rect 75177 181386 75243 181389
rect 332685 181386 332751 181389
rect 75177 181384 332751 181386
rect 75177 181328 75182 181384
rect 75238 181328 332690 181384
rect 332746 181328 332751 181384
rect 75177 181326 332751 181328
rect 75177 181323 75243 181326
rect 332685 181323 332751 181326
rect 239489 180162 239555 180165
rect 256734 180162 256740 180164
rect 239489 180160 256740 180162
rect 239489 180104 239494 180160
rect 239550 180104 256740 180160
rect 239489 180102 256740 180104
rect 239489 180099 239555 180102
rect 256734 180100 256740 180102
rect 256804 180100 256810 180164
rect 53741 180026 53807 180029
rect 249006 180026 249012 180028
rect 53741 180024 249012 180026
rect 53741 179968 53746 180024
rect 53802 179968 249012 180024
rect 53741 179966 249012 179968
rect 53741 179963 53807 179966
rect 249006 179964 249012 179966
rect 249076 179964 249082 180028
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect 313917 178802 313983 178805
rect 334014 178802 334020 178804
rect 313917 178800 334020 178802
rect 313917 178744 313922 178800
rect 313978 178744 334020 178800
rect 313917 178742 334020 178744
rect 313917 178739 313983 178742
rect 334014 178740 334020 178742
rect 334084 178740 334090 178804
rect 55121 178666 55187 178669
rect 336917 178666 336983 178669
rect 55121 178664 336983 178666
rect 55121 178608 55126 178664
rect 55182 178608 336922 178664
rect 336978 178608 336983 178664
rect 55121 178606 336983 178608
rect 55121 178603 55187 178606
rect 336917 178603 336983 178606
rect 247769 177714 247835 177717
rect 249190 177714 249196 177716
rect 247769 177712 249196 177714
rect 247769 177656 247774 177712
rect 247830 177656 249196 177712
rect 247769 177654 249196 177656
rect 247769 177651 247835 177654
rect 249190 177652 249196 177654
rect 249260 177652 249266 177716
rect 99414 177516 99420 177580
rect 99484 177578 99490 177580
rect 100661 177578 100727 177581
rect 102041 177580 102107 177581
rect 101990 177578 101996 177580
rect 99484 177576 100727 177578
rect 99484 177520 100666 177576
rect 100722 177520 100727 177576
rect 99484 177518 100727 177520
rect 101950 177518 101996 177578
rect 102060 177576 102107 177580
rect 102102 177520 102107 177576
rect 99484 177516 99490 177518
rect 100661 177515 100727 177518
rect 101990 177516 101996 177518
rect 102060 177516 102107 177520
rect 106038 177516 106044 177580
rect 106108 177578 106114 177580
rect 106181 177578 106247 177581
rect 106108 177576 106247 177578
rect 106108 177520 106186 177576
rect 106242 177520 106247 177576
rect 106108 177518 106247 177520
rect 106108 177516 106114 177518
rect 102041 177515 102107 177516
rect 106181 177515 106247 177518
rect 106958 177516 106964 177580
rect 107028 177578 107034 177580
rect 107561 177578 107627 177581
rect 107028 177576 107627 177578
rect 107028 177520 107566 177576
rect 107622 177520 107627 177576
rect 107028 177518 107627 177520
rect 107028 177516 107034 177518
rect 107561 177515 107627 177518
rect 112110 177516 112116 177580
rect 112180 177578 112186 177580
rect 112989 177578 113055 177581
rect 112180 177576 113055 177578
rect 112180 177520 112994 177576
rect 113050 177520 113055 177576
rect 112180 177518 113055 177520
rect 112180 177516 112186 177518
rect 112989 177515 113055 177518
rect 114134 177516 114140 177580
rect 114204 177578 114210 177580
rect 114461 177578 114527 177581
rect 116945 177580 117011 177581
rect 116894 177578 116900 177580
rect 114204 177576 114527 177578
rect 114204 177520 114466 177576
rect 114522 177520 114527 177576
rect 114204 177518 114527 177520
rect 116854 177518 116900 177578
rect 116964 177576 117011 177580
rect 117006 177520 117011 177576
rect 114204 177516 114210 177518
rect 114461 177515 114527 177518
rect 116894 177516 116900 177518
rect 116964 177516 117011 177520
rect 118366 177516 118372 177580
rect 118436 177578 118442 177580
rect 118601 177578 118667 177581
rect 118436 177576 118667 177578
rect 118436 177520 118606 177576
rect 118662 177520 118667 177576
rect 118436 177518 118667 177520
rect 118436 177516 118442 177518
rect 116945 177515 117011 177516
rect 118601 177515 118667 177518
rect 127014 177516 127020 177580
rect 127084 177578 127090 177580
rect 127801 177578 127867 177581
rect 129457 177580 129523 177581
rect 129406 177578 129412 177580
rect 127084 177576 127867 177578
rect 127084 177520 127806 177576
rect 127862 177520 127867 177576
rect 127084 177518 127867 177520
rect 129366 177518 129412 177578
rect 129476 177576 129523 177580
rect 129518 177520 129523 177576
rect 127084 177516 127090 177518
rect 127801 177515 127867 177518
rect 129406 177516 129412 177518
rect 129476 177516 129523 177520
rect 133086 177516 133092 177580
rect 133156 177578 133162 177580
rect 133781 177578 133847 177581
rect 133156 177576 133847 177578
rect 133156 177520 133786 177576
rect 133842 177520 133847 177576
rect 133156 177518 133847 177520
rect 133156 177516 133162 177518
rect 129457 177515 129523 177516
rect 133781 177515 133847 177518
rect 311157 177442 311223 177445
rect 331438 177442 331444 177444
rect 311157 177440 331444 177442
rect 311157 177384 311162 177440
rect 311218 177384 331444 177440
rect 311157 177382 331444 177384
rect 311157 177379 311223 177382
rect 331438 177380 331444 177382
rect 331508 177380 331514 177444
rect 239397 177306 239463 177309
rect 257838 177306 257844 177308
rect 239397 177304 257844 177306
rect 239397 177248 239402 177304
rect 239458 177248 257844 177304
rect 239397 177246 257844 177248
rect 239397 177243 239463 177246
rect 257838 177244 257844 177246
rect 257908 177244 257914 177308
rect 315297 177306 315363 177309
rect 336774 177306 336780 177308
rect 315297 177304 336780 177306
rect 315297 177248 315302 177304
rect 315358 177248 336780 177304
rect 315297 177246 336780 177248
rect 315297 177243 315363 177246
rect 336774 177244 336780 177246
rect 336844 177244 336850 177308
rect 110689 177172 110755 177173
rect 110638 177170 110644 177172
rect 110598 177110 110644 177170
rect 110708 177168 110755 177172
rect 110750 177112 110755 177168
rect 110638 177108 110644 177110
rect 110708 177108 110755 177112
rect 113214 177108 113220 177172
rect 113284 177170 113290 177172
rect 113909 177170 113975 177173
rect 113284 177168 113975 177170
rect 113284 177112 113914 177168
rect 113970 177112 113975 177168
rect 113284 177110 113975 177112
rect 113284 177108 113290 177110
rect 110689 177107 110755 177108
rect 113909 177107 113975 177110
rect 103278 176972 103284 177036
rect 103348 177034 103354 177036
rect 169109 177034 169175 177037
rect 103348 177032 169175 177034
rect 103348 176976 169114 177032
rect 169170 176976 169175 177032
rect 103348 176974 169175 176976
rect 103348 176972 103354 176974
rect 169109 176971 169175 176974
rect 97022 176836 97028 176900
rect 97092 176898 97098 176900
rect 97809 176898 97875 176901
rect 97092 176896 97875 176898
rect 97092 176840 97814 176896
rect 97870 176840 97875 176896
rect 97092 176838 97875 176840
rect 97092 176836 97098 176838
rect 97809 176835 97875 176838
rect 100702 176836 100708 176900
rect 100772 176898 100778 176900
rect 166206 176898 166212 176900
rect 100772 176838 166212 176898
rect 100772 176836 100778 176838
rect 166206 176836 166212 176838
rect 166276 176836 166282 176900
rect 108113 176764 108179 176765
rect 108062 176762 108068 176764
rect 108022 176702 108068 176762
rect 108132 176760 108179 176764
rect 108174 176704 108179 176760
rect 108062 176700 108068 176702
rect 108132 176700 108179 176704
rect 109534 176700 109540 176764
rect 109604 176762 109610 176764
rect 109861 176762 109927 176765
rect 119705 176764 119771 176765
rect 119654 176762 119660 176764
rect 109604 176760 109927 176762
rect 109604 176704 109866 176760
rect 109922 176704 109927 176760
rect 109604 176702 109927 176704
rect 119614 176702 119660 176762
rect 119724 176760 119771 176764
rect 119766 176704 119771 176760
rect 109604 176700 109610 176702
rect 108113 176699 108179 176700
rect 109861 176699 109927 176702
rect 119654 176700 119660 176702
rect 119724 176700 119771 176704
rect 121862 176700 121868 176764
rect 121932 176762 121938 176764
rect 122005 176762 122071 176765
rect 123017 176764 123083 176765
rect 122966 176762 122972 176764
rect 121932 176760 122071 176762
rect 121932 176704 122010 176760
rect 122066 176704 122071 176760
rect 121932 176702 122071 176704
rect 122926 176702 122972 176762
rect 123036 176760 123083 176764
rect 123078 176704 123083 176760
rect 121932 176700 121938 176702
rect 119705 176699 119771 176700
rect 122005 176699 122071 176702
rect 122966 176700 122972 176702
rect 123036 176700 123083 176704
rect 124438 176700 124444 176764
rect 124508 176762 124514 176764
rect 124949 176762 125015 176765
rect 124508 176760 125015 176762
rect 124508 176704 124954 176760
rect 125010 176704 125015 176760
rect 124508 176702 125015 176704
rect 124508 176700 124514 176702
rect 123017 176699 123083 176700
rect 124949 176699 125015 176702
rect 125726 176700 125732 176764
rect 125796 176762 125802 176764
rect 125869 176762 125935 176765
rect 128261 176762 128327 176765
rect 132033 176764 132099 176765
rect 134425 176764 134491 176765
rect 135713 176764 135779 176765
rect 148225 176764 148291 176765
rect 131982 176762 131988 176764
rect 125796 176760 125935 176762
rect 125796 176704 125874 176760
rect 125930 176704 125935 176760
rect 125796 176702 125935 176704
rect 125796 176700 125802 176702
rect 125869 176699 125935 176702
rect 128126 176760 128327 176762
rect 128126 176704 128266 176760
rect 128322 176704 128327 176760
rect 128126 176702 128327 176704
rect 131942 176702 131988 176762
rect 132052 176760 132099 176764
rect 134374 176762 134380 176764
rect 132094 176704 132099 176760
rect 128126 176492 128186 176702
rect 128261 176699 128327 176702
rect 131982 176700 131988 176702
rect 132052 176700 132099 176704
rect 134334 176702 134380 176762
rect 134444 176760 134491 176764
rect 135662 176762 135668 176764
rect 134486 176704 134491 176760
rect 134374 176700 134380 176702
rect 134444 176700 134491 176704
rect 135622 176702 135668 176762
rect 135732 176760 135779 176764
rect 148174 176762 148180 176764
rect 135774 176704 135779 176760
rect 135662 176700 135668 176702
rect 135732 176700 135779 176704
rect 148134 176702 148180 176762
rect 148244 176760 148291 176764
rect 148286 176704 148291 176760
rect 148174 176700 148180 176702
rect 148244 176700 148291 176704
rect 158846 176700 158852 176764
rect 158916 176762 158922 176764
rect 158989 176762 159055 176765
rect 158916 176760 159055 176762
rect 158916 176704 158994 176760
rect 159050 176704 159055 176760
rect 158916 176702 159055 176704
rect 158916 176700 158922 176702
rect 132033 176699 132099 176700
rect 134425 176699 134491 176700
rect 135713 176699 135779 176700
rect 148225 176699 148291 176700
rect 158989 176699 159055 176702
rect 264094 176700 264100 176764
rect 264164 176762 264170 176764
rect 316033 176762 316099 176765
rect 320173 176764 320239 176765
rect 320173 176762 320220 176764
rect 264164 176760 316099 176762
rect 264164 176704 316038 176760
rect 316094 176704 316099 176760
rect 264164 176702 316099 176704
rect 320128 176760 320220 176762
rect 320128 176704 320178 176760
rect 320128 176702 320220 176704
rect 264164 176700 264170 176702
rect 316033 176699 316099 176702
rect 320173 176700 320220 176702
rect 320284 176700 320290 176764
rect 320817 176762 320883 176765
rect 321645 176762 321711 176765
rect 320817 176760 321711 176762
rect 320817 176704 320822 176760
rect 320878 176704 321650 176760
rect 321706 176704 321711 176760
rect 320817 176702 321711 176704
rect 320173 176699 320239 176700
rect 320817 176699 320883 176702
rect 321645 176699 321711 176702
rect 128118 176428 128124 176492
rect 128188 176428 128194 176492
rect 319437 176218 319503 176221
rect 321502 176218 321508 176220
rect 319437 176216 321508 176218
rect 319437 176160 319442 176216
rect 319498 176160 321508 176216
rect 319437 176158 321508 176160
rect 319437 176155 319503 176158
rect 321502 176156 321508 176158
rect 321572 176156 321578 176220
rect 244917 176082 244983 176085
rect 252502 176082 252508 176084
rect 244917 176080 252508 176082
rect -960 175796 480 176036
rect 244917 176024 244922 176080
rect 244978 176024 252508 176080
rect 244917 176022 252508 176024
rect 244917 176019 244983 176022
rect 252502 176020 252508 176022
rect 252572 176020 252578 176084
rect 155217 175946 155283 175949
rect 173893 175946 173959 175949
rect 155217 175944 173959 175946
rect 155217 175888 155222 175944
rect 155278 175888 173898 175944
rect 173954 175888 173959 175944
rect 155217 175886 173959 175888
rect 155217 175883 155283 175886
rect 173893 175883 173959 175886
rect 186957 175946 187023 175949
rect 338389 175946 338455 175949
rect 186957 175944 338455 175946
rect 186957 175888 186962 175944
rect 187018 175888 338394 175944
rect 338450 175888 338455 175944
rect 186957 175886 338455 175888
rect 186957 175883 187023 175886
rect 338389 175883 338455 175886
rect 248045 175810 248111 175813
rect 321461 175810 321527 175813
rect 248045 175808 248338 175810
rect 248045 175752 248050 175808
rect 248106 175752 248338 175808
rect 248045 175750 248338 175752
rect 248045 175747 248111 175750
rect 213913 175674 213979 175677
rect 213913 175672 217212 175674
rect 213913 175616 213918 175672
rect 213974 175616 217212 175672
rect 248278 175644 248338 175750
rect 321461 175808 321570 175810
rect 321461 175752 321466 175808
rect 321522 175752 321570 175808
rect 321461 175747 321570 175752
rect 307569 175674 307635 175677
rect 307569 175672 310132 175674
rect 213913 175614 217212 175616
rect 307569 175616 307574 175672
rect 307630 175616 310132 175672
rect 307569 175614 310132 175616
rect 213913 175611 213979 175614
rect 307569 175611 307635 175614
rect 104617 175540 104683 175541
rect 120809 175540 120875 175541
rect 130745 175540 130811 175541
rect 98310 175476 98316 175540
rect 98380 175538 98386 175540
rect 104566 175538 104572 175540
rect 98380 175478 103530 175538
rect 104526 175478 104572 175538
rect 104636 175536 104683 175540
rect 120758 175538 120764 175540
rect 104678 175480 104683 175536
rect 98380 175476 98386 175478
rect 103470 175402 103530 175478
rect 104566 175476 104572 175478
rect 104636 175476 104683 175480
rect 120718 175478 120764 175538
rect 120828 175536 120875 175540
rect 130694 175538 130700 175540
rect 120870 175480 120875 175536
rect 120758 175476 120764 175478
rect 120828 175476 120875 175480
rect 130654 175478 130700 175538
rect 130764 175536 130811 175540
rect 130806 175480 130811 175536
rect 321510 175508 321570 175747
rect 130694 175476 130700 175478
rect 130764 175476 130811 175480
rect 104617 175475 104683 175476
rect 120809 175475 120875 175476
rect 130745 175475 130811 175476
rect 170489 175402 170555 175405
rect 103470 175400 170555 175402
rect 103470 175344 170494 175400
rect 170550 175344 170555 175400
rect 103470 175342 170555 175344
rect 170489 175339 170555 175342
rect 250069 175266 250135 175269
rect 248860 175264 250135 175266
rect 248860 175208 250074 175264
rect 250130 175208 250135 175264
rect 248860 175206 250135 175208
rect 250069 175203 250135 175206
rect 307109 175266 307175 175269
rect 321829 175266 321895 175269
rect 307109 175264 310132 175266
rect 307109 175208 307114 175264
rect 307170 175208 310132 175264
rect 307109 175206 310132 175208
rect 321829 175264 321938 175266
rect 321829 175208 321834 175264
rect 321890 175208 321938 175264
rect 307109 175203 307175 175206
rect 321829 175203 321938 175208
rect 115749 174996 115815 174997
rect 115720 174994 115726 174996
rect 115658 174934 115726 174994
rect 115790 174992 115815 174996
rect 115810 174936 115815 174992
rect 115720 174932 115726 174934
rect 115790 174932 115815 174936
rect 115749 174931 115815 174932
rect 213913 174994 213979 174997
rect 213913 174992 217212 174994
rect 213913 174936 213918 174992
rect 213974 174936 217212 174992
rect 213913 174934 217212 174936
rect 213913 174931 213979 174934
rect 306741 174858 306807 174861
rect 306741 174856 310132 174858
rect 306741 174800 306746 174856
rect 306802 174800 310132 174856
rect 306741 174798 310132 174800
rect 306741 174795 306807 174798
rect 249149 174722 249215 174725
rect 248860 174720 249215 174722
rect 248860 174664 249154 174720
rect 249210 174664 249215 174720
rect 321878 174692 321938 175203
rect 248860 174662 249215 174664
rect 249149 174659 249215 174662
rect 165521 174586 165587 174589
rect 214414 174586 214420 174588
rect 165521 174584 214420 174586
rect 165521 174528 165526 174584
rect 165582 174528 214420 174584
rect 165521 174526 214420 174528
rect 165521 174523 165587 174526
rect 214414 174524 214420 174526
rect 214484 174524 214490 174588
rect 307661 174450 307727 174453
rect 307661 174448 310132 174450
rect 307661 174392 307666 174448
rect 307722 174392 310132 174448
rect 307661 174390 310132 174392
rect 307661 174387 307727 174390
rect 214649 174314 214715 174317
rect 249190 174314 249196 174316
rect 214649 174312 217212 174314
rect 214649 174256 214654 174312
rect 214710 174256 217212 174312
rect 214649 174254 217212 174256
rect 248860 174254 249196 174314
rect 214649 174251 214715 174254
rect 249190 174252 249196 174254
rect 249260 174252 249266 174316
rect 307569 174042 307635 174045
rect 324405 174042 324471 174045
rect 307569 174040 310132 174042
rect 307569 173984 307574 174040
rect 307630 173984 310132 174040
rect 307569 173982 310132 173984
rect 321908 174040 324471 174042
rect 321908 173984 324410 174040
rect 324466 173984 324471 174040
rect 321908 173982 324471 173984
rect 307569 173979 307635 173982
rect 324405 173979 324471 173982
rect 249374 173770 249380 173772
rect 248860 173710 249380 173770
rect 249374 173708 249380 173710
rect 249444 173708 249450 173772
rect 213913 173634 213979 173637
rect 306557 173634 306623 173637
rect 213913 173632 217212 173634
rect 213913 173576 213918 173632
rect 213974 173576 217212 173632
rect 213913 173574 217212 173576
rect 306557 173632 310132 173634
rect 306557 173576 306562 173632
rect 306618 173576 310132 173632
rect 306557 173574 310132 173576
rect 213913 173571 213979 173574
rect 306557 173571 306623 173574
rect 249333 173362 249399 173365
rect 248860 173360 249399 173362
rect 248860 173304 249338 173360
rect 249394 173304 249399 173360
rect 248860 173302 249399 173304
rect 249333 173299 249399 173302
rect 306925 173226 306991 173229
rect 324313 173226 324379 173229
rect 306925 173224 310132 173226
rect 306925 173168 306930 173224
rect 306986 173168 310132 173224
rect 306925 173166 310132 173168
rect 321908 173224 324379 173226
rect 321908 173168 324318 173224
rect 324374 173168 324379 173224
rect 321908 173166 324379 173168
rect 306925 173163 306991 173166
rect 324313 173163 324379 173166
rect 214005 172954 214071 172957
rect 214005 172952 217212 172954
rect 214005 172896 214010 172952
rect 214066 172896 217212 172952
rect 214005 172894 217212 172896
rect 214005 172891 214071 172894
rect 252093 172818 252159 172821
rect 248860 172816 252159 172818
rect 248860 172760 252098 172816
rect 252154 172760 252159 172816
rect 248860 172758 252159 172760
rect 252093 172755 252159 172758
rect 307293 172682 307359 172685
rect 321277 172682 321343 172685
rect 307293 172680 310132 172682
rect 307293 172624 307298 172680
rect 307354 172624 310132 172680
rect 307293 172622 310132 172624
rect 321277 172680 321386 172682
rect 321277 172624 321282 172680
rect 321338 172624 321386 172680
rect 307293 172619 307359 172622
rect 321277 172619 321386 172624
rect 249241 172410 249307 172413
rect 248860 172408 249307 172410
rect 248860 172352 249246 172408
rect 249302 172352 249307 172408
rect 321326 172380 321386 172619
rect 248860 172350 249307 172352
rect 249241 172347 249307 172350
rect 213913 172274 213979 172277
rect 306925 172274 306991 172277
rect 213913 172272 217212 172274
rect 213913 172216 213918 172272
rect 213974 172216 217212 172272
rect 213913 172214 217212 172216
rect 306925 172272 310132 172274
rect 306925 172216 306930 172272
rect 306986 172216 310132 172272
rect 306925 172214 310132 172216
rect 213913 172211 213979 172214
rect 306925 172211 306991 172214
rect 321502 172076 321508 172140
rect 321572 172076 321578 172140
rect 252461 171866 252527 171869
rect 248860 171864 252527 171866
rect 248860 171808 252466 171864
rect 252522 171808 252527 171864
rect 248860 171806 252527 171808
rect 252461 171803 252527 171806
rect 307569 171866 307635 171869
rect 307569 171864 310132 171866
rect 307569 171808 307574 171864
rect 307630 171808 310132 171864
rect 307569 171806 310132 171808
rect 307569 171803 307635 171806
rect 321510 171700 321570 172076
rect 168005 171594 168071 171597
rect 164694 171592 168071 171594
rect 164694 171536 168010 171592
rect 168066 171536 168071 171592
rect 164694 171534 168071 171536
rect -960 162890 480 162980
rect 3509 162890 3575 162893
rect -960 162888 3575 162890
rect -960 162832 3514 162888
rect 3570 162832 3575 162888
rect -960 162830 3575 162832
rect -960 162740 480 162830
rect 3509 162827 3575 162830
rect -960 149834 480 149924
rect 3509 149834 3575 149837
rect -960 149832 3575 149834
rect -960 149776 3514 149832
rect 3570 149776 3575 149832
rect -960 149774 3575 149776
rect -960 149684 480 149774
rect 3509 149771 3575 149774
rect -960 136778 480 136868
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 168005 171531 168071 171534
rect 214741 171594 214807 171597
rect 214741 171592 217212 171594
rect 214741 171536 214746 171592
rect 214802 171536 217212 171592
rect 214741 171534 217212 171536
rect 214741 171531 214807 171534
rect 252553 171458 252619 171461
rect 248860 171456 252619 171458
rect 248860 171400 252558 171456
rect 252614 171400 252619 171456
rect 248860 171398 252619 171400
rect 252553 171395 252619 171398
rect 307661 171458 307727 171461
rect 307661 171456 310132 171458
rect 307661 171400 307666 171456
rect 307722 171400 310132 171456
rect 307661 171398 310132 171400
rect 307661 171395 307727 171398
rect 321318 171396 321324 171460
rect 321388 171458 321394 171460
rect 321461 171458 321527 171461
rect 321388 171456 321527 171458
rect 321388 171400 321466 171456
rect 321522 171400 321527 171456
rect 321388 171398 321527 171400
rect 321388 171396 321394 171398
rect 321461 171395 321527 171398
rect 321921 171186 321987 171189
rect 321878 171184 321987 171186
rect 321878 171128 321926 171184
rect 321982 171128 321987 171184
rect 321878 171123 321987 171128
rect 213913 171050 213979 171053
rect 307201 171050 307267 171053
rect 213913 171048 217212 171050
rect 213913 170992 213918 171048
rect 213974 170992 217212 171048
rect 213913 170990 217212 170992
rect 307201 171048 310132 171050
rect 307201 170992 307206 171048
rect 307262 170992 310132 171048
rect 307201 170990 310132 170992
rect 213913 170987 213979 170990
rect 307201 170987 307267 170990
rect 251725 170914 251791 170917
rect 248860 170912 251791 170914
rect 248860 170856 251730 170912
rect 251786 170856 251791 170912
rect 321878 170884 321938 171123
rect 248860 170854 251791 170856
rect 251725 170851 251791 170854
rect 306741 170642 306807 170645
rect 306741 170640 310132 170642
rect 306741 170584 306746 170640
rect 306802 170584 310132 170640
rect 306741 170582 310132 170584
rect 306741 170579 306807 170582
rect 321318 170580 321324 170644
rect 321388 170580 321394 170644
rect 251817 170506 251883 170509
rect 248860 170504 251883 170506
rect 248860 170448 251822 170504
rect 251878 170448 251883 170504
rect 248860 170446 251883 170448
rect 251817 170443 251883 170446
rect 214005 170370 214071 170373
rect 214005 170368 217212 170370
rect 214005 170312 214010 170368
rect 214066 170312 217212 170368
rect 214005 170310 217212 170312
rect 214005 170307 214071 170310
rect 307661 170234 307727 170237
rect 307661 170232 310132 170234
rect 307661 170176 307666 170232
rect 307722 170176 310132 170232
rect 307661 170174 310132 170176
rect 307661 170171 307727 170174
rect 251357 170098 251423 170101
rect 248860 170096 251423 170098
rect 248860 170040 251362 170096
rect 251418 170040 251423 170096
rect 321326 170068 321386 170580
rect 248860 170038 251423 170040
rect 251357 170035 251423 170038
rect 306925 169826 306991 169829
rect 306925 169824 310132 169826
rect 306925 169768 306930 169824
rect 306986 169768 310132 169824
rect 306925 169766 310132 169768
rect 306925 169763 306991 169766
rect 214925 169690 214991 169693
rect 321461 169690 321527 169693
rect 214925 169688 217212 169690
rect 214925 169632 214930 169688
rect 214986 169632 217212 169688
rect 214925 169630 217212 169632
rect 321461 169688 321570 169690
rect 321461 169632 321466 169688
rect 321522 169632 321570 169688
rect 214925 169627 214991 169630
rect 321461 169627 321570 169632
rect 252461 169554 252527 169557
rect 248860 169552 252527 169554
rect 248860 169496 252466 169552
rect 252522 169496 252527 169552
rect 248860 169494 252527 169496
rect 252461 169491 252527 169494
rect 321510 169388 321570 169627
rect 307477 169282 307543 169285
rect 307477 169280 310132 169282
rect 307477 169224 307482 169280
rect 307538 169224 310132 169280
rect 307477 169222 310132 169224
rect 307477 169219 307543 169222
rect 252277 169146 252343 169149
rect 248860 169144 252343 169146
rect 248860 169088 252282 169144
rect 252338 169088 252343 169144
rect 248860 169086 252343 169088
rect 252277 169083 252343 169086
rect 214414 168948 214420 169012
rect 214484 169010 214490 169012
rect 214484 168950 217212 169010
rect 214484 168948 214490 168950
rect 307569 168874 307635 168877
rect 307569 168872 310132 168874
rect 307569 168816 307574 168872
rect 307630 168816 310132 168872
rect 307569 168814 310132 168816
rect 307569 168811 307635 168814
rect 256918 168602 256924 168604
rect 248860 168542 256924 168602
rect 256918 168540 256924 168542
rect 256988 168540 256994 168604
rect 324313 168602 324379 168605
rect 321908 168600 324379 168602
rect 321908 168544 324318 168600
rect 324374 168544 324379 168600
rect 321908 168542 324379 168544
rect 324313 168539 324379 168542
rect 307661 168466 307727 168469
rect 307661 168464 310132 168466
rect 307661 168408 307666 168464
rect 307722 168408 310132 168464
rect 307661 168406 310132 168408
rect 307661 168403 307727 168406
rect 213913 168330 213979 168333
rect 213913 168328 217212 168330
rect 213913 168272 213918 168328
rect 213974 168272 217212 168328
rect 213913 168270 217212 168272
rect 213913 168267 213979 168270
rect 252461 168194 252527 168197
rect 248860 168192 252527 168194
rect 248860 168136 252466 168192
rect 252522 168136 252527 168192
rect 248860 168134 252527 168136
rect 252461 168131 252527 168134
rect 307477 168058 307543 168061
rect 307477 168056 310132 168058
rect 307477 168000 307482 168056
rect 307538 168000 310132 168056
rect 307477 167998 310132 168000
rect 307477 167995 307543 167998
rect 324313 167786 324379 167789
rect 321908 167784 324379 167786
rect 321908 167728 324318 167784
rect 324374 167728 324379 167784
rect 321908 167726 324379 167728
rect 324313 167723 324379 167726
rect 214005 167650 214071 167653
rect 252461 167650 252527 167653
rect 214005 167648 217212 167650
rect 214005 167592 214010 167648
rect 214066 167592 217212 167648
rect 214005 167590 217212 167592
rect 248860 167648 252527 167650
rect 248860 167592 252466 167648
rect 252522 167592 252527 167648
rect 248860 167590 252527 167592
rect 214005 167587 214071 167590
rect 252461 167587 252527 167590
rect 307661 167650 307727 167653
rect 307661 167648 310132 167650
rect 307661 167592 307666 167648
rect 307722 167592 310132 167648
rect 307661 167590 310132 167592
rect 307661 167587 307727 167590
rect 321737 167514 321803 167517
rect 321694 167512 321803 167514
rect 321694 167456 321742 167512
rect 321798 167456 321803 167512
rect 321694 167451 321803 167456
rect 251909 167242 251975 167245
rect 248860 167240 251975 167242
rect 248860 167184 251914 167240
rect 251970 167184 251975 167240
rect 248860 167182 251975 167184
rect 251909 167179 251975 167182
rect 307293 167242 307359 167245
rect 307293 167240 310132 167242
rect 307293 167184 307298 167240
rect 307354 167184 310132 167240
rect 307293 167182 310132 167184
rect 307293 167179 307359 167182
rect 321694 167076 321754 167451
rect 214097 166970 214163 166973
rect 214097 166968 217212 166970
rect 214097 166912 214102 166968
rect 214158 166912 217212 166968
rect 214097 166910 217212 166912
rect 214097 166907 214163 166910
rect 307569 166834 307635 166837
rect 307569 166832 310132 166834
rect 307569 166776 307574 166832
rect 307630 166776 310132 166832
rect 307569 166774 310132 166776
rect 307569 166771 307635 166774
rect 252093 166698 252159 166701
rect 248860 166696 252159 166698
rect 248860 166640 252098 166696
rect 252154 166640 252159 166696
rect 248860 166638 252159 166640
rect 252093 166635 252159 166638
rect 213913 166426 213979 166429
rect 252369 166426 252435 166429
rect 213913 166424 217212 166426
rect 213913 166368 213918 166424
rect 213974 166368 217212 166424
rect 213913 166366 217212 166368
rect 250854 166424 252435 166426
rect 250854 166368 252374 166424
rect 252430 166368 252435 166424
rect 250854 166366 252435 166368
rect 213913 166363 213979 166366
rect 250854 166290 250914 166366
rect 252369 166363 252435 166366
rect 307477 166426 307543 166429
rect 307477 166424 310132 166426
rect 307477 166368 307482 166424
rect 307538 166368 310132 166424
rect 307477 166366 310132 166368
rect 307477 166363 307543 166366
rect 248860 166230 250914 166290
rect 251030 166228 251036 166292
rect 251100 166290 251106 166292
rect 287697 166290 287763 166293
rect 324681 166290 324747 166293
rect 251100 166288 287763 166290
rect 251100 166232 287702 166288
rect 287758 166232 287763 166288
rect 251100 166230 287763 166232
rect 321908 166288 324747 166290
rect 321908 166232 324686 166288
rect 324742 166232 324747 166288
rect 321908 166230 324747 166232
rect 251100 166228 251106 166230
rect 287697 166227 287763 166230
rect 324681 166227 324747 166230
rect 307661 165882 307727 165885
rect 580257 165882 580323 165885
rect 583520 165882 584960 165972
rect 307661 165880 310132 165882
rect 307661 165824 307666 165880
rect 307722 165824 310132 165880
rect 307661 165822 310132 165824
rect 580257 165880 584960 165882
rect 580257 165824 580262 165880
rect 580318 165824 584960 165880
rect 580257 165822 584960 165824
rect 307661 165819 307727 165822
rect 580257 165819 580323 165822
rect 214005 165746 214071 165749
rect 252461 165746 252527 165749
rect 214005 165744 217212 165746
rect 214005 165688 214010 165744
rect 214066 165688 217212 165744
rect 214005 165686 217212 165688
rect 248860 165744 252527 165746
rect 248860 165688 252466 165744
rect 252522 165688 252527 165744
rect 583520 165732 584960 165822
rect 248860 165686 252527 165688
rect 214005 165683 214071 165686
rect 252461 165683 252527 165686
rect 307385 165474 307451 165477
rect 323117 165474 323183 165477
rect 307385 165472 310132 165474
rect 307385 165416 307390 165472
rect 307446 165416 310132 165472
rect 307385 165414 310132 165416
rect 321908 165472 323183 165474
rect 321908 165416 323122 165472
rect 323178 165416 323183 165472
rect 321908 165414 323183 165416
rect 307385 165411 307451 165414
rect 323117 165411 323183 165414
rect 252461 165338 252527 165341
rect 248860 165336 252527 165338
rect 248860 165280 252466 165336
rect 252522 165280 252527 165336
rect 248860 165278 252527 165280
rect 252461 165275 252527 165278
rect 213913 165066 213979 165069
rect 307017 165066 307083 165069
rect 213913 165064 217212 165066
rect 213913 165008 213918 165064
rect 213974 165008 217212 165064
rect 213913 165006 217212 165008
rect 307017 165064 310132 165066
rect 307017 165008 307022 165064
rect 307078 165008 310132 165064
rect 307017 165006 310132 165008
rect 213913 165003 213979 165006
rect 307017 165003 307083 165006
rect 251725 164794 251791 164797
rect 324313 164794 324379 164797
rect 248860 164792 251791 164794
rect 248860 164736 251730 164792
rect 251786 164736 251791 164792
rect 248860 164734 251791 164736
rect 321908 164792 324379 164794
rect 321908 164736 324318 164792
rect 324374 164736 324379 164792
rect 321908 164734 324379 164736
rect 251725 164731 251791 164734
rect 324313 164731 324379 164734
rect 307661 164658 307727 164661
rect 307661 164656 310132 164658
rect 307661 164600 307666 164656
rect 307722 164600 310132 164656
rect 307661 164598 310132 164600
rect 307661 164595 307727 164598
rect 214005 164386 214071 164389
rect 252093 164386 252159 164389
rect 214005 164384 217212 164386
rect 214005 164328 214010 164384
rect 214066 164328 217212 164384
rect 214005 164326 217212 164328
rect 248860 164384 252159 164386
rect 248860 164328 252098 164384
rect 252154 164328 252159 164384
rect 248860 164326 252159 164328
rect 214005 164323 214071 164326
rect 252093 164323 252159 164326
rect 307293 164250 307359 164253
rect 307293 164248 310132 164250
rect 307293 164192 307298 164248
rect 307354 164192 310132 164248
rect 307293 164190 310132 164192
rect 307293 164187 307359 164190
rect 253197 163978 253263 163981
rect 324313 163978 324379 163981
rect 248860 163976 253263 163978
rect 248860 163920 253202 163976
rect 253258 163920 253263 163976
rect 248860 163918 253263 163920
rect 321908 163976 324379 163978
rect 321908 163920 324318 163976
rect 324374 163920 324379 163976
rect 321908 163918 324379 163920
rect 253197 163915 253263 163918
rect 324313 163915 324379 163918
rect 306741 163842 306807 163845
rect 306741 163840 310132 163842
rect 306741 163784 306746 163840
rect 306802 163784 310132 163840
rect 306741 163782 310132 163784
rect 306741 163779 306807 163782
rect 213913 163706 213979 163709
rect 213913 163704 217212 163706
rect 213913 163648 213918 163704
rect 213974 163648 217212 163704
rect 213913 163646 217212 163648
rect 213913 163643 213979 163646
rect 307661 163434 307727 163437
rect 248860 163374 258090 163434
rect 258030 163162 258090 163374
rect 307661 163432 310132 163434
rect 307661 163376 307666 163432
rect 307722 163376 310132 163432
rect 307661 163374 310132 163376
rect 307661 163371 307727 163374
rect 269062 163162 269068 163164
rect 258030 163102 269068 163162
rect 269062 163100 269068 163102
rect 269132 163100 269138 163164
rect 324405 163162 324471 163165
rect 321908 163160 324471 163162
rect 321908 163104 324410 163160
rect 324466 163104 324471 163160
rect 321908 163102 324471 163104
rect 324405 163099 324471 163102
rect 214005 163026 214071 163029
rect 252185 163026 252251 163029
rect 214005 163024 217212 163026
rect 214005 162968 214010 163024
rect 214066 162968 217212 163024
rect 214005 162966 217212 162968
rect 248860 163024 252251 163026
rect 248860 162968 252190 163024
rect 252246 162968 252251 163024
rect 248860 162966 252251 162968
rect 214005 162963 214071 162966
rect 252185 162963 252251 162966
rect 253197 163026 253263 163029
rect 266302 163026 266308 163028
rect 253197 163024 266308 163026
rect 253197 162968 253202 163024
rect 253258 162968 266308 163024
rect 253197 162966 266308 162968
rect 253197 162963 253263 162966
rect 266302 162964 266308 162966
rect 266372 162964 266378 163028
rect 307293 163026 307359 163029
rect 307293 163024 310132 163026
rect 307293 162968 307298 163024
rect 307354 162968 310132 163024
rect 307293 162966 310132 162968
rect 307293 162963 307359 162966
rect 252461 162482 252527 162485
rect 248860 162480 252527 162482
rect 248860 162424 252466 162480
rect 252522 162424 252527 162480
rect 248860 162422 252527 162424
rect 252461 162419 252527 162422
rect 307477 162482 307543 162485
rect 324313 162482 324379 162485
rect 307477 162480 310132 162482
rect 307477 162424 307482 162480
rect 307538 162424 310132 162480
rect 307477 162422 310132 162424
rect 321908 162480 324379 162482
rect 321908 162424 324318 162480
rect 324374 162424 324379 162480
rect 321908 162422 324379 162424
rect 307477 162419 307543 162422
rect 324313 162419 324379 162422
rect 213913 162346 213979 162349
rect 213913 162344 217212 162346
rect 213913 162288 213918 162344
rect 213974 162288 217212 162344
rect 213913 162286 217212 162288
rect 213913 162283 213979 162286
rect 265014 162210 265020 162212
rect 258030 162150 265020 162210
rect 258030 162074 258090 162150
rect 265014 162148 265020 162150
rect 265084 162148 265090 162212
rect 248860 162014 258090 162074
rect 262213 162074 262279 162077
rect 275134 162074 275140 162076
rect 262213 162072 275140 162074
rect 262213 162016 262218 162072
rect 262274 162016 275140 162072
rect 262213 162014 275140 162016
rect 262213 162011 262279 162014
rect 275134 162012 275140 162014
rect 275204 162012 275210 162076
rect 307661 162074 307727 162077
rect 307661 162072 310132 162074
rect 307661 162016 307666 162072
rect 307722 162016 310132 162072
rect 307661 162014 310132 162016
rect 307661 162011 307727 162014
rect 214005 161802 214071 161805
rect 214005 161800 217212 161802
rect 214005 161744 214010 161800
rect 214066 161744 217212 161800
rect 214005 161742 217212 161744
rect 214005 161739 214071 161742
rect 306465 161666 306531 161669
rect 324405 161666 324471 161669
rect 306465 161664 310132 161666
rect 306465 161608 306470 161664
rect 306526 161608 310132 161664
rect 306465 161606 310132 161608
rect 321908 161664 324471 161666
rect 321908 161608 324410 161664
rect 324466 161608 324471 161664
rect 321908 161606 324471 161608
rect 306465 161603 306531 161606
rect 324405 161603 324471 161606
rect 260782 161530 260788 161532
rect 248860 161470 260788 161530
rect 260782 161468 260788 161470
rect 260852 161468 260858 161532
rect 307569 161258 307635 161261
rect 307569 161256 310132 161258
rect 307569 161200 307574 161256
rect 307630 161200 310132 161256
rect 307569 161198 310132 161200
rect 307569 161195 307635 161198
rect 214557 161122 214623 161125
rect 256734 161122 256740 161124
rect 214557 161120 217212 161122
rect 214557 161064 214562 161120
rect 214618 161064 217212 161120
rect 214557 161062 217212 161064
rect 248860 161062 256740 161122
rect 214557 161059 214623 161062
rect 256734 161060 256740 161062
rect 256804 161060 256810 161124
rect 307661 160850 307727 160853
rect 324313 160850 324379 160853
rect 307661 160848 310132 160850
rect 307661 160792 307666 160848
rect 307722 160792 310132 160848
rect 307661 160790 310132 160792
rect 321908 160848 324379 160850
rect 321908 160792 324318 160848
rect 324374 160792 324379 160848
rect 321908 160790 324379 160792
rect 307661 160787 307727 160790
rect 324313 160787 324379 160790
rect 166206 160652 166212 160716
rect 166276 160714 166282 160716
rect 214097 160714 214163 160717
rect 166276 160712 214163 160714
rect 166276 160656 214102 160712
rect 214158 160656 214163 160712
rect 166276 160654 214163 160656
rect 166276 160652 166282 160654
rect 214097 160651 214163 160654
rect 252461 160578 252527 160581
rect 248860 160576 252527 160578
rect 248860 160520 252466 160576
rect 252522 160520 252527 160576
rect 248860 160518 252527 160520
rect 252461 160515 252527 160518
rect 213913 160442 213979 160445
rect 306557 160442 306623 160445
rect 213913 160440 217212 160442
rect 213913 160384 213918 160440
rect 213974 160384 217212 160440
rect 213913 160382 217212 160384
rect 306557 160440 310132 160442
rect 306557 160384 306562 160440
rect 306618 160384 310132 160440
rect 306557 160382 310132 160384
rect 213913 160379 213979 160382
rect 306557 160379 306623 160382
rect 251357 160170 251423 160173
rect 324405 160170 324471 160173
rect 248860 160168 251423 160170
rect 248860 160112 251362 160168
rect 251418 160112 251423 160168
rect 248860 160110 251423 160112
rect 321908 160168 324471 160170
rect 321908 160112 324410 160168
rect 324466 160112 324471 160168
rect 321908 160110 324471 160112
rect 251357 160107 251423 160110
rect 324405 160107 324471 160110
rect 306925 160034 306991 160037
rect 306925 160032 310132 160034
rect 306925 159976 306930 160032
rect 306986 159976 310132 160032
rect 306925 159974 310132 159976
rect 306925 159971 306991 159974
rect 213913 159762 213979 159765
rect 213913 159760 217212 159762
rect 213913 159704 213918 159760
rect 213974 159704 217212 159760
rect 213913 159702 217212 159704
rect 213913 159699 213979 159702
rect 251265 159626 251331 159629
rect 248860 159624 251331 159626
rect 248860 159568 251270 159624
rect 251326 159568 251331 159624
rect 248860 159566 251331 159568
rect 251265 159563 251331 159566
rect 307109 159626 307175 159629
rect 307109 159624 310132 159626
rect 307109 159568 307114 159624
rect 307170 159568 310132 159624
rect 307109 159566 310132 159568
rect 307109 159563 307175 159566
rect 324313 159354 324379 159357
rect 321908 159352 324379 159354
rect 321908 159296 324318 159352
rect 324374 159296 324379 159352
rect 321908 159294 324379 159296
rect 324313 159291 324379 159294
rect 250069 159218 250135 159221
rect 248860 159216 250135 159218
rect 248860 159160 250074 159216
rect 250130 159160 250135 159216
rect 248860 159158 250135 159160
rect 250069 159155 250135 159158
rect 214005 159082 214071 159085
rect 307661 159082 307727 159085
rect 214005 159080 217212 159082
rect 214005 159024 214010 159080
rect 214066 159024 217212 159080
rect 214005 159022 217212 159024
rect 307661 159080 310132 159082
rect 307661 159024 307666 159080
rect 307722 159024 310132 159080
rect 307661 159022 310132 159024
rect 214005 159019 214071 159022
rect 307661 159019 307727 159022
rect 251173 158810 251239 158813
rect 248860 158808 251239 158810
rect 248860 158752 251178 158808
rect 251234 158752 251239 158808
rect 248860 158750 251239 158752
rect 251173 158747 251239 158750
rect 306925 158674 306991 158677
rect 306925 158672 310132 158674
rect 306925 158616 306930 158672
rect 306986 158616 310132 158672
rect 306925 158614 310132 158616
rect 306925 158611 306991 158614
rect 324313 158538 324379 158541
rect 321908 158536 324379 158538
rect 321908 158480 324318 158536
rect 324374 158480 324379 158536
rect 321908 158478 324379 158480
rect 324313 158475 324379 158478
rect 214649 158402 214715 158405
rect 214649 158400 217212 158402
rect 214649 158344 214654 158400
rect 214710 158344 217212 158400
rect 214649 158342 217212 158344
rect 214649 158339 214715 158342
rect 255446 158266 255452 158268
rect 248860 158206 255452 158266
rect 255446 158204 255452 158206
rect 255516 158204 255522 158268
rect 307477 158266 307543 158269
rect 307477 158264 310132 158266
rect 307477 158208 307482 158264
rect 307538 158208 310132 158264
rect 307477 158206 310132 158208
rect 307477 158203 307543 158206
rect 251909 157858 251975 157861
rect 248860 157856 251975 157858
rect 248860 157800 251914 157856
rect 251970 157800 251975 157856
rect 248860 157798 251975 157800
rect 251909 157795 251975 157798
rect 307661 157858 307727 157861
rect 324405 157858 324471 157861
rect 307661 157856 310132 157858
rect 307661 157800 307666 157856
rect 307722 157800 310132 157856
rect 307661 157798 310132 157800
rect 321908 157856 324471 157858
rect 321908 157800 324410 157856
rect 324466 157800 324471 157856
rect 321908 157798 324471 157800
rect 307661 157795 307727 157798
rect 324405 157795 324471 157798
rect 213913 157722 213979 157725
rect 213913 157720 217212 157722
rect 213913 157664 213918 157720
rect 213974 157664 217212 157720
rect 213913 157662 217212 157664
rect 213913 157659 213979 157662
rect 307150 157388 307156 157452
rect 307220 157450 307226 157452
rect 307220 157390 310132 157450
rect 307220 157388 307226 157390
rect 252461 157314 252527 157317
rect 248860 157312 252527 157314
rect 248860 157256 252466 157312
rect 252522 157256 252527 157312
rect 248860 157254 252527 157256
rect 252461 157251 252527 157254
rect 214097 157178 214163 157181
rect 214097 157176 217212 157178
rect 214097 157120 214102 157176
rect 214158 157120 217212 157176
rect 214097 157118 217212 157120
rect 214097 157115 214163 157118
rect 307477 157042 307543 157045
rect 324313 157042 324379 157045
rect 307477 157040 310132 157042
rect 307477 156984 307482 157040
rect 307538 156984 310132 157040
rect 307477 156982 310132 156984
rect 321908 157040 324379 157042
rect 321908 156984 324318 157040
rect 324374 156984 324379 157040
rect 321908 156982 324379 156984
rect 307477 156979 307543 156982
rect 324313 156979 324379 156982
rect 251541 156906 251607 156909
rect 248860 156904 251607 156906
rect 248860 156848 251546 156904
rect 251602 156848 251607 156904
rect 248860 156846 251607 156848
rect 251541 156843 251607 156846
rect 307569 156634 307635 156637
rect 307569 156632 310132 156634
rect 307569 156576 307574 156632
rect 307630 156576 310132 156632
rect 307569 156574 310132 156576
rect 307569 156571 307635 156574
rect 213913 156498 213979 156501
rect 213913 156496 217212 156498
rect 213913 156440 213918 156496
rect 213974 156440 217212 156496
rect 213913 156438 217212 156440
rect 213913 156435 213979 156438
rect 252369 156362 252435 156365
rect 325877 156362 325943 156365
rect 248860 156360 252435 156362
rect 248860 156304 252374 156360
rect 252430 156304 252435 156360
rect 248860 156302 252435 156304
rect 321908 156360 325943 156362
rect 321908 156304 325882 156360
rect 325938 156304 325943 156360
rect 321908 156302 325943 156304
rect 252369 156299 252435 156302
rect 325877 156299 325943 156302
rect 307661 156226 307727 156229
rect 307661 156224 310132 156226
rect 307661 156168 307666 156224
rect 307722 156168 310132 156224
rect 307661 156166 310132 156168
rect 307661 156163 307727 156166
rect 251909 155954 251975 155957
rect 248860 155952 251975 155954
rect 248860 155896 251914 155952
rect 251970 155896 251975 155952
rect 248860 155894 251975 155896
rect 251909 155891 251975 155894
rect 213913 155818 213979 155821
rect 213913 155816 217212 155818
rect 213913 155760 213918 155816
rect 213974 155760 217212 155816
rect 213913 155758 217212 155760
rect 213913 155755 213979 155758
rect 307661 155682 307727 155685
rect 307661 155680 310132 155682
rect 307661 155624 307666 155680
rect 307722 155624 310132 155680
rect 307661 155622 310132 155624
rect 307661 155619 307727 155622
rect 324313 155546 324379 155549
rect 321908 155544 324379 155546
rect 321908 155488 324318 155544
rect 324374 155488 324379 155544
rect 321908 155486 324379 155488
rect 324313 155483 324379 155486
rect 251173 155410 251239 155413
rect 248860 155408 251239 155410
rect 248860 155352 251178 155408
rect 251234 155352 251239 155408
rect 248860 155350 251239 155352
rect 251173 155347 251239 155350
rect 307477 155274 307543 155277
rect 307477 155272 310132 155274
rect 307477 155216 307482 155272
rect 307538 155216 310132 155272
rect 307477 155214 310132 155216
rect 307477 155211 307543 155214
rect 214005 155138 214071 155141
rect 214005 155136 217212 155138
rect 214005 155080 214010 155136
rect 214066 155080 217212 155136
rect 214005 155078 217212 155080
rect 214005 155075 214071 155078
rect 252461 155002 252527 155005
rect 248860 155000 252527 155002
rect 248860 154944 252466 155000
rect 252522 154944 252527 155000
rect 248860 154942 252527 154944
rect 252461 154939 252527 154942
rect 306966 154804 306972 154868
rect 307036 154866 307042 154868
rect 307036 154806 310132 154866
rect 307036 154804 307042 154806
rect 324405 154730 324471 154733
rect 321908 154728 324471 154730
rect 321908 154672 324410 154728
rect 324466 154672 324471 154728
rect 321908 154670 324471 154672
rect 324405 154667 324471 154670
rect 214005 154458 214071 154461
rect 251081 154458 251147 154461
rect 214005 154456 217212 154458
rect 214005 154400 214010 154456
rect 214066 154400 217212 154456
rect 214005 154398 217212 154400
rect 248860 154456 251147 154458
rect 248860 154400 251086 154456
rect 251142 154400 251147 154456
rect 248860 154398 251147 154400
rect 214005 154395 214071 154398
rect 251081 154395 251147 154398
rect 307569 154458 307635 154461
rect 307569 154456 310132 154458
rect 307569 154400 307574 154456
rect 307630 154400 310132 154456
rect 307569 154398 310132 154400
rect 307569 154395 307635 154398
rect 251633 154050 251699 154053
rect 248860 154048 251699 154050
rect 248860 153992 251638 154048
rect 251694 153992 251699 154048
rect 248860 153990 251699 153992
rect 251633 153987 251699 153990
rect 307477 154050 307543 154053
rect 324313 154050 324379 154053
rect 307477 154048 310132 154050
rect 307477 153992 307482 154048
rect 307538 153992 310132 154048
rect 307477 153990 310132 153992
rect 321908 154048 324379 154050
rect 321908 153992 324318 154048
rect 324374 153992 324379 154048
rect 321908 153990 324379 153992
rect 307477 153987 307543 153990
rect 324313 153987 324379 153990
rect 213913 153778 213979 153781
rect 213913 153776 217212 153778
rect 213913 153720 213918 153776
rect 213974 153720 217212 153776
rect 213913 153718 217212 153720
rect 213913 153715 213979 153718
rect 307661 153642 307727 153645
rect 307661 153640 310132 153642
rect 307661 153584 307666 153640
rect 307722 153584 310132 153640
rect 307661 153582 310132 153584
rect 307661 153579 307727 153582
rect 252461 153506 252527 153509
rect 248860 153504 252527 153506
rect 248860 153448 252466 153504
rect 252522 153448 252527 153504
rect 248860 153446 252527 153448
rect 252461 153443 252527 153446
rect 307201 153234 307267 153237
rect 324313 153234 324379 153237
rect 307201 153232 310132 153234
rect 307201 153176 307206 153232
rect 307262 153176 310132 153232
rect 307201 153174 310132 153176
rect 321908 153232 324379 153234
rect 321908 153176 324318 153232
rect 324374 153176 324379 153232
rect 321908 153174 324379 153176
rect 307201 153171 307267 153174
rect 324313 153171 324379 153174
rect 213913 153098 213979 153101
rect 252461 153098 252527 153101
rect 213913 153096 217212 153098
rect 213913 153040 213918 153096
rect 213974 153040 217212 153096
rect 213913 153038 217212 153040
rect 248860 153096 252527 153098
rect 248860 153040 252466 153096
rect 252522 153040 252527 153096
rect 248860 153038 252527 153040
rect 213913 153035 213979 153038
rect 252461 153035 252527 153038
rect 250529 152962 250595 152965
rect 257838 152962 257844 152964
rect 250529 152960 257844 152962
rect 250529 152904 250534 152960
rect 250590 152904 257844 152960
rect 250529 152902 257844 152904
rect 250529 152899 250595 152902
rect 257838 152900 257844 152902
rect 257908 152900 257914 152964
rect 252369 152690 252435 152693
rect 248860 152688 252435 152690
rect 248860 152632 252374 152688
rect 252430 152632 252435 152688
rect 248860 152630 252435 152632
rect 252369 152627 252435 152630
rect 306649 152690 306715 152693
rect 580349 152690 580415 152693
rect 583520 152690 584960 152780
rect 306649 152688 310132 152690
rect 306649 152632 306654 152688
rect 306710 152632 310132 152688
rect 306649 152630 310132 152632
rect 580349 152688 584960 152690
rect 580349 152632 580354 152688
rect 580410 152632 584960 152688
rect 580349 152630 584960 152632
rect 306649 152627 306715 152630
rect 580349 152627 580415 152630
rect 214005 152554 214071 152557
rect 214005 152552 217212 152554
rect 214005 152496 214010 152552
rect 214066 152496 217212 152552
rect 583520 152540 584960 152630
rect 214005 152494 217212 152496
rect 214005 152491 214071 152494
rect 324497 152418 324563 152421
rect 321908 152416 324563 152418
rect 321908 152360 324502 152416
rect 324558 152360 324563 152416
rect 321908 152358 324563 152360
rect 324497 152355 324563 152358
rect 307569 152282 307635 152285
rect 307569 152280 310132 152282
rect 307569 152224 307574 152280
rect 307630 152224 310132 152280
rect 307569 152222 310132 152224
rect 307569 152219 307635 152222
rect 251909 152146 251975 152149
rect 248860 152144 251975 152146
rect 248860 152088 251914 152144
rect 251970 152088 251975 152144
rect 248860 152086 251975 152088
rect 251909 152083 251975 152086
rect 214373 151874 214439 151877
rect 307661 151874 307727 151877
rect 214373 151872 217212 151874
rect 214373 151816 214378 151872
rect 214434 151816 217212 151872
rect 214373 151814 217212 151816
rect 307661 151872 310132 151874
rect 307661 151816 307666 151872
rect 307722 151816 310132 151872
rect 307661 151814 310132 151816
rect 214373 151811 214439 151814
rect 307661 151811 307727 151814
rect 252461 151738 252527 151741
rect 324313 151738 324379 151741
rect 248860 151736 252527 151738
rect 248860 151680 252466 151736
rect 252522 151680 252527 151736
rect 248860 151678 252527 151680
rect 321908 151736 324379 151738
rect 321908 151680 324318 151736
rect 324374 151680 324379 151736
rect 321908 151678 324379 151680
rect 252461 151675 252527 151678
rect 324313 151675 324379 151678
rect 307477 151466 307543 151469
rect 307477 151464 310132 151466
rect 307477 151408 307482 151464
rect 307538 151408 310132 151464
rect 307477 151406 310132 151408
rect 307477 151403 307543 151406
rect 214005 151194 214071 151197
rect 252369 151194 252435 151197
rect 214005 151192 217212 151194
rect 214005 151136 214010 151192
rect 214066 151136 217212 151192
rect 214005 151134 217212 151136
rect 248860 151192 252435 151194
rect 248860 151136 252374 151192
rect 252430 151136 252435 151192
rect 248860 151134 252435 151136
rect 214005 151131 214071 151134
rect 252369 151131 252435 151134
rect 307661 151058 307727 151061
rect 307661 151056 310132 151058
rect 307661 151000 307666 151056
rect 307722 151000 310132 151056
rect 307661 150998 310132 151000
rect 307661 150995 307727 150998
rect 323025 150922 323091 150925
rect 321908 150920 323091 150922
rect 321908 150864 323030 150920
rect 323086 150864 323091 150920
rect 321908 150862 323091 150864
rect 323025 150859 323091 150862
rect 251909 150786 251975 150789
rect 248860 150784 251975 150786
rect 248860 150728 251914 150784
rect 251970 150728 251975 150784
rect 248860 150726 251975 150728
rect 251909 150723 251975 150726
rect 306741 150650 306807 150653
rect 306741 150648 310132 150650
rect 306741 150592 306746 150648
rect 306802 150592 310132 150648
rect 306741 150590 310132 150592
rect 306741 150587 306807 150590
rect 213913 150514 213979 150517
rect 213913 150512 217212 150514
rect 213913 150456 213918 150512
rect 213974 150456 217212 150512
rect 213913 150454 217212 150456
rect 213913 150451 213979 150454
rect 321645 150378 321711 150381
rect 321645 150376 321754 150378
rect 321645 150320 321650 150376
rect 321706 150320 321754 150376
rect 321645 150315 321754 150320
rect 252461 150242 252527 150245
rect 248860 150240 252527 150242
rect 248860 150184 252466 150240
rect 252522 150184 252527 150240
rect 248860 150182 252527 150184
rect 252461 150179 252527 150182
rect 307569 150242 307635 150245
rect 307569 150240 310132 150242
rect 307569 150184 307574 150240
rect 307630 150184 310132 150240
rect 307569 150182 310132 150184
rect 307569 150179 307635 150182
rect 321694 150076 321754 150315
rect 214005 149834 214071 149837
rect 251173 149834 251239 149837
rect 214005 149832 217212 149834
rect 214005 149776 214010 149832
rect 214066 149776 217212 149832
rect 214005 149774 217212 149776
rect 248860 149832 251239 149834
rect 248860 149776 251178 149832
rect 251234 149776 251239 149832
rect 248860 149774 251239 149776
rect 214005 149771 214071 149774
rect 251173 149771 251239 149774
rect 306741 149834 306807 149837
rect 306741 149832 310132 149834
rect 306741 149776 306746 149832
rect 306802 149776 310132 149832
rect 306741 149774 310132 149776
rect 306741 149771 306807 149774
rect 251950 149636 251956 149700
rect 252020 149698 252026 149700
rect 300761 149698 300827 149701
rect 252020 149696 300827 149698
rect 252020 149640 300766 149696
rect 300822 149640 300827 149696
rect 252020 149638 300827 149640
rect 252020 149636 252026 149638
rect 300761 149635 300827 149638
rect 324313 149426 324379 149429
rect 321908 149424 324379 149426
rect 321908 149368 324318 149424
rect 324374 149368 324379 149424
rect 321908 149366 324379 149368
rect 324313 149363 324379 149366
rect 252001 149290 252067 149293
rect 248860 149288 252067 149290
rect 248860 149232 252006 149288
rect 252062 149232 252067 149288
rect 248860 149230 252067 149232
rect 252001 149227 252067 149230
rect 307661 149290 307727 149293
rect 307661 149288 310132 149290
rect 307661 149232 307666 149288
rect 307722 149232 310132 149288
rect 307661 149230 310132 149232
rect 307661 149227 307727 149230
rect 213913 149154 213979 149157
rect 213913 149152 217212 149154
rect 213913 149096 213918 149152
rect 213974 149096 217212 149152
rect 213913 149094 217212 149096
rect 213913 149091 213979 149094
rect 251909 148882 251975 148885
rect 248860 148880 251975 148882
rect 248860 148824 251914 148880
rect 251970 148824 251975 148880
rect 248860 148822 251975 148824
rect 251909 148819 251975 148822
rect 307569 148882 307635 148885
rect 307569 148880 310132 148882
rect 307569 148824 307574 148880
rect 307630 148824 310132 148880
rect 307569 148822 310132 148824
rect 307569 148819 307635 148822
rect 324313 148610 324379 148613
rect 321908 148608 324379 148610
rect 321908 148552 324318 148608
rect 324374 148552 324379 148608
rect 321908 148550 324379 148552
rect 324313 148547 324379 148550
rect 213913 148474 213979 148477
rect 307385 148474 307451 148477
rect 213913 148472 217212 148474
rect 213913 148416 213918 148472
rect 213974 148416 217212 148472
rect 213913 148414 217212 148416
rect 307385 148472 310132 148474
rect 307385 148416 307390 148472
rect 307446 148416 310132 148472
rect 307385 148414 310132 148416
rect 213913 148411 213979 148414
rect 307385 148411 307451 148414
rect 252461 148338 252527 148341
rect 248860 148336 252527 148338
rect 248860 148280 252466 148336
rect 252522 148280 252527 148336
rect 248860 148278 252527 148280
rect 252461 148275 252527 148278
rect 257521 148338 257587 148341
rect 307150 148338 307156 148340
rect 257521 148336 307156 148338
rect 257521 148280 257526 148336
rect 257582 148280 307156 148336
rect 257521 148278 307156 148280
rect 257521 148275 257587 148278
rect 307150 148276 307156 148278
rect 307220 148276 307226 148340
rect 307661 148066 307727 148069
rect 307661 148064 310132 148066
rect 307661 148008 307666 148064
rect 307722 148008 310132 148064
rect 307661 148006 310132 148008
rect 307661 148003 307727 148006
rect 213913 147930 213979 147933
rect 252502 147930 252508 147932
rect 213913 147928 217212 147930
rect 213913 147872 213918 147928
rect 213974 147872 217212 147928
rect 213913 147870 217212 147872
rect 248860 147870 252508 147930
rect 213913 147867 213979 147870
rect 252502 147868 252508 147870
rect 252572 147868 252578 147932
rect 324405 147794 324471 147797
rect 321908 147792 324471 147794
rect 321908 147736 324410 147792
rect 324466 147736 324471 147792
rect 321908 147734 324471 147736
rect 324405 147731 324471 147734
rect 307293 147658 307359 147661
rect 307293 147656 310132 147658
rect 307293 147600 307298 147656
rect 307354 147600 310132 147656
rect 307293 147598 310132 147600
rect 307293 147595 307359 147598
rect 252461 147522 252527 147525
rect 248860 147520 252527 147522
rect 248860 147464 252466 147520
rect 252522 147464 252527 147520
rect 248860 147462 252527 147464
rect 252461 147459 252527 147462
rect 214005 147250 214071 147253
rect 307477 147250 307543 147253
rect 214005 147248 217212 147250
rect 214005 147192 214010 147248
rect 214066 147192 217212 147248
rect 214005 147190 217212 147192
rect 307477 147248 310132 147250
rect 307477 147192 307482 147248
rect 307538 147192 310132 147248
rect 307477 147190 310132 147192
rect 214005 147187 214071 147190
rect 307477 147187 307543 147190
rect 324313 147114 324379 147117
rect 321908 147112 324379 147114
rect 321908 147056 324318 147112
rect 324374 147056 324379 147112
rect 321908 147054 324379 147056
rect 324313 147051 324379 147054
rect 254526 146978 254532 146980
rect 248860 146918 254532 146978
rect 254526 146916 254532 146918
rect 254596 146916 254602 146980
rect 307569 146842 307635 146845
rect 307569 146840 310132 146842
rect 307569 146784 307574 146840
rect 307630 146784 310132 146840
rect 307569 146782 310132 146784
rect 307569 146779 307635 146782
rect 213913 146570 213979 146573
rect 252369 146570 252435 146573
rect 213913 146568 217212 146570
rect 213913 146512 213918 146568
rect 213974 146512 217212 146568
rect 213913 146510 217212 146512
rect 248860 146568 252435 146570
rect 248860 146512 252374 146568
rect 252430 146512 252435 146568
rect 248860 146510 252435 146512
rect 213913 146507 213979 146510
rect 252369 146507 252435 146510
rect 307661 146434 307727 146437
rect 307661 146432 310132 146434
rect 307661 146376 307666 146432
rect 307722 146376 310132 146432
rect 307661 146374 310132 146376
rect 307661 146371 307727 146374
rect 252461 146026 252527 146029
rect 248860 146024 252527 146026
rect 248860 145968 252466 146024
rect 252522 145968 252527 146024
rect 248860 145966 252527 145968
rect 252461 145963 252527 145966
rect 214005 145890 214071 145893
rect 307477 145890 307543 145893
rect 214005 145888 217212 145890
rect 214005 145832 214010 145888
rect 214066 145832 217212 145888
rect 214005 145830 217212 145832
rect 307477 145888 310132 145890
rect 307477 145832 307482 145888
rect 307538 145832 310132 145888
rect 307477 145830 310132 145832
rect 214005 145827 214071 145830
rect 307477 145827 307543 145830
rect 252277 145618 252343 145621
rect 248860 145616 252343 145618
rect 248860 145560 252282 145616
rect 252338 145560 252343 145616
rect 248860 145558 252343 145560
rect 321878 145618 321938 146268
rect 335670 145618 335676 145620
rect 321878 145558 335676 145618
rect 252277 145555 252343 145558
rect 335670 145556 335676 145558
rect 335740 145556 335746 145620
rect 307661 145482 307727 145485
rect 327206 145482 327212 145484
rect 307661 145480 310132 145482
rect 307661 145424 307666 145480
rect 307722 145424 310132 145480
rect 307661 145422 310132 145424
rect 321908 145422 327212 145482
rect 307661 145419 307727 145422
rect 327206 145420 327212 145422
rect 327276 145420 327282 145484
rect 213913 145210 213979 145213
rect 213913 145208 217212 145210
rect 213913 145152 213918 145208
rect 213974 145152 217212 145208
rect 213913 145150 217212 145152
rect 213913 145147 213979 145150
rect 252093 145074 252159 145077
rect 248860 145072 252159 145074
rect 248860 145016 252098 145072
rect 252154 145016 252159 145072
rect 248860 145014 252159 145016
rect 252093 145011 252159 145014
rect 307109 145074 307175 145077
rect 307109 145072 310132 145074
rect 307109 145016 307114 145072
rect 307170 145016 310132 145072
rect 307109 145014 310132 145016
rect 307109 145011 307175 145014
rect 321908 144742 322122 144802
rect 263542 144666 263548 144668
rect 248860 144606 263548 144666
rect 263542 144604 263548 144606
rect 263612 144604 263618 144668
rect 307569 144666 307635 144669
rect 322062 144668 322122 144742
rect 307569 144664 310132 144666
rect 307569 144608 307574 144664
rect 307630 144608 310132 144664
rect 307569 144606 310132 144608
rect 307569 144603 307635 144606
rect 322054 144604 322060 144668
rect 322124 144604 322130 144668
rect 214005 144530 214071 144533
rect 214005 144528 217212 144530
rect 214005 144472 214010 144528
rect 214066 144472 217212 144528
rect 214005 144470 217212 144472
rect 214005 144467 214071 144470
rect 307661 144258 307727 144261
rect 307661 144256 310132 144258
rect 307661 144200 307666 144256
rect 307722 144200 310132 144256
rect 307661 144198 310132 144200
rect 307661 144195 307727 144198
rect 252461 144122 252527 144125
rect 248860 144120 252527 144122
rect 248860 144064 252466 144120
rect 252522 144064 252527 144120
rect 248860 144062 252527 144064
rect 252461 144059 252527 144062
rect 258993 144122 259059 144125
rect 306966 144122 306972 144124
rect 258993 144120 306972 144122
rect 258993 144064 258998 144120
rect 259054 144064 306972 144120
rect 258993 144062 306972 144064
rect 258993 144059 259059 144062
rect 306966 144060 306972 144062
rect 307036 144060 307042 144124
rect 324313 143986 324379 143989
rect 321908 143984 324379 143986
rect 321908 143928 324318 143984
rect 324374 143928 324379 143984
rect 321908 143926 324379 143928
rect 324313 143923 324379 143926
rect 213913 143850 213979 143853
rect 306649 143850 306715 143853
rect 213913 143848 217212 143850
rect 213913 143792 213918 143848
rect 213974 143792 217212 143848
rect 213913 143790 217212 143792
rect 306649 143848 310132 143850
rect 306649 143792 306654 143848
rect 306710 143792 310132 143848
rect 306649 143790 310132 143792
rect 213913 143787 213979 143790
rect 306649 143787 306715 143790
rect 252093 143714 252159 143717
rect 248860 143712 252159 143714
rect 248860 143656 252098 143712
rect 252154 143656 252159 143712
rect 248860 143654 252159 143656
rect 252093 143651 252159 143654
rect 305729 143714 305795 143717
rect 307569 143714 307635 143717
rect 305729 143712 307635 143714
rect 305729 143656 305734 143712
rect 305790 143656 307574 143712
rect 307630 143656 307635 143712
rect 305729 143654 307635 143656
rect 305729 143651 305795 143654
rect 307569 143651 307635 143654
rect 306557 143442 306623 143445
rect 306557 143440 310132 143442
rect 306557 143384 306562 143440
rect 306618 143384 310132 143440
rect 306557 143382 310132 143384
rect 306557 143379 306623 143382
rect 213913 143306 213979 143309
rect 213913 143304 217212 143306
rect 213913 143248 213918 143304
rect 213974 143248 217212 143304
rect 213913 143246 217212 143248
rect 213913 143243 213979 143246
rect 251817 143170 251883 143173
rect 324313 143170 324379 143173
rect 248860 143168 251883 143170
rect 248860 143112 251822 143168
rect 251878 143112 251883 143168
rect 248860 143110 251883 143112
rect 321908 143168 324379 143170
rect 321908 143112 324318 143168
rect 324374 143112 324379 143168
rect 321908 143110 324379 143112
rect 251817 143107 251883 143110
rect 324313 143107 324379 143110
rect 307569 143034 307635 143037
rect 307569 143032 310132 143034
rect 307569 142976 307574 143032
rect 307630 142976 310132 143032
rect 307569 142974 310132 142976
rect 307569 142971 307635 142974
rect 252277 142762 252343 142765
rect 248860 142760 252343 142762
rect 248860 142704 252282 142760
rect 252338 142704 252343 142760
rect 248860 142702 252343 142704
rect 252277 142699 252343 142702
rect 214741 142626 214807 142629
rect 214741 142624 217212 142626
rect 214741 142568 214746 142624
rect 214802 142568 217212 142624
rect 214741 142566 217212 142568
rect 214741 142563 214807 142566
rect 307661 142490 307727 142493
rect 324589 142490 324655 142493
rect 307661 142488 310132 142490
rect 307661 142432 307666 142488
rect 307722 142432 310132 142488
rect 307661 142430 310132 142432
rect 321908 142488 324655 142490
rect 321908 142432 324594 142488
rect 324650 142432 324655 142488
rect 321908 142430 324655 142432
rect 307661 142427 307727 142430
rect 324589 142427 324655 142430
rect 306005 142354 306071 142357
rect 306557 142354 306623 142357
rect 306005 142352 306623 142354
rect 306005 142296 306010 142352
rect 306066 142296 306562 142352
rect 306618 142296 306623 142352
rect 306005 142294 306623 142296
rect 306005 142291 306071 142294
rect 306557 142291 306623 142294
rect 259678 142218 259684 142220
rect 248860 142158 259684 142218
rect 259678 142156 259684 142158
rect 259748 142156 259754 142220
rect 306925 142082 306991 142085
rect 306925 142080 310132 142082
rect 306925 142024 306930 142080
rect 306986 142024 310132 142080
rect 306925 142022 310132 142024
rect 306925 142019 306991 142022
rect 213913 141946 213979 141949
rect 213913 141944 217212 141946
rect 213913 141888 213918 141944
rect 213974 141888 217212 141944
rect 213913 141886 217212 141888
rect 213913 141883 213979 141886
rect 248860 141750 253306 141810
rect 249977 141402 250043 141405
rect 248860 141400 250043 141402
rect 248860 141344 249982 141400
rect 250038 141344 250043 141400
rect 248860 141342 250043 141344
rect 249977 141339 250043 141342
rect 214005 141266 214071 141269
rect 253246 141266 253306 141750
rect 307293 141674 307359 141677
rect 324313 141674 324379 141677
rect 307293 141672 310132 141674
rect 307293 141616 307298 141672
rect 307354 141616 310132 141672
rect 307293 141614 310132 141616
rect 321908 141672 324379 141674
rect 321908 141616 324318 141672
rect 324374 141616 324379 141672
rect 321908 141614 324379 141616
rect 307293 141611 307359 141614
rect 324313 141611 324379 141614
rect 253422 141340 253428 141404
rect 253492 141402 253498 141404
rect 306557 141402 306623 141405
rect 253492 141400 306623 141402
rect 253492 141344 306562 141400
rect 306618 141344 306623 141400
rect 253492 141342 306623 141344
rect 253492 141340 253498 141342
rect 306557 141339 306623 141342
rect 260966 141266 260972 141268
rect 214005 141264 217212 141266
rect 214005 141208 214010 141264
rect 214066 141208 217212 141264
rect 214005 141206 217212 141208
rect 253246 141206 260972 141266
rect 214005 141203 214071 141206
rect 260966 141204 260972 141206
rect 261036 141204 261042 141268
rect 307385 141266 307451 141269
rect 307385 141264 310132 141266
rect 307385 141208 307390 141264
rect 307446 141208 310132 141264
rect 307385 141206 310132 141208
rect 307385 141203 307451 141206
rect 251214 140858 251220 140860
rect 248860 140798 251220 140858
rect 251214 140796 251220 140798
rect 251284 140796 251290 140860
rect 306097 140858 306163 140861
rect 324589 140858 324655 140861
rect 306097 140856 310132 140858
rect 306097 140800 306102 140856
rect 306158 140800 310132 140856
rect 306097 140798 310132 140800
rect 321908 140856 324655 140858
rect 321908 140800 324594 140856
rect 324650 140800 324655 140856
rect 321908 140798 324655 140800
rect 306097 140795 306163 140798
rect 324589 140795 324655 140798
rect 213913 140586 213979 140589
rect 213913 140584 217212 140586
rect 213913 140528 213918 140584
rect 213974 140528 217212 140584
rect 213913 140526 217212 140528
rect 213913 140523 213979 140526
rect 252093 140450 252159 140453
rect 248860 140448 252159 140450
rect 248860 140392 252098 140448
rect 252154 140392 252159 140448
rect 248860 140390 252159 140392
rect 252093 140387 252159 140390
rect 307477 140450 307543 140453
rect 307477 140448 310132 140450
rect 307477 140392 307482 140448
rect 307538 140392 310132 140448
rect 307477 140390 310132 140392
rect 307477 140387 307543 140390
rect 324313 140178 324379 140181
rect 321908 140176 324379 140178
rect 321908 140120 324318 140176
rect 324374 140120 324379 140176
rect 321908 140118 324379 140120
rect 324313 140115 324379 140118
rect 307569 140042 307635 140045
rect 307569 140040 310132 140042
rect 307569 139984 307574 140040
rect 307630 139984 310132 140040
rect 307569 139982 310132 139984
rect 307569 139979 307635 139982
rect 213177 139906 213243 139909
rect 213177 139904 217212 139906
rect 213177 139848 213182 139904
rect 213238 139848 217212 139904
rect 213177 139846 217212 139848
rect 248860 139846 258090 139906
rect 213177 139843 213243 139846
rect 258030 139770 258090 139846
rect 270534 139770 270540 139772
rect 258030 139710 270540 139770
rect 270534 139708 270540 139710
rect 270604 139708 270610 139772
rect 307661 139634 307727 139637
rect 307661 139632 310132 139634
rect 307661 139576 307666 139632
rect 307722 139576 310132 139632
rect 307661 139574 310132 139576
rect 307661 139571 307727 139574
rect 255262 139498 255268 139500
rect 248860 139438 255268 139498
rect 255262 139436 255268 139438
rect 255332 139436 255338 139500
rect 324313 139362 324379 139365
rect 321908 139360 324379 139362
rect 321908 139304 324318 139360
rect 324374 139304 324379 139360
rect 321908 139302 324379 139304
rect 324313 139299 324379 139302
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 214005 139226 214071 139229
rect 214005 139224 217212 139226
rect 214005 139168 214010 139224
rect 214066 139168 217212 139224
rect 583520 139212 584960 139302
rect 214005 139166 217212 139168
rect 214005 139163 214071 139166
rect 307477 139090 307543 139093
rect 307477 139088 310132 139090
rect 307477 139032 307482 139088
rect 307538 139032 310132 139088
rect 307477 139030 310132 139032
rect 307477 139027 307543 139030
rect 248860 138894 253306 138954
rect 213913 138682 213979 138685
rect 213913 138680 217212 138682
rect 213913 138624 213918 138680
rect 213974 138624 217212 138680
rect 213913 138622 217212 138624
rect 213913 138619 213979 138622
rect 249793 138546 249859 138549
rect 248860 138544 249859 138546
rect 248860 138488 249798 138544
rect 249854 138488 249859 138544
rect 248860 138486 249859 138488
rect 253246 138546 253306 138894
rect 256693 138682 256759 138685
rect 273846 138682 273852 138684
rect 256693 138680 273852 138682
rect 256693 138624 256698 138680
rect 256754 138624 273852 138680
rect 256693 138622 273852 138624
rect 256693 138619 256759 138622
rect 273846 138620 273852 138622
rect 273916 138620 273922 138684
rect 307569 138682 307635 138685
rect 307569 138680 310132 138682
rect 307569 138624 307574 138680
rect 307630 138624 310132 138680
rect 307569 138622 310132 138624
rect 307569 138619 307635 138622
rect 259494 138546 259500 138548
rect 253246 138486 259500 138546
rect 249793 138483 249859 138486
rect 259494 138484 259500 138486
rect 259564 138484 259570 138548
rect 307661 138274 307727 138277
rect 307661 138272 310132 138274
rect 307661 138216 307666 138272
rect 307722 138216 310132 138272
rect 307661 138214 310132 138216
rect 307661 138211 307727 138214
rect 321878 138138 321938 138516
rect 334014 138138 334020 138140
rect 321878 138078 334020 138138
rect 334014 138076 334020 138078
rect 334084 138076 334090 138140
rect 214649 138002 214715 138005
rect 252461 138002 252527 138005
rect 214649 138000 217212 138002
rect 214649 137944 214654 138000
rect 214710 137944 217212 138000
rect 214649 137942 217212 137944
rect 248860 138000 252527 138002
rect 248860 137944 252466 138000
rect 252522 137944 252527 138000
rect 248860 137942 252527 137944
rect 214649 137939 214715 137942
rect 252461 137939 252527 137942
rect 307569 137866 307635 137869
rect 324313 137866 324379 137869
rect 307569 137864 310132 137866
rect 307569 137808 307574 137864
rect 307630 137808 310132 137864
rect 307569 137806 310132 137808
rect 321908 137864 324379 137866
rect 321908 137808 324318 137864
rect 324374 137808 324379 137864
rect 321908 137806 324379 137808
rect 307569 137803 307635 137806
rect 324313 137803 324379 137806
rect 252093 137594 252159 137597
rect 248860 137592 252159 137594
rect 248860 137536 252098 137592
rect 252154 137536 252159 137592
rect 248860 137534 252159 137536
rect 252093 137531 252159 137534
rect 306557 137458 306623 137461
rect 306557 137456 310132 137458
rect 306557 137400 306562 137456
rect 306618 137400 310132 137456
rect 306557 137398 310132 137400
rect 306557 137395 306623 137398
rect 213913 137322 213979 137325
rect 213913 137320 217212 137322
rect 213913 137264 213918 137320
rect 213974 137264 217212 137320
rect 213913 137262 217212 137264
rect 213913 137259 213979 137262
rect 252369 137050 252435 137053
rect 248860 137048 252435 137050
rect 248860 136992 252374 137048
rect 252430 136992 252435 137048
rect 248860 136990 252435 136992
rect 252369 136987 252435 136990
rect 307661 137050 307727 137053
rect 324405 137050 324471 137053
rect 307661 137048 310132 137050
rect 307661 136992 307666 137048
rect 307722 136992 310132 137048
rect 307661 136990 310132 136992
rect 321908 137048 324471 137050
rect 321908 136992 324410 137048
rect 324466 136992 324471 137048
rect 321908 136990 324471 136992
rect 307661 136987 307727 136990
rect 324405 136987 324471 136990
rect 214557 136642 214623 136645
rect 250529 136642 250595 136645
rect 214557 136640 217212 136642
rect 214557 136584 214562 136640
rect 214618 136584 217212 136640
rect 214557 136582 217212 136584
rect 248860 136640 250595 136642
rect 248860 136584 250534 136640
rect 250590 136584 250595 136640
rect 248860 136582 250595 136584
rect 214557 136579 214623 136582
rect 250529 136579 250595 136582
rect 307477 136642 307543 136645
rect 307477 136640 310132 136642
rect 307477 136584 307482 136640
rect 307538 136584 310132 136640
rect 307477 136582 310132 136584
rect 307477 136579 307543 136582
rect 324313 136370 324379 136373
rect 321908 136368 324379 136370
rect 321908 136312 324318 136368
rect 324374 136312 324379 136368
rect 321908 136310 324379 136312
rect 324313 136307 324379 136310
rect 252093 136234 252159 136237
rect 248860 136232 252159 136234
rect 248860 136176 252098 136232
rect 252154 136176 252159 136232
rect 248860 136174 252159 136176
rect 252093 136171 252159 136174
rect 307569 136234 307635 136237
rect 307569 136232 310132 136234
rect 307569 136176 307574 136232
rect 307630 136176 310132 136232
rect 307569 136174 310132 136176
rect 307569 136171 307635 136174
rect 214005 135962 214071 135965
rect 214005 135960 217212 135962
rect 214005 135904 214010 135960
rect 214066 135904 217212 135960
rect 214005 135902 217212 135904
rect 214005 135899 214071 135902
rect 252369 135690 252435 135693
rect 248860 135688 252435 135690
rect 248860 135632 252374 135688
rect 252430 135632 252435 135688
rect 248860 135630 252435 135632
rect 252369 135627 252435 135630
rect 307661 135690 307727 135693
rect 307661 135688 310132 135690
rect 307661 135632 307666 135688
rect 307722 135632 310132 135688
rect 307661 135630 310132 135632
rect 307661 135627 307727 135630
rect 324405 135554 324471 135557
rect 321908 135552 324471 135554
rect 321908 135496 324410 135552
rect 324466 135496 324471 135552
rect 321908 135494 324471 135496
rect 324405 135491 324471 135494
rect 213913 135282 213979 135285
rect 252461 135282 252527 135285
rect 213913 135280 217212 135282
rect 213913 135224 213918 135280
rect 213974 135224 217212 135280
rect 213913 135222 217212 135224
rect 248860 135280 252527 135282
rect 248860 135224 252466 135280
rect 252522 135224 252527 135280
rect 248860 135222 252527 135224
rect 213913 135219 213979 135222
rect 252461 135219 252527 135222
rect 307661 135282 307727 135285
rect 307661 135280 310132 135282
rect 307661 135224 307666 135280
rect 307722 135224 310132 135280
rect 307661 135222 310132 135224
rect 307661 135219 307727 135222
rect 307477 134874 307543 134877
rect 307477 134872 310132 134874
rect 307477 134816 307482 134872
rect 307538 134816 310132 134872
rect 307477 134814 310132 134816
rect 307477 134811 307543 134814
rect 251633 134738 251699 134741
rect 248860 134736 251699 134738
rect 248860 134680 251638 134736
rect 251694 134680 251699 134736
rect 248860 134678 251699 134680
rect 251633 134675 251699 134678
rect 167494 134132 167500 134196
rect 167564 134194 167570 134196
rect 217182 134194 217242 134572
rect 307661 134466 307727 134469
rect 307661 134464 310132 134466
rect 307661 134408 307666 134464
rect 307722 134408 310132 134464
rect 307661 134406 310132 134408
rect 307661 134403 307727 134406
rect 252461 134330 252527 134333
rect 248860 134328 252527 134330
rect 248860 134272 252466 134328
rect 252522 134272 252527 134328
rect 248860 134270 252527 134272
rect 252461 134267 252527 134270
rect 167564 134134 217242 134194
rect 321878 134194 321938 134708
rect 331438 134194 331444 134196
rect 321878 134134 331444 134194
rect 167564 134132 167570 134134
rect 331438 134132 331444 134134
rect 331508 134132 331514 134196
rect 307569 134058 307635 134061
rect 307569 134056 310132 134058
rect 307569 134000 307574 134056
rect 307630 134000 310132 134056
rect 307569 133998 310132 134000
rect 321908 133998 325710 134058
rect 307569 133995 307635 133998
rect 213913 133922 213979 133925
rect 325650 133922 325710 133998
rect 332726 133922 332732 133924
rect 213913 133920 217212 133922
rect 213913 133864 213918 133920
rect 213974 133864 217212 133920
rect 213913 133862 217212 133864
rect 325650 133862 332732 133922
rect 213913 133859 213979 133862
rect 332726 133860 332732 133862
rect 332796 133860 332802 133924
rect 252461 133786 252527 133789
rect 248860 133784 252527 133786
rect 248860 133728 252466 133784
rect 252522 133728 252527 133784
rect 248860 133726 252527 133728
rect 252461 133723 252527 133726
rect 307385 133650 307451 133653
rect 307385 133648 310132 133650
rect 307385 133592 307390 133648
rect 307446 133592 310132 133648
rect 307385 133590 310132 133592
rect 307385 133587 307451 133590
rect 213913 133378 213979 133381
rect 251449 133378 251515 133381
rect 213913 133376 217212 133378
rect 213913 133320 213918 133376
rect 213974 133320 217212 133376
rect 213913 133318 217212 133320
rect 248860 133376 251515 133378
rect 248860 133320 251454 133376
rect 251510 133320 251515 133376
rect 248860 133318 251515 133320
rect 213913 133315 213979 133318
rect 251449 133315 251515 133318
rect 307569 133242 307635 133245
rect 324497 133242 324563 133245
rect 307569 133240 310132 133242
rect 307569 133184 307574 133240
rect 307630 133184 310132 133240
rect 307569 133182 310132 133184
rect 321908 133240 324563 133242
rect 321908 133184 324502 133240
rect 324558 133184 324563 133240
rect 321908 133182 324563 133184
rect 307569 133179 307635 133182
rect 324497 133179 324563 133182
rect 252001 132834 252067 132837
rect 248860 132832 252067 132834
rect 248860 132776 252006 132832
rect 252062 132776 252067 132832
rect 248860 132774 252067 132776
rect 252001 132771 252067 132774
rect 307661 132698 307727 132701
rect 321553 132698 321619 132701
rect 200070 132638 217212 132698
rect 307661 132696 310132 132698
rect 307661 132640 307666 132696
rect 307722 132640 310132 132696
rect 307661 132638 310132 132640
rect 321510 132696 321619 132698
rect 321510 132640 321558 132696
rect 321614 132640 321619 132696
rect 166390 132500 166396 132564
rect 166460 132562 166466 132564
rect 200070 132562 200130 132638
rect 307661 132635 307727 132638
rect 321510 132635 321619 132640
rect 166460 132502 200130 132562
rect 166460 132500 166466 132502
rect 252461 132426 252527 132429
rect 248860 132424 252527 132426
rect 248860 132368 252466 132424
rect 252522 132368 252527 132424
rect 321510 132396 321570 132635
rect 248860 132366 252527 132368
rect 252461 132363 252527 132366
rect 307661 132290 307727 132293
rect 307661 132288 310132 132290
rect 307661 132232 307666 132288
rect 307722 132232 310132 132288
rect 307661 132230 310132 132232
rect 307661 132227 307727 132230
rect 169150 131412 169156 131476
rect 169220 131474 169226 131476
rect 217182 131474 217242 131988
rect 251541 131882 251607 131885
rect 248860 131880 251607 131882
rect 248860 131824 251546 131880
rect 251602 131824 251607 131880
rect 248860 131822 251607 131824
rect 251541 131819 251607 131822
rect 307017 131882 307083 131885
rect 307017 131880 310132 131882
rect 307017 131824 307022 131880
rect 307078 131824 310132 131880
rect 307017 131822 310132 131824
rect 307017 131819 307083 131822
rect 251766 131684 251772 131748
rect 251836 131746 251842 131748
rect 305637 131746 305703 131749
rect 324313 131746 324379 131749
rect 251836 131744 305703 131746
rect 251836 131688 305642 131744
rect 305698 131688 305703 131744
rect 251836 131686 305703 131688
rect 321908 131744 324379 131746
rect 321908 131688 324318 131744
rect 324374 131688 324379 131744
rect 321908 131686 324379 131688
rect 251836 131684 251842 131686
rect 305637 131683 305703 131686
rect 324313 131683 324379 131686
rect 252277 131474 252343 131477
rect 169220 131414 217242 131474
rect 248860 131472 252343 131474
rect 248860 131416 252282 131472
rect 252338 131416 252343 131472
rect 248860 131414 252343 131416
rect 169220 131412 169226 131414
rect 252277 131411 252343 131414
rect 295926 131412 295932 131476
rect 295996 131474 296002 131476
rect 295996 131414 310132 131474
rect 295996 131412 296002 131414
rect 213913 131338 213979 131341
rect 213913 131336 217212 131338
rect 213913 131280 213918 131336
rect 213974 131280 217212 131336
rect 213913 131278 217212 131280
rect 213913 131275 213979 131278
rect 306741 131066 306807 131069
rect 306741 131064 310132 131066
rect 306741 131008 306746 131064
rect 306802 131008 310132 131064
rect 306741 131006 310132 131008
rect 306741 131003 306807 131006
rect 251541 130930 251607 130933
rect 324313 130930 324379 130933
rect 248860 130928 251607 130930
rect 248860 130872 251546 130928
rect 251602 130872 251607 130928
rect 248860 130870 251607 130872
rect 321908 130928 324379 130930
rect 321908 130872 324318 130928
rect 324374 130872 324379 130928
rect 321908 130870 324379 130872
rect 251541 130867 251607 130870
rect 324313 130867 324379 130870
rect 214925 130658 214991 130661
rect 214925 130656 217212 130658
rect 214925 130600 214930 130656
rect 214986 130600 217212 130656
rect 214925 130598 217212 130600
rect 214925 130595 214991 130598
rect 307150 130596 307156 130660
rect 307220 130658 307226 130660
rect 307220 130598 310132 130658
rect 307220 130596 307226 130598
rect 252461 130522 252527 130525
rect 248860 130520 252527 130522
rect 248860 130464 252466 130520
rect 252522 130464 252527 130520
rect 248860 130462 252527 130464
rect 252461 130459 252527 130462
rect 307569 130250 307635 130253
rect 307569 130248 310132 130250
rect 307569 130192 307574 130248
rect 307630 130192 310132 130248
rect 307569 130190 310132 130192
rect 307569 130187 307635 130190
rect 251817 130114 251883 130117
rect 324405 130114 324471 130117
rect 248860 130112 251883 130114
rect 248860 130056 251822 130112
rect 251878 130056 251883 130112
rect 248860 130054 251883 130056
rect 321908 130112 324471 130114
rect 321908 130056 324410 130112
rect 324466 130056 324471 130112
rect 321908 130054 324471 130056
rect 251817 130051 251883 130054
rect 324405 130051 324471 130054
rect 213913 129978 213979 129981
rect 213913 129976 217212 129978
rect 213913 129920 213918 129976
rect 213974 129920 217212 129976
rect 213913 129918 217212 129920
rect 213913 129915 213979 129918
rect 307661 129842 307727 129845
rect 307661 129840 310132 129842
rect 307661 129784 307666 129840
rect 307722 129784 310132 129840
rect 307661 129782 310132 129784
rect 307661 129779 307727 129782
rect 252461 129570 252527 129573
rect 248860 129568 252527 129570
rect 248860 129512 252466 129568
rect 252522 129512 252527 129568
rect 248860 129510 252527 129512
rect 252461 129507 252527 129510
rect 324313 129434 324379 129437
rect 321908 129432 324379 129434
rect 321908 129376 324318 129432
rect 324374 129376 324379 129432
rect 321908 129374 324379 129376
rect 324313 129371 324379 129374
rect 66069 129298 66135 129301
rect 68142 129298 68816 129304
rect 66069 129296 68816 129298
rect 66069 129240 66074 129296
rect 66130 129244 68816 129296
rect 66130 129240 68202 129244
rect 66069 129238 68202 129240
rect 66069 129235 66135 129238
rect 213913 129298 213979 129301
rect 307385 129298 307451 129301
rect 213913 129296 217212 129298
rect 213913 129240 213918 129296
rect 213974 129240 217212 129296
rect 213913 129238 217212 129240
rect 307385 129296 310132 129298
rect 307385 129240 307390 129296
rect 307446 129240 310132 129296
rect 307385 129238 310132 129240
rect 213913 129235 213979 129238
rect 307385 129235 307451 129238
rect 251725 129162 251791 129165
rect 248860 129160 251791 129162
rect 248860 129104 251730 129160
rect 251786 129104 251791 129160
rect 248860 129102 251791 129104
rect 251725 129099 251791 129102
rect 307661 128890 307727 128893
rect 307661 128888 310132 128890
rect 307661 128832 307666 128888
rect 307722 128832 310132 128888
rect 307661 128830 310132 128832
rect 307661 128827 307727 128830
rect 200070 128694 217212 128754
rect 166206 128556 166212 128620
rect 166276 128618 166282 128620
rect 200070 128618 200130 128694
rect 252001 128618 252067 128621
rect 324405 128618 324471 128621
rect 166276 128558 200130 128618
rect 248860 128616 252067 128618
rect 248860 128560 252006 128616
rect 252062 128560 252067 128616
rect 248860 128558 252067 128560
rect 321908 128616 324471 128618
rect 321908 128560 324410 128616
rect 324466 128560 324471 128616
rect 321908 128558 324471 128560
rect 166276 128556 166282 128558
rect 252001 128555 252067 128558
rect 324405 128555 324471 128558
rect 307569 128482 307635 128485
rect 307569 128480 310132 128482
rect 307569 128424 307574 128480
rect 307630 128424 310132 128480
rect 307569 128422 310132 128424
rect 307569 128419 307635 128422
rect 252461 128210 252527 128213
rect 248860 128208 252527 128210
rect 248860 128152 252466 128208
rect 252522 128152 252527 128208
rect 248860 128150 252527 128152
rect 252461 128147 252527 128150
rect 67633 128074 67699 128077
rect 68142 128074 68816 128080
rect 67633 128072 68816 128074
rect 67633 128016 67638 128072
rect 67694 128020 68816 128072
rect 67694 128016 68202 128020
rect 67633 128014 68202 128016
rect 67633 128011 67699 128014
rect 214005 128074 214071 128077
rect 307661 128074 307727 128077
rect 214005 128072 217212 128074
rect 214005 128016 214010 128072
rect 214066 128016 217212 128072
rect 214005 128014 217212 128016
rect 307661 128072 310132 128074
rect 307661 128016 307666 128072
rect 307722 128016 310132 128072
rect 307661 128014 310132 128016
rect 214005 128011 214071 128014
rect 307661 128011 307727 128014
rect 324313 127802 324379 127805
rect 321908 127800 324379 127802
rect 321908 127744 324318 127800
rect 324374 127744 324379 127800
rect 321908 127742 324379 127744
rect 324313 127739 324379 127742
rect 252369 127666 252435 127669
rect 248860 127664 252435 127666
rect 248860 127608 252374 127664
rect 252430 127608 252435 127664
rect 248860 127606 252435 127608
rect 252369 127603 252435 127606
rect 307109 127666 307175 127669
rect 307109 127664 310132 127666
rect 307109 127608 307114 127664
rect 307170 127608 310132 127664
rect 307109 127606 310132 127608
rect 307109 127603 307175 127606
rect 213913 127394 213979 127397
rect 213913 127392 217212 127394
rect 213913 127336 213918 127392
rect 213974 127336 217212 127392
rect 213913 127334 217212 127336
rect 213913 127331 213979 127334
rect 252001 127258 252067 127261
rect 248860 127256 252067 127258
rect 248860 127200 252006 127256
rect 252062 127200 252067 127256
rect 248860 127198 252067 127200
rect 252001 127195 252067 127198
rect 306741 127258 306807 127261
rect 306741 127256 310132 127258
rect 306741 127200 306746 127256
rect 306802 127200 310132 127256
rect 306741 127198 310132 127200
rect 306741 127195 306807 127198
rect 324405 127122 324471 127125
rect 321908 127120 324471 127122
rect 321908 127064 324410 127120
rect 324466 127064 324471 127120
rect 321908 127062 324471 127064
rect 324405 127059 324471 127062
rect 306741 126850 306807 126853
rect 306741 126848 310132 126850
rect 306741 126792 306746 126848
rect 306802 126792 310132 126848
rect 306741 126790 310132 126792
rect 306741 126787 306807 126790
rect 213913 126714 213979 126717
rect 252461 126714 252527 126717
rect 213913 126712 217212 126714
rect 213913 126656 213918 126712
rect 213974 126656 217212 126712
rect 213913 126654 217212 126656
rect 248860 126712 252527 126714
rect 248860 126656 252466 126712
rect 252522 126656 252527 126712
rect 248860 126654 252527 126656
rect 213913 126651 213979 126654
rect 252461 126651 252527 126654
rect 300158 126380 300164 126444
rect 300228 126442 300234 126444
rect 300228 126382 310132 126442
rect 300228 126380 300234 126382
rect 66161 126306 66227 126309
rect 68142 126306 68816 126312
rect 66161 126304 68816 126306
rect 66161 126248 66166 126304
rect 66222 126252 68816 126304
rect 251909 126306 251975 126309
rect 66222 126248 68202 126252
rect 66161 126246 68202 126248
rect 66161 126243 66227 126246
rect 248860 126304 251975 126306
rect 248860 126248 251914 126304
rect 251970 126248 251975 126304
rect 248860 126246 251975 126248
rect 251909 126243 251975 126246
rect 214465 126034 214531 126037
rect 214465 126032 217212 126034
rect 214465 125976 214470 126032
rect 214526 125976 217212 126032
rect 214465 125974 217212 125976
rect 214465 125971 214531 125974
rect 307661 125898 307727 125901
rect 307661 125896 310132 125898
rect 307661 125840 307666 125896
rect 307722 125840 310132 125896
rect 307661 125838 310132 125840
rect 307661 125835 307727 125838
rect 252185 125762 252251 125765
rect 248860 125760 252251 125762
rect 248860 125704 252190 125760
rect 252246 125704 252251 125760
rect 248860 125702 252251 125704
rect 252185 125699 252251 125702
rect 321878 125626 321938 126276
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect 328494 125626 328500 125628
rect 321878 125566 328500 125626
rect 328494 125564 328500 125566
rect 328564 125564 328570 125628
rect 307569 125490 307635 125493
rect 325785 125490 325851 125493
rect 307569 125488 310132 125490
rect 307569 125432 307574 125488
rect 307630 125432 310132 125488
rect 307569 125430 310132 125432
rect 321908 125488 325851 125490
rect 321908 125432 325790 125488
rect 325846 125432 325851 125488
rect 321908 125430 325851 125432
rect 307569 125427 307635 125430
rect 325785 125427 325851 125430
rect 214005 125354 214071 125357
rect 251173 125354 251239 125357
rect 214005 125352 217212 125354
rect 214005 125296 214010 125352
rect 214066 125296 217212 125352
rect 214005 125294 217212 125296
rect 248860 125352 251239 125354
rect 248860 125296 251178 125352
rect 251234 125296 251239 125352
rect 248860 125294 251239 125296
rect 214005 125291 214071 125294
rect 251173 125291 251239 125294
rect 65517 125218 65583 125221
rect 68142 125218 68816 125224
rect 65517 125216 68816 125218
rect 65517 125160 65522 125216
rect 65578 125164 68816 125216
rect 65578 125160 68202 125164
rect 65517 125158 68202 125160
rect 65517 125155 65583 125158
rect -960 123572 480 123812
rect 306741 125082 306807 125085
rect 306741 125080 310132 125082
rect 306741 125024 306746 125080
rect 306802 125024 310132 125080
rect 306741 125022 310132 125024
rect 306741 125019 306807 125022
rect 251265 124810 251331 124813
rect 324313 124810 324379 124813
rect 248860 124808 251331 124810
rect 248860 124752 251270 124808
rect 251326 124752 251331 124808
rect 248860 124750 251331 124752
rect 321908 124808 324379 124810
rect 321908 124752 324318 124808
rect 324374 124752 324379 124808
rect 321908 124750 324379 124752
rect 251265 124747 251331 124750
rect 324313 124747 324379 124750
rect 213913 124674 213979 124677
rect 307661 124674 307727 124677
rect 213913 124672 217212 124674
rect 213913 124616 213918 124672
rect 213974 124616 217212 124672
rect 213913 124614 217212 124616
rect 307661 124672 310132 124674
rect 307661 124616 307666 124672
rect 307722 124616 310132 124672
rect 307661 124614 310132 124616
rect 213913 124611 213979 124614
rect 307661 124611 307727 124614
rect 252185 124402 252251 124405
rect 248860 124400 252251 124402
rect 248860 124344 252190 124400
rect 252246 124344 252251 124400
rect 248860 124342 252251 124344
rect 252185 124339 252251 124342
rect 307109 124266 307175 124269
rect 307109 124264 310132 124266
rect 307109 124208 307114 124264
rect 307170 124208 310132 124264
rect 307109 124206 310132 124208
rect 307109 124203 307175 124206
rect 214005 124130 214071 124133
rect 214005 124128 217212 124130
rect 214005 124072 214010 124128
rect 214066 124072 217212 124128
rect 214005 124070 217212 124072
rect 214005 124067 214071 124070
rect 252461 123994 252527 123997
rect 248860 123992 252527 123994
rect 248860 123936 252466 123992
rect 252522 123936 252527 123992
rect 248860 123934 252527 123936
rect 252461 123931 252527 123934
rect 306557 123858 306623 123861
rect 306557 123856 310132 123858
rect 306557 123800 306562 123856
rect 306618 123800 310132 123856
rect 306557 123798 310132 123800
rect 306557 123795 306623 123798
rect 66069 123586 66135 123589
rect 68142 123586 68816 123592
rect 66069 123584 68816 123586
rect 66069 123528 66074 123584
rect 66130 123532 68816 123584
rect 66130 123528 68202 123532
rect 66069 123526 68202 123528
rect 66069 123523 66135 123526
rect 213913 123450 213979 123453
rect 252093 123450 252159 123453
rect 213913 123448 217212 123450
rect 213913 123392 213918 123448
rect 213974 123392 217212 123448
rect 213913 123390 217212 123392
rect 248860 123448 252159 123450
rect 248860 123392 252098 123448
rect 252154 123392 252159 123448
rect 248860 123390 252159 123392
rect 213913 123387 213979 123390
rect 252093 123387 252159 123390
rect 307569 123450 307635 123453
rect 307569 123448 310132 123450
rect 307569 123392 307574 123448
rect 307630 123392 310132 123448
rect 307569 123390 310132 123392
rect 307569 123387 307635 123390
rect 321878 123314 321938 123964
rect 329782 123314 329788 123316
rect 321878 123254 329788 123314
rect 329782 123252 329788 123254
rect 329852 123252 329858 123316
rect 324313 123178 324379 123181
rect 321908 123176 324379 123178
rect 321908 123120 324318 123176
rect 324374 123120 324379 123176
rect 321908 123118 324379 123120
rect 324313 123115 324379 123118
rect 251725 123042 251791 123045
rect 248860 123040 251791 123042
rect 248860 122984 251730 123040
rect 251786 122984 251791 123040
rect 248860 122982 251791 122984
rect 251725 122979 251791 122982
rect 307661 123042 307727 123045
rect 307661 123040 310132 123042
rect 307661 122984 307666 123040
rect 307722 122984 310132 123040
rect 307661 122982 310132 122984
rect 307661 122979 307727 122982
rect 214005 122770 214071 122773
rect 214005 122768 217212 122770
rect 214005 122712 214010 122768
rect 214066 122712 217212 122768
rect 214005 122710 217212 122712
rect 214005 122707 214071 122710
rect 66069 122634 66135 122637
rect 68142 122634 68816 122640
rect 66069 122632 68816 122634
rect 66069 122576 66074 122632
rect 66130 122580 68816 122632
rect 66130 122576 68202 122580
rect 66069 122574 68202 122576
rect 66069 122571 66135 122574
rect 252461 122498 252527 122501
rect 248860 122496 252527 122498
rect 248860 122440 252466 122496
rect 252522 122440 252527 122496
rect 248860 122438 252527 122440
rect 252461 122435 252527 122438
rect 306741 122498 306807 122501
rect 324313 122498 324379 122501
rect 306741 122496 310132 122498
rect 306741 122440 306746 122496
rect 306802 122440 310132 122496
rect 306741 122438 310132 122440
rect 321908 122496 324379 122498
rect 321908 122440 324318 122496
rect 324374 122440 324379 122496
rect 321908 122438 324379 122440
rect 306741 122435 306807 122438
rect 324313 122435 324379 122438
rect 213913 122090 213979 122093
rect 252369 122090 252435 122093
rect 213913 122088 217212 122090
rect 213913 122032 213918 122088
rect 213974 122032 217212 122088
rect 213913 122030 217212 122032
rect 248860 122088 252435 122090
rect 248860 122032 252374 122088
rect 252430 122032 252435 122088
rect 248860 122030 252435 122032
rect 213913 122027 213979 122030
rect 252369 122027 252435 122030
rect 307569 122090 307635 122093
rect 307569 122088 310132 122090
rect 307569 122032 307574 122088
rect 307630 122032 310132 122088
rect 307569 122030 310132 122032
rect 307569 122027 307635 122030
rect 307661 121682 307727 121685
rect 327022 121682 327028 121684
rect 307661 121680 310132 121682
rect 307661 121624 307666 121680
rect 307722 121624 310132 121680
rect 307661 121622 310132 121624
rect 321908 121622 327028 121682
rect 307661 121619 307727 121622
rect 327022 121620 327028 121622
rect 327092 121620 327098 121684
rect 252461 121546 252527 121549
rect 248860 121544 252527 121546
rect 248860 121488 252466 121544
rect 252522 121488 252527 121544
rect 248860 121486 252527 121488
rect 252461 121483 252527 121486
rect 214005 121410 214071 121413
rect 214005 121408 217212 121410
rect 214005 121352 214010 121408
rect 214066 121352 217212 121408
rect 214005 121350 217212 121352
rect 214005 121347 214071 121350
rect 306741 121274 306807 121277
rect 306741 121272 310132 121274
rect 306741 121216 306746 121272
rect 306802 121216 310132 121272
rect 306741 121214 310132 121216
rect 306741 121211 306807 121214
rect 252461 121138 252527 121141
rect 248860 121136 252527 121138
rect 248860 121080 252466 121136
rect 252522 121080 252527 121136
rect 248860 121078 252527 121080
rect 252461 121075 252527 121078
rect 67449 120866 67515 120869
rect 68142 120866 68816 120872
rect 67449 120864 68816 120866
rect 67449 120808 67454 120864
rect 67510 120812 68816 120864
rect 67510 120808 68202 120812
rect 67449 120806 68202 120808
rect 67449 120803 67515 120806
rect 307569 120866 307635 120869
rect 324313 120866 324379 120869
rect 307569 120864 310132 120866
rect 307569 120808 307574 120864
rect 307630 120808 310132 120864
rect 307569 120806 310132 120808
rect 321908 120864 324379 120866
rect 321908 120808 324318 120864
rect 324374 120808 324379 120864
rect 321908 120806 324379 120808
rect 307569 120803 307635 120806
rect 324313 120803 324379 120806
rect 213913 120730 213979 120733
rect 213913 120728 217212 120730
rect 213913 120672 213918 120728
rect 213974 120672 217212 120728
rect 213913 120670 217212 120672
rect 213913 120667 213979 120670
rect 251909 120594 251975 120597
rect 248860 120592 251975 120594
rect 248860 120536 251914 120592
rect 251970 120536 251975 120592
rect 248860 120534 251975 120536
rect 251909 120531 251975 120534
rect 307661 120458 307727 120461
rect 307661 120456 310132 120458
rect 307661 120400 307666 120456
rect 307722 120400 310132 120456
rect 307661 120398 310132 120400
rect 307661 120395 307727 120398
rect 252093 120186 252159 120189
rect 324405 120186 324471 120189
rect 248860 120184 252159 120186
rect 248860 120128 252098 120184
rect 252154 120128 252159 120184
rect 248860 120126 252159 120128
rect 321908 120184 324471 120186
rect 321908 120128 324410 120184
rect 324466 120128 324471 120184
rect 321908 120126 324471 120128
rect 252093 120123 252159 120126
rect 324405 120123 324471 120126
rect 214097 120050 214163 120053
rect 307661 120050 307727 120053
rect 214097 120048 217212 120050
rect 214097 119992 214102 120048
rect 214158 119992 217212 120048
rect 214097 119990 217212 119992
rect 307661 120048 310132 120050
rect 307661 119992 307666 120048
rect 307722 119992 310132 120048
rect 307661 119990 310132 119992
rect 214097 119987 214163 119990
rect 307661 119987 307727 119990
rect 252461 119642 252527 119645
rect 248860 119640 252527 119642
rect 248860 119584 252466 119640
rect 252522 119584 252527 119640
rect 248860 119582 252527 119584
rect 252461 119579 252527 119582
rect 306741 119642 306807 119645
rect 306741 119640 310132 119642
rect 306741 119584 306746 119640
rect 306802 119584 310132 119640
rect 306741 119582 310132 119584
rect 306741 119579 306807 119582
rect 214005 119506 214071 119509
rect 214005 119504 217212 119506
rect 214005 119448 214010 119504
rect 214066 119448 217212 119504
rect 214005 119446 217212 119448
rect 214005 119443 214071 119446
rect 324313 119370 324379 119373
rect 321908 119368 324379 119370
rect 321908 119312 324318 119368
rect 324374 119312 324379 119368
rect 321908 119310 324379 119312
rect 324313 119307 324379 119310
rect 252369 119234 252435 119237
rect 248860 119232 252435 119234
rect 248860 119176 252374 119232
rect 252430 119176 252435 119232
rect 248860 119174 252435 119176
rect 252369 119171 252435 119174
rect 304206 119036 304212 119100
rect 304276 119098 304282 119100
rect 304276 119038 310132 119098
rect 304276 119036 304282 119038
rect 213913 118826 213979 118829
rect 251817 118826 251883 118829
rect 213913 118824 217212 118826
rect 213913 118768 213918 118824
rect 213974 118768 217212 118824
rect 213913 118766 217212 118768
rect 248860 118824 251883 118826
rect 248860 118768 251822 118824
rect 251878 118768 251883 118824
rect 248860 118766 251883 118768
rect 213913 118763 213979 118766
rect 251817 118763 251883 118766
rect 305494 118628 305500 118692
rect 305564 118690 305570 118692
rect 305564 118630 310132 118690
rect 305564 118628 305570 118630
rect 324313 118554 324379 118557
rect 321908 118552 324379 118554
rect 321908 118496 324318 118552
rect 324374 118496 324379 118552
rect 321908 118494 324379 118496
rect 324313 118491 324379 118494
rect 251541 118282 251607 118285
rect 248860 118280 251607 118282
rect 248860 118224 251546 118280
rect 251602 118224 251607 118280
rect 248860 118222 251607 118224
rect 251541 118219 251607 118222
rect 307477 118282 307543 118285
rect 307477 118280 310132 118282
rect 307477 118224 307482 118280
rect 307538 118224 310132 118280
rect 307477 118222 310132 118224
rect 307477 118219 307543 118222
rect 214005 118146 214071 118149
rect 214005 118144 217212 118146
rect 214005 118088 214010 118144
rect 214066 118088 217212 118144
rect 214005 118086 217212 118088
rect 214005 118083 214071 118086
rect 252461 117874 252527 117877
rect 248860 117872 252527 117874
rect 248860 117816 252466 117872
rect 252522 117816 252527 117872
rect 248860 117814 252527 117816
rect 252461 117811 252527 117814
rect 307661 117874 307727 117877
rect 324405 117874 324471 117877
rect 307661 117872 310132 117874
rect 307661 117816 307666 117872
rect 307722 117816 310132 117872
rect 307661 117814 310132 117816
rect 321908 117872 324471 117874
rect 321908 117816 324410 117872
rect 324466 117816 324471 117872
rect 321908 117814 324471 117816
rect 307661 117811 307727 117814
rect 324405 117811 324471 117814
rect 213913 117466 213979 117469
rect 213913 117464 217212 117466
rect 213913 117408 213918 117464
rect 213974 117408 217212 117464
rect 213913 117406 217212 117408
rect 213913 117403 213979 117406
rect 299974 117404 299980 117468
rect 300044 117466 300050 117468
rect 300044 117406 310132 117466
rect 300044 117404 300050 117406
rect 252093 117330 252159 117333
rect 248860 117328 252159 117330
rect 248860 117272 252098 117328
rect 252154 117272 252159 117328
rect 248860 117270 252159 117272
rect 252093 117267 252159 117270
rect 307661 117058 307727 117061
rect 324313 117058 324379 117061
rect 307661 117056 310132 117058
rect 307661 117000 307666 117056
rect 307722 117000 310132 117056
rect 307661 116998 310132 117000
rect 321908 117056 324379 117058
rect 321908 117000 324318 117056
rect 324374 117000 324379 117056
rect 321908 116998 324379 117000
rect 307661 116995 307727 116998
rect 324313 116995 324379 116998
rect 251541 116922 251607 116925
rect 248860 116920 251607 116922
rect 248860 116864 251546 116920
rect 251602 116864 251607 116920
rect 248860 116862 251607 116864
rect 251541 116859 251607 116862
rect 214005 116786 214071 116789
rect 214005 116784 217212 116786
rect 214005 116728 214010 116784
rect 214066 116728 217212 116784
rect 214005 116726 217212 116728
rect 214005 116723 214071 116726
rect 307477 116650 307543 116653
rect 307477 116648 310132 116650
rect 307477 116592 307482 116648
rect 307538 116592 310132 116648
rect 307477 116590 310132 116592
rect 307477 116587 307543 116590
rect 252369 116378 252435 116381
rect 324405 116378 324471 116381
rect 248860 116376 252435 116378
rect 248860 116320 252374 116376
rect 252430 116320 252435 116376
rect 248860 116318 252435 116320
rect 321908 116376 324471 116378
rect 321908 116320 324410 116376
rect 324466 116320 324471 116376
rect 321908 116318 324471 116320
rect 252369 116315 252435 116318
rect 324405 116315 324471 116318
rect 307017 116242 307083 116245
rect 307017 116240 310132 116242
rect 307017 116184 307022 116240
rect 307078 116184 310132 116240
rect 307017 116182 310132 116184
rect 307017 116179 307083 116182
rect 213913 116106 213979 116109
rect 213913 116104 217212 116106
rect 213913 116048 213918 116104
rect 213974 116048 217212 116104
rect 213913 116046 217212 116048
rect 213913 116043 213979 116046
rect 252277 115970 252343 115973
rect 248860 115968 252343 115970
rect 248860 115912 252282 115968
rect 252338 115912 252343 115968
rect 248860 115910 252343 115912
rect 252277 115907 252343 115910
rect 307477 115698 307543 115701
rect 307477 115696 310132 115698
rect 307477 115640 307482 115696
rect 307538 115640 310132 115696
rect 307477 115638 310132 115640
rect 307477 115635 307543 115638
rect 324313 115562 324379 115565
rect 321908 115560 324379 115562
rect 321908 115504 324318 115560
rect 324374 115504 324379 115560
rect 321908 115502 324379 115504
rect 324313 115499 324379 115502
rect 214005 115426 214071 115429
rect 251633 115426 251699 115429
rect 214005 115424 217212 115426
rect 214005 115368 214010 115424
rect 214066 115368 217212 115424
rect 214005 115366 217212 115368
rect 248860 115424 251699 115426
rect 248860 115368 251638 115424
rect 251694 115368 251699 115424
rect 248860 115366 251699 115368
rect 214005 115363 214071 115366
rect 251633 115363 251699 115366
rect 307569 115290 307635 115293
rect 307569 115288 310132 115290
rect 307569 115232 307574 115288
rect 307630 115232 310132 115288
rect 307569 115230 310132 115232
rect 307569 115227 307635 115230
rect 252369 115018 252435 115021
rect 248860 115016 252435 115018
rect 248860 114960 252374 115016
rect 252430 114960 252435 115016
rect 248860 114958 252435 114960
rect 252369 114955 252435 114958
rect 213913 114882 213979 114885
rect 307661 114882 307727 114885
rect 213913 114880 217212 114882
rect 213913 114824 213918 114880
rect 213974 114824 217212 114880
rect 213913 114822 217212 114824
rect 307661 114880 310132 114882
rect 307661 114824 307666 114880
rect 307722 114824 310132 114880
rect 307661 114822 310132 114824
rect 213913 114819 213979 114822
rect 307661 114819 307727 114822
rect 321908 114686 325710 114746
rect 325650 114610 325710 114686
rect 340822 114610 340828 114612
rect 325650 114550 340828 114610
rect 340822 114548 340828 114550
rect 340892 114548 340898 114612
rect 252461 114474 252527 114477
rect 248860 114472 252527 114474
rect 248860 114416 252466 114472
rect 252522 114416 252527 114472
rect 248860 114414 252527 114416
rect 252461 114411 252527 114414
rect 309133 114474 309199 114477
rect 309133 114472 310132 114474
rect 309133 114416 309138 114472
rect 309194 114416 310132 114472
rect 309133 114414 310132 114416
rect 309133 114411 309199 114414
rect 214005 114202 214071 114205
rect 214005 114200 217212 114202
rect 214005 114144 214010 114200
rect 214066 114144 217212 114200
rect 214005 114142 217212 114144
rect 214005 114139 214071 114142
rect 252461 114066 252527 114069
rect 248860 114064 252527 114066
rect 248860 114008 252466 114064
rect 252522 114008 252527 114064
rect 248860 114006 252527 114008
rect 252461 114003 252527 114006
rect 306966 114004 306972 114068
rect 307036 114066 307042 114068
rect 324313 114066 324379 114069
rect 307036 114006 310132 114066
rect 321908 114064 324379 114066
rect 321908 114008 324318 114064
rect 324374 114008 324379 114064
rect 321908 114006 324379 114008
rect 307036 114004 307042 114006
rect 324313 114003 324379 114006
rect 307661 113658 307727 113661
rect 307661 113656 310132 113658
rect 307661 113600 307666 113656
rect 307722 113600 310132 113656
rect 307661 113598 310132 113600
rect 307661 113595 307727 113598
rect 213913 113522 213979 113525
rect 252001 113522 252067 113525
rect 213913 113520 217212 113522
rect 213913 113464 213918 113520
rect 213974 113464 217212 113520
rect 213913 113462 217212 113464
rect 248860 113520 252067 113522
rect 248860 113464 252006 113520
rect 252062 113464 252067 113520
rect 248860 113462 252067 113464
rect 213913 113459 213979 113462
rect 252001 113459 252067 113462
rect 282126 113460 282132 113524
rect 282196 113522 282202 113524
rect 282196 113462 309426 113522
rect 282196 113460 282202 113462
rect 307569 113250 307635 113253
rect 309366 113250 309426 113462
rect 324405 113250 324471 113253
rect 307569 113248 309150 113250
rect 307569 113192 307574 113248
rect 307630 113192 309150 113248
rect 307569 113190 309150 113192
rect 309366 113190 310132 113250
rect 321908 113248 324471 113250
rect 321908 113192 324410 113248
rect 324466 113192 324471 113248
rect 321908 113190 324471 113192
rect 307569 113187 307635 113190
rect 309090 113117 309150 113190
rect 324405 113187 324471 113190
rect 252185 113114 252251 113117
rect 248860 113112 252251 113114
rect 248860 113056 252190 113112
rect 252246 113056 252251 113112
rect 248860 113054 252251 113056
rect 309090 113112 309199 113117
rect 309090 113056 309138 113112
rect 309194 113056 309199 113112
rect 309090 113054 309199 113056
rect 252185 113051 252251 113054
rect 309133 113051 309199 113054
rect 213913 112842 213979 112845
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 213913 112840 217212 112842
rect 213913 112784 213918 112840
rect 213974 112784 217212 112840
rect 213913 112782 217212 112784
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 213913 112779 213979 112782
rect 579797 112779 579863 112782
rect 251909 112706 251975 112709
rect 248860 112704 251975 112706
rect 248860 112648 251914 112704
rect 251970 112648 251975 112704
rect 248860 112646 251975 112648
rect 251909 112643 251975 112646
rect 306557 112706 306623 112709
rect 306557 112704 310132 112706
rect 306557 112648 306562 112704
rect 306618 112648 310132 112704
rect 583520 112692 584960 112782
rect 306557 112646 310132 112648
rect 306557 112643 306623 112646
rect 324313 112434 324379 112437
rect 321908 112432 324379 112434
rect 321908 112376 324318 112432
rect 324374 112376 324379 112432
rect 321908 112374 324379 112376
rect 324313 112371 324379 112374
rect 307661 112298 307727 112301
rect 307661 112296 310132 112298
rect 307661 112240 307666 112296
rect 307722 112240 310132 112296
rect 307661 112238 310132 112240
rect 307661 112235 307727 112238
rect 214741 112162 214807 112165
rect 252093 112162 252159 112165
rect 214741 112160 217212 112162
rect 214741 112104 214746 112160
rect 214802 112104 217212 112160
rect 214741 112102 217212 112104
rect 248860 112160 252159 112162
rect 248860 112104 252098 112160
rect 252154 112104 252159 112160
rect 248860 112102 252159 112104
rect 214741 112099 214807 112102
rect 252093 112099 252159 112102
rect 307293 111890 307359 111893
rect 307293 111888 310132 111890
rect 307293 111832 307298 111888
rect 307354 111832 310132 111888
rect 307293 111830 310132 111832
rect 307293 111827 307359 111830
rect 167729 111754 167795 111757
rect 252369 111754 252435 111757
rect 324313 111754 324379 111757
rect 164694 111752 167795 111754
rect 164694 111696 167734 111752
rect 167790 111696 167795 111752
rect 164694 111694 167795 111696
rect 248860 111752 252435 111754
rect 248860 111696 252374 111752
rect 252430 111696 252435 111752
rect 248860 111694 252435 111696
rect 321908 111752 324379 111754
rect 321908 111696 324318 111752
rect 324374 111696 324379 111752
rect 321908 111694 324379 111696
rect -960 110666 480 110756
rect 3141 110666 3207 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 167729 111691 167795 111694
rect 252369 111691 252435 111694
rect 324313 111691 324379 111694
rect 214005 111482 214071 111485
rect 306741 111482 306807 111485
rect 214005 111480 217212 111482
rect 214005 111424 214010 111480
rect 214066 111424 217212 111480
rect 214005 111422 217212 111424
rect 306741 111480 310132 111482
rect 306741 111424 306746 111480
rect 306802 111424 310132 111480
rect 306741 111422 310132 111424
rect 214005 111419 214071 111422
rect 306741 111419 306807 111422
rect 251950 111210 251956 111212
rect 248860 111150 251956 111210
rect 251950 111148 251956 111150
rect 252020 111148 252026 111212
rect 306557 111074 306623 111077
rect 306557 111072 310132 111074
rect 306557 111016 306562 111072
rect 306618 111016 310132 111072
rect 306557 111014 310132 111016
rect 306557 111011 306623 111014
rect 213913 110802 213979 110805
rect 251725 110802 251791 110805
rect 213913 110800 217212 110802
rect 213913 110744 213918 110800
rect 213974 110744 217212 110800
rect 213913 110742 217212 110744
rect 248860 110800 251791 110802
rect 248860 110744 251730 110800
rect 251786 110744 251791 110800
rect 248860 110742 251791 110744
rect 213913 110739 213979 110742
rect 251725 110739 251791 110742
rect 307293 110666 307359 110669
rect 307293 110664 310132 110666
rect 307293 110608 307298 110664
rect 307354 110608 310132 110664
rect 307293 110606 310132 110608
rect 307293 110603 307359 110606
rect 321878 110530 321938 110908
rect 335670 110530 335676 110532
rect 321878 110470 335676 110530
rect 335670 110468 335676 110470
rect 335740 110468 335746 110532
rect 213913 110258 213979 110261
rect 251541 110258 251607 110261
rect 213913 110256 217212 110258
rect 213913 110200 213918 110256
rect 213974 110200 217212 110256
rect 213913 110198 217212 110200
rect 248860 110256 251607 110258
rect 248860 110200 251546 110256
rect 251602 110200 251607 110256
rect 248860 110198 251607 110200
rect 213913 110195 213979 110198
rect 251541 110195 251607 110198
rect 306741 110258 306807 110261
rect 306741 110256 310132 110258
rect 306741 110200 306746 110256
rect 306802 110200 310132 110256
rect 306741 110198 310132 110200
rect 306741 110195 306807 110198
rect 167545 110122 167611 110125
rect 164694 110120 167611 110122
rect 164694 110064 167550 110120
rect 167606 110064 167611 110120
rect 164694 110062 167611 110064
rect 167545 110059 167611 110062
rect 252461 109850 252527 109853
rect 248860 109848 252527 109850
rect 248860 109792 252466 109848
rect 252522 109792 252527 109848
rect 248860 109790 252527 109792
rect 252461 109787 252527 109790
rect 307569 109850 307635 109853
rect 307569 109848 310132 109850
rect 307569 109792 307574 109848
rect 307630 109792 310132 109848
rect 307569 109790 310132 109792
rect 307569 109787 307635 109790
rect 321878 109578 321938 110092
rect 167862 109108 167868 109172
rect 167932 109170 167938 109172
rect 217182 109170 217242 109548
rect 321878 109518 325710 109578
rect 324313 109442 324379 109445
rect 321908 109440 324379 109442
rect 321908 109384 324318 109440
rect 324374 109384 324379 109440
rect 321908 109382 324379 109384
rect 324313 109379 324379 109382
rect 251449 109306 251515 109309
rect 248860 109304 251515 109306
rect 248860 109248 251454 109304
rect 251510 109248 251515 109304
rect 248860 109246 251515 109248
rect 251449 109243 251515 109246
rect 307661 109306 307727 109309
rect 307661 109304 310132 109306
rect 307661 109248 307666 109304
rect 307722 109248 310132 109304
rect 307661 109246 310132 109248
rect 307661 109243 307727 109246
rect 167932 109110 217242 109170
rect 325650 109170 325710 109518
rect 336958 109170 336964 109172
rect 325650 109110 336964 109170
rect 167932 109108 167938 109110
rect 336958 109108 336964 109110
rect 337028 109108 337034 109172
rect 214005 108898 214071 108901
rect 251173 108898 251239 108901
rect 214005 108896 217212 108898
rect 214005 108840 214010 108896
rect 214066 108840 217212 108896
rect 214005 108838 217212 108840
rect 248860 108896 251239 108898
rect 248860 108840 251178 108896
rect 251234 108840 251239 108896
rect 248860 108838 251239 108840
rect 214005 108835 214071 108838
rect 251173 108835 251239 108838
rect 307569 108898 307635 108901
rect 307569 108896 310132 108898
rect 307569 108840 307574 108896
rect 307630 108840 310132 108896
rect 307569 108838 310132 108840
rect 307569 108835 307635 108838
rect 167729 108762 167795 108765
rect 164694 108760 167795 108762
rect 164694 108704 167734 108760
rect 167790 108704 167795 108760
rect 164694 108702 167795 108704
rect 167729 108699 167795 108702
rect 324313 108626 324379 108629
rect 321908 108624 324379 108626
rect 321908 108568 324318 108624
rect 324374 108568 324379 108624
rect 321908 108566 324379 108568
rect 324313 108563 324379 108566
rect 307477 108490 307543 108493
rect 307477 108488 310132 108490
rect 307477 108432 307482 108488
rect 307538 108432 310132 108488
rect 307477 108430 310132 108432
rect 307477 108427 307543 108430
rect 251817 108354 251883 108357
rect 248860 108352 251883 108354
rect 248860 108296 251822 108352
rect 251878 108296 251883 108352
rect 248860 108294 251883 108296
rect 251817 108291 251883 108294
rect 213913 108218 213979 108221
rect 213913 108216 217212 108218
rect 213913 108160 213918 108216
rect 213974 108160 217212 108216
rect 213913 108158 217212 108160
rect 213913 108155 213979 108158
rect 307661 108082 307727 108085
rect 307661 108080 310132 108082
rect 307661 108024 307666 108080
rect 307722 108024 310132 108080
rect 307661 108022 310132 108024
rect 307661 108019 307727 108022
rect 251909 107946 251975 107949
rect 248860 107944 251975 107946
rect 248860 107888 251914 107944
rect 251970 107888 251975 107944
rect 248860 107886 251975 107888
rect 251909 107883 251975 107886
rect 305821 107810 305887 107813
rect 307569 107810 307635 107813
rect 325601 107810 325667 107813
rect 305821 107808 307635 107810
rect 305821 107752 305826 107808
rect 305882 107752 307574 107808
rect 307630 107752 307635 107808
rect 305821 107750 307635 107752
rect 321908 107808 325667 107810
rect 321908 107752 325606 107808
rect 325662 107752 325667 107808
rect 321908 107750 325667 107752
rect 305821 107747 305887 107750
rect 307569 107747 307635 107750
rect 325601 107747 325667 107750
rect 307293 107674 307359 107677
rect 307293 107672 310132 107674
rect 307293 107616 307298 107672
rect 307354 107616 310132 107672
rect 307293 107614 310132 107616
rect 307293 107611 307359 107614
rect 213913 107538 213979 107541
rect 252461 107538 252527 107541
rect 213913 107536 217212 107538
rect 213913 107480 213918 107536
rect 213974 107480 217212 107536
rect 213913 107478 217212 107480
rect 248860 107536 252527 107538
rect 248860 107480 252466 107536
rect 252522 107480 252527 107536
rect 248860 107478 252527 107480
rect 213913 107475 213979 107478
rect 252461 107475 252527 107478
rect 307477 107266 307543 107269
rect 307477 107264 310132 107266
rect 307477 107208 307482 107264
rect 307538 107208 310132 107264
rect 307477 107206 310132 107208
rect 307477 107203 307543 107206
rect 323025 107130 323091 107133
rect 321908 107128 323091 107130
rect 321908 107072 323030 107128
rect 323086 107072 323091 107128
rect 321908 107070 323091 107072
rect 323025 107067 323091 107070
rect 252369 106994 252435 106997
rect 248860 106992 252435 106994
rect 248860 106936 252374 106992
rect 252430 106936 252435 106992
rect 248860 106934 252435 106936
rect 252369 106931 252435 106934
rect 214465 106858 214531 106861
rect 307293 106858 307359 106861
rect 214465 106856 217212 106858
rect 214465 106800 214470 106856
rect 214526 106800 217212 106856
rect 214465 106798 217212 106800
rect 307293 106856 310132 106858
rect 307293 106800 307298 106856
rect 307354 106800 310132 106856
rect 307293 106798 310132 106800
rect 214465 106795 214531 106798
rect 307293 106795 307359 106798
rect 251541 106586 251607 106589
rect 248860 106584 251607 106586
rect 248860 106528 251546 106584
rect 251602 106528 251607 106584
rect 248860 106526 251607 106528
rect 251541 106523 251607 106526
rect 307661 106450 307727 106453
rect 328678 106450 328684 106452
rect 307661 106448 310132 106450
rect 307661 106392 307666 106448
rect 307722 106392 310132 106448
rect 307661 106390 310132 106392
rect 321878 106390 328684 106450
rect 307661 106387 307727 106390
rect 321878 106284 321938 106390
rect 328678 106388 328684 106390
rect 328748 106388 328754 106452
rect 214005 106178 214071 106181
rect 214005 106176 217212 106178
rect 214005 106120 214010 106176
rect 214066 106120 217212 106176
rect 214005 106118 217212 106120
rect 214005 106115 214071 106118
rect 251173 106042 251239 106045
rect 248860 106040 251239 106042
rect 248860 105984 251178 106040
rect 251234 105984 251239 106040
rect 248860 105982 251239 105984
rect 251173 105979 251239 105982
rect 306741 105906 306807 105909
rect 306741 105904 310132 105906
rect 306741 105848 306746 105904
rect 306802 105848 310132 105904
rect 306741 105846 310132 105848
rect 306741 105843 306807 105846
rect 213913 105634 213979 105637
rect 252369 105634 252435 105637
rect 213913 105632 217212 105634
rect 213913 105576 213918 105632
rect 213974 105576 217212 105632
rect 213913 105574 217212 105576
rect 248860 105632 252435 105634
rect 248860 105576 252374 105632
rect 252430 105576 252435 105632
rect 248860 105574 252435 105576
rect 213913 105571 213979 105574
rect 252369 105571 252435 105574
rect 307661 105498 307727 105501
rect 324313 105498 324379 105501
rect 307661 105496 310132 105498
rect 307661 105440 307666 105496
rect 307722 105440 310132 105496
rect 307661 105438 310132 105440
rect 321908 105496 324379 105498
rect 321908 105440 324318 105496
rect 324374 105440 324379 105496
rect 321908 105438 324379 105440
rect 307661 105435 307727 105438
rect 324313 105435 324379 105438
rect 252277 105090 252343 105093
rect 248860 105088 252343 105090
rect 248860 105032 252282 105088
rect 252338 105032 252343 105088
rect 248860 105030 252343 105032
rect 252277 105027 252343 105030
rect 305913 105090 305979 105093
rect 306741 105090 306807 105093
rect 305913 105088 306807 105090
rect 305913 105032 305918 105088
rect 305974 105032 306746 105088
rect 306802 105032 306807 105088
rect 305913 105030 306807 105032
rect 305913 105027 305979 105030
rect 306741 105027 306807 105030
rect 308262 105030 310132 105090
rect 214414 104892 214420 104956
rect 214484 104954 214490 104956
rect 305637 104954 305703 104957
rect 308262 104954 308322 105030
rect 214484 104894 217212 104954
rect 305637 104952 308322 104954
rect 305637 104896 305642 104952
rect 305698 104896 308322 104952
rect 305637 104894 308322 104896
rect 214484 104892 214490 104894
rect 305637 104891 305703 104894
rect 324313 104818 324379 104821
rect 321908 104816 324379 104818
rect 321908 104760 324318 104816
rect 324374 104760 324379 104816
rect 321908 104758 324379 104760
rect 324313 104755 324379 104758
rect 251725 104682 251791 104685
rect 248860 104680 251791 104682
rect 248860 104624 251730 104680
rect 251786 104624 251791 104680
rect 248860 104622 251791 104624
rect 251725 104619 251791 104622
rect 307477 104682 307543 104685
rect 307477 104680 310132 104682
rect 307477 104624 307482 104680
rect 307538 104624 310132 104680
rect 307477 104622 310132 104624
rect 307477 104619 307543 104622
rect 214005 104274 214071 104277
rect 307661 104274 307727 104277
rect 214005 104272 217212 104274
rect 214005 104216 214010 104272
rect 214066 104216 217212 104272
rect 214005 104214 217212 104216
rect 307661 104272 310132 104274
rect 307661 104216 307666 104272
rect 307722 104216 310132 104272
rect 307661 104214 310132 104216
rect 214005 104211 214071 104214
rect 307661 104211 307727 104214
rect 252461 104138 252527 104141
rect 248860 104136 252527 104138
rect 248860 104080 252466 104136
rect 252522 104080 252527 104136
rect 248860 104078 252527 104080
rect 252461 104075 252527 104078
rect 324313 104002 324379 104005
rect 321908 104000 324379 104002
rect 321908 103944 324318 104000
rect 324374 103944 324379 104000
rect 321908 103942 324379 103944
rect 324313 103939 324379 103942
rect 307569 103866 307635 103869
rect 307569 103864 310132 103866
rect 307569 103808 307574 103864
rect 307630 103808 310132 103864
rect 307569 103806 310132 103808
rect 307569 103803 307635 103806
rect 252001 103730 252067 103733
rect 248860 103728 252067 103730
rect 248860 103672 252006 103728
rect 252062 103672 252067 103728
rect 248860 103670 252067 103672
rect 252001 103667 252067 103670
rect 213913 103594 213979 103597
rect 213913 103592 217212 103594
rect 213913 103536 213918 103592
rect 213974 103536 217212 103592
rect 213913 103534 217212 103536
rect 213913 103531 213979 103534
rect 307569 103458 307635 103461
rect 307569 103456 310132 103458
rect 307569 103400 307574 103456
rect 307630 103400 310132 103456
rect 307569 103398 310132 103400
rect 307569 103395 307635 103398
rect 252461 103186 252527 103189
rect 322933 103186 322999 103189
rect 248860 103184 252527 103186
rect 248860 103128 252466 103184
rect 252522 103128 252527 103184
rect 248860 103126 252527 103128
rect 321908 103184 322999 103186
rect 321908 103128 322938 103184
rect 322994 103128 322999 103184
rect 321908 103126 322999 103128
rect 252461 103123 252527 103126
rect 322933 103123 322999 103126
rect 306557 103050 306623 103053
rect 306557 103048 310132 103050
rect 306557 102992 306562 103048
rect 306618 102992 310132 103048
rect 306557 102990 310132 102992
rect 306557 102987 306623 102990
rect 214005 102914 214071 102917
rect 214005 102912 217212 102914
rect 214005 102856 214010 102912
rect 214066 102856 217212 102912
rect 214005 102854 217212 102856
rect 214005 102851 214071 102854
rect 252277 102778 252343 102781
rect 248860 102776 252343 102778
rect 248860 102720 252282 102776
rect 252338 102720 252343 102776
rect 248860 102718 252343 102720
rect 252277 102715 252343 102718
rect 307661 102506 307727 102509
rect 307661 102504 310132 102506
rect 307661 102448 307666 102504
rect 307722 102448 310132 102504
rect 307661 102446 310132 102448
rect 307661 102443 307727 102446
rect 66069 102370 66135 102373
rect 68142 102370 68816 102376
rect 66069 102368 68816 102370
rect 66069 102312 66074 102368
rect 66130 102316 68816 102368
rect 66130 102312 68202 102316
rect 66069 102310 68202 102312
rect 66069 102307 66135 102310
rect 213913 102234 213979 102237
rect 252369 102234 252435 102237
rect 213913 102232 217212 102234
rect 213913 102176 213918 102232
rect 213974 102176 217212 102232
rect 213913 102174 217212 102176
rect 248860 102232 252435 102234
rect 248860 102176 252374 102232
rect 252430 102176 252435 102232
rect 248860 102174 252435 102176
rect 321878 102234 321938 102476
rect 346342 102234 346348 102236
rect 321878 102174 346348 102234
rect 213913 102171 213979 102174
rect 252369 102171 252435 102174
rect 346342 102172 346348 102174
rect 346412 102172 346418 102236
rect 307477 102098 307543 102101
rect 307477 102096 310132 102098
rect 307477 102040 307482 102096
rect 307538 102040 310132 102096
rect 307477 102038 310132 102040
rect 307477 102035 307543 102038
rect 253054 101826 253060 101828
rect 248860 101766 253060 101826
rect 253054 101764 253060 101766
rect 253124 101764 253130 101828
rect 306557 101690 306623 101693
rect 306557 101688 310132 101690
rect 306557 101632 306562 101688
rect 306618 101632 310132 101688
rect 306557 101630 310132 101632
rect 306557 101627 306623 101630
rect 214833 101554 214899 101557
rect 214833 101552 217212 101554
rect 214833 101496 214838 101552
rect 214894 101496 217212 101552
rect 214833 101494 217212 101496
rect 214833 101491 214899 101494
rect 252185 101418 252251 101421
rect 248860 101416 252251 101418
rect 248860 101360 252190 101416
rect 252246 101360 252251 101416
rect 248860 101358 252251 101360
rect 252185 101355 252251 101358
rect 307661 101282 307727 101285
rect 307661 101280 310132 101282
rect 307661 101224 307666 101280
rect 307722 101224 310132 101280
rect 307661 101222 310132 101224
rect 307661 101219 307727 101222
rect 321510 101149 321570 101660
rect 321510 101144 321619 101149
rect 321510 101088 321558 101144
rect 321614 101088 321619 101144
rect 321510 101086 321619 101088
rect 321553 101083 321619 101086
rect 213913 101010 213979 101013
rect 213913 101008 217212 101010
rect 213913 100952 213918 101008
rect 213974 100952 217212 101008
rect 213913 100950 217212 100952
rect 213913 100947 213979 100950
rect 252461 100874 252527 100877
rect 248860 100872 252527 100874
rect 248860 100816 252466 100872
rect 252522 100816 252527 100872
rect 248860 100814 252527 100816
rect 252461 100811 252527 100814
rect 305729 100874 305795 100877
rect 307477 100874 307543 100877
rect 305729 100872 307543 100874
rect 305729 100816 305734 100872
rect 305790 100816 307482 100872
rect 307538 100816 307543 100872
rect 305729 100814 307543 100816
rect 305729 100811 305795 100814
rect 307477 100811 307543 100814
rect 307661 100874 307727 100877
rect 324497 100874 324563 100877
rect 307661 100872 310132 100874
rect 307661 100816 307666 100872
rect 307722 100816 310132 100872
rect 307661 100814 310132 100816
rect 321908 100872 324563 100874
rect 321908 100816 324502 100872
rect 324558 100816 324563 100872
rect 321908 100814 324563 100816
rect 307661 100811 307727 100814
rect 324497 100811 324563 100814
rect 67725 100738 67791 100741
rect 68142 100738 68816 100744
rect 67725 100736 68816 100738
rect 67725 100680 67730 100736
rect 67786 100684 68816 100736
rect 67786 100680 68202 100684
rect 67725 100678 68202 100680
rect 67725 100675 67791 100678
rect -960 97610 480 97700
rect 2773 97610 2839 97613
rect -960 97608 2839 97610
rect -960 97552 2778 97608
rect 2834 97552 2839 97608
rect -960 97550 2839 97552
rect -960 97460 480 97550
rect 2773 97547 2839 97550
rect 252001 100466 252067 100469
rect 248860 100464 252067 100466
rect 248860 100408 252006 100464
rect 252062 100408 252067 100464
rect 248860 100406 252067 100408
rect 252001 100403 252067 100406
rect 306741 100466 306807 100469
rect 306741 100464 310132 100466
rect 306741 100408 306746 100464
rect 306802 100408 310132 100464
rect 306741 100406 310132 100408
rect 306741 100403 306807 100406
rect 214097 100330 214163 100333
rect 214097 100328 217212 100330
rect 214097 100272 214102 100328
rect 214158 100272 217212 100328
rect 214097 100270 217212 100272
rect 214097 100267 214163 100270
rect 324405 100194 324471 100197
rect 321908 100192 324471 100194
rect 321908 100136 324410 100192
rect 324466 100136 324471 100192
rect 321908 100134 324471 100136
rect 324405 100131 324471 100134
rect 306230 99996 306236 100060
rect 306300 100058 306306 100060
rect 306557 100058 306623 100061
rect 306300 99998 306436 100058
rect 306300 99996 306306 99998
rect 252461 99922 252527 99925
rect 248860 99920 252527 99922
rect 248860 99864 252466 99920
rect 252522 99864 252527 99920
rect 248860 99862 252527 99864
rect 306376 99922 306436 99998
rect 306557 100056 310132 100058
rect 306557 100000 306562 100056
rect 306618 100000 310132 100056
rect 306557 99998 310132 100000
rect 306557 99995 306623 99998
rect 309174 99922 309180 99924
rect 306376 99862 309180 99922
rect 252461 99859 252527 99862
rect 309174 99860 309180 99862
rect 309244 99860 309250 99924
rect 213913 99650 213979 99653
rect 307661 99650 307727 99653
rect 213913 99648 217212 99650
rect 213913 99592 213918 99648
rect 213974 99592 217212 99648
rect 213913 99590 217212 99592
rect 307661 99648 310132 99650
rect 307661 99592 307666 99648
rect 307722 99592 310132 99648
rect 307661 99590 310132 99592
rect 213913 99587 213979 99590
rect 307661 99587 307727 99590
rect 252093 99514 252159 99517
rect 248860 99512 252159 99514
rect 248860 99456 252098 99512
rect 252154 99456 252159 99512
rect 248860 99454 252159 99456
rect 252093 99451 252159 99454
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect 306741 99106 306807 99109
rect 306741 99104 310132 99106
rect 306741 99048 306746 99104
rect 306802 99048 310132 99104
rect 306741 99046 310132 99048
rect 306741 99043 306807 99046
rect 214005 98970 214071 98973
rect 252461 98970 252527 98973
rect 214005 98968 217212 98970
rect 214005 98912 214010 98968
rect 214066 98912 217212 98968
rect 214005 98910 217212 98912
rect 248860 98968 252527 98970
rect 248860 98912 252466 98968
rect 252522 98912 252527 98968
rect 248860 98910 252527 98912
rect 214005 98907 214071 98910
rect 252461 98907 252527 98910
rect 321694 98837 321754 99348
rect 321645 98832 321754 98837
rect 321645 98776 321650 98832
rect 321706 98776 321754 98832
rect 321645 98774 321754 98776
rect 321645 98771 321711 98774
rect 307201 98698 307267 98701
rect 307201 98696 310132 98698
rect 307201 98640 307206 98696
rect 307262 98640 310132 98696
rect 307201 98638 310132 98640
rect 307201 98635 307267 98638
rect 252369 98562 252435 98565
rect 324262 98562 324268 98564
rect 248860 98560 252435 98562
rect 248860 98504 252374 98560
rect 252430 98504 252435 98560
rect 248860 98502 252435 98504
rect 321908 98502 324268 98562
rect 252369 98499 252435 98502
rect 324262 98500 324268 98502
rect 324332 98500 324338 98564
rect 213913 98290 213979 98293
rect 307661 98290 307727 98293
rect 213913 98288 217212 98290
rect 213913 98232 213918 98288
rect 213974 98232 217212 98288
rect 213913 98230 217212 98232
rect 307661 98288 310132 98290
rect 307661 98232 307666 98288
rect 307722 98232 310132 98288
rect 307661 98230 310132 98232
rect 213913 98227 213979 98230
rect 307661 98227 307727 98230
rect 251633 98018 251699 98021
rect 248860 98016 251699 98018
rect 248860 97960 251638 98016
rect 251694 97960 251699 98016
rect 248860 97958 251699 97960
rect 251633 97955 251699 97958
rect 307569 97882 307635 97885
rect 307569 97880 310132 97882
rect 307569 97824 307574 97880
rect 307630 97824 310132 97880
rect 307569 97822 310132 97824
rect 307569 97819 307635 97822
rect 213913 97610 213979 97613
rect 252461 97610 252527 97613
rect 213913 97608 217212 97610
rect 213913 97552 213918 97608
rect 213974 97552 217212 97608
rect 213913 97550 217212 97552
rect 248860 97608 252527 97610
rect 248860 97552 252466 97608
rect 252522 97552 252527 97608
rect 248860 97550 252527 97552
rect 213913 97547 213979 97550
rect 252461 97547 252527 97550
rect 307293 97474 307359 97477
rect 307293 97472 310132 97474
rect 307293 97416 307298 97472
rect 307354 97416 310132 97472
rect 307293 97414 310132 97416
rect 307293 97411 307359 97414
rect 321510 97341 321570 97852
rect 321461 97336 321570 97341
rect 321461 97280 321466 97336
rect 321522 97280 321570 97336
rect 321461 97278 321570 97280
rect 321461 97275 321527 97278
rect 249149 97066 249215 97069
rect 264094 97066 264100 97068
rect 248860 97064 264100 97066
rect 248860 97008 249154 97064
rect 249210 97008 264100 97064
rect 248860 97006 264100 97008
rect 249149 97003 249215 97006
rect 264094 97004 264100 97006
rect 264164 97004 264170 97068
rect 307661 97066 307727 97069
rect 324589 97066 324655 97069
rect 307661 97064 310132 97066
rect 307661 97008 307666 97064
rect 307722 97008 310132 97064
rect 307661 97006 310132 97008
rect 321908 97064 324655 97066
rect 321908 97008 324594 97064
rect 324650 97008 324655 97064
rect 321908 97006 324655 97008
rect 307661 97003 307727 97006
rect 324589 97003 324655 97006
rect 214649 96930 214715 96933
rect 214649 96928 217212 96930
rect 214649 96872 214654 96928
rect 214710 96872 217212 96928
rect 214649 96870 217212 96872
rect 214649 96867 214715 96870
rect 251173 96658 251239 96661
rect 251766 96658 251772 96660
rect 248860 96656 251772 96658
rect 248860 96600 251178 96656
rect 251234 96600 251772 96656
rect 248860 96598 251772 96600
rect 251173 96595 251239 96598
rect 251766 96596 251772 96598
rect 251836 96596 251842 96660
rect 307661 96658 307727 96661
rect 307661 96656 310132 96658
rect 307661 96600 307666 96656
rect 307722 96600 310132 96656
rect 307661 96598 310132 96600
rect 307661 96595 307727 96598
rect 214557 96386 214623 96389
rect 214557 96384 217212 96386
rect 214557 96328 214562 96384
rect 214618 96328 217212 96384
rect 214557 96326 217212 96328
rect 214557 96323 214623 96326
rect 251265 96250 251331 96253
rect 248860 96248 251331 96250
rect 248860 96192 251270 96248
rect 251326 96192 251331 96248
rect 248860 96190 251331 96192
rect 251265 96187 251331 96190
rect 306925 96250 306991 96253
rect 306925 96248 310132 96250
rect 306925 96192 306930 96248
rect 306986 96192 310132 96248
rect 306925 96190 310132 96192
rect 306925 96187 306991 96190
rect 170254 95372 170260 95436
rect 170324 95434 170330 95436
rect 321326 95434 321386 96356
rect 170324 95374 321386 95434
rect 170324 95372 170330 95374
rect 66161 94890 66227 94893
rect 196893 94890 196959 94893
rect 66161 94888 196959 94890
rect 66161 94832 66166 94888
rect 66222 94832 196898 94888
rect 196954 94832 196959 94888
rect 66161 94830 196959 94832
rect 66161 94827 66227 94830
rect 196893 94827 196959 94830
rect 102041 94756 102107 94757
rect 113725 94756 113791 94757
rect 115473 94756 115539 94757
rect 133137 94756 133203 94757
rect 101984 94692 101990 94756
rect 102054 94754 102107 94756
rect 102054 94752 102146 94754
rect 102102 94696 102146 94752
rect 102054 94694 102146 94696
rect 102054 94692 102107 94694
rect 113680 94692 113686 94756
rect 113750 94754 113791 94756
rect 113750 94752 113842 94754
rect 113786 94696 113842 94752
rect 113750 94694 113842 94696
rect 113750 94692 113791 94694
rect 115448 94692 115454 94756
rect 115518 94754 115539 94756
rect 115518 94752 115610 94754
rect 115534 94696 115610 94752
rect 115518 94694 115610 94696
rect 115518 94692 115539 94694
rect 119392 94692 119398 94756
rect 119462 94754 119468 94756
rect 119654 94754 119660 94756
rect 119462 94694 119660 94754
rect 119462 94692 119468 94694
rect 119654 94692 119660 94694
rect 119724 94692 119730 94756
rect 133128 94692 133134 94756
rect 133198 94754 133204 94756
rect 133198 94694 133290 94754
rect 133198 94692 133204 94694
rect 151302 94692 151308 94756
rect 151372 94754 151378 94756
rect 151760 94754 151766 94756
rect 151372 94694 151766 94754
rect 151372 94692 151378 94694
rect 151760 94692 151766 94694
rect 151830 94692 151836 94756
rect 102041 94691 102107 94692
rect 113725 94691 113791 94692
rect 115473 94691 115539 94692
rect 133137 94691 133203 94692
rect 241513 94482 241579 94485
rect 269614 94482 269620 94484
rect 241513 94480 269620 94482
rect 241513 94424 241518 94480
rect 241574 94424 269620 94480
rect 241513 94422 269620 94424
rect 241513 94419 241579 94422
rect 269614 94420 269620 94422
rect 269684 94420 269690 94484
rect 67633 93802 67699 93805
rect 214414 93802 214420 93804
rect 67633 93800 214420 93802
rect 67633 93744 67638 93800
rect 67694 93744 214420 93800
rect 67633 93742 214420 93744
rect 67633 93739 67699 93742
rect 214414 93740 214420 93742
rect 214484 93740 214490 93804
rect 134425 93668 134491 93669
rect 151721 93668 151787 93669
rect 134374 93666 134380 93668
rect 134334 93606 134380 93666
rect 134444 93664 134491 93668
rect 151670 93666 151676 93668
rect 134486 93608 134491 93664
rect 134374 93604 134380 93606
rect 134444 93604 134491 93608
rect 151630 93606 151676 93666
rect 151740 93664 151787 93668
rect 151782 93608 151787 93664
rect 151670 93604 151676 93606
rect 151740 93604 151787 93608
rect 134425 93603 134491 93604
rect 151721 93603 151787 93604
rect 110137 93532 110203 93533
rect 118049 93532 118115 93533
rect 119521 93532 119587 93533
rect 110086 93530 110092 93532
rect 110046 93470 110092 93530
rect 110156 93528 110203 93532
rect 117998 93530 118004 93532
rect 110198 93472 110203 93528
rect 110086 93468 110092 93470
rect 110156 93468 110203 93472
rect 117958 93470 118004 93530
rect 118068 93528 118115 93532
rect 119470 93530 119476 93532
rect 118110 93472 118115 93528
rect 117998 93468 118004 93470
rect 118068 93468 118115 93472
rect 119430 93470 119476 93530
rect 119540 93528 119587 93532
rect 119582 93472 119587 93528
rect 119470 93468 119476 93470
rect 119540 93468 119587 93472
rect 110137 93467 110203 93468
rect 118049 93467 118115 93468
rect 119521 93467 119587 93468
rect 128169 93260 128235 93261
rect 128118 93258 128124 93260
rect 128078 93198 128124 93258
rect 128188 93256 128235 93260
rect 128230 93200 128235 93256
rect 128118 93196 128124 93198
rect 128188 93196 128235 93200
rect 128169 93195 128235 93196
rect 74809 92444 74875 92445
rect 74758 92442 74764 92444
rect 74718 92382 74764 92442
rect 74828 92440 74875 92444
rect 74870 92384 74875 92440
rect 74758 92380 74764 92382
rect 74828 92380 74875 92384
rect 85614 92380 85620 92444
rect 85684 92442 85690 92444
rect 85757 92442 85823 92445
rect 88057 92444 88123 92445
rect 88977 92444 89043 92445
rect 100569 92444 100635 92445
rect 109217 92444 109283 92445
rect 88006 92442 88012 92444
rect 85684 92440 85823 92442
rect 85684 92384 85762 92440
rect 85818 92384 85823 92440
rect 85684 92382 85823 92384
rect 87966 92382 88012 92442
rect 88076 92440 88123 92444
rect 88926 92442 88932 92444
rect 88118 92384 88123 92440
rect 85684 92380 85690 92382
rect 74809 92379 74875 92380
rect 85757 92379 85823 92382
rect 88006 92380 88012 92382
rect 88076 92380 88123 92384
rect 88886 92382 88932 92442
rect 88996 92440 89043 92444
rect 100518 92442 100524 92444
rect 89038 92384 89043 92440
rect 88926 92380 88932 92382
rect 88996 92380 89043 92384
rect 100478 92382 100524 92442
rect 100588 92440 100635 92444
rect 109166 92442 109172 92444
rect 100630 92384 100635 92440
rect 100518 92380 100524 92382
rect 100588 92380 100635 92384
rect 109126 92382 109172 92442
rect 109236 92440 109283 92444
rect 109278 92384 109283 92440
rect 109166 92380 109172 92382
rect 109236 92380 109283 92384
rect 111926 92380 111932 92444
rect 111996 92442 112002 92444
rect 112161 92442 112227 92445
rect 111996 92440 112227 92442
rect 111996 92384 112166 92440
rect 112222 92384 112227 92440
rect 111996 92382 112227 92384
rect 111996 92380 112002 92382
rect 88057 92379 88123 92380
rect 88977 92379 89043 92380
rect 100569 92379 100635 92380
rect 109217 92379 109283 92380
rect 112161 92379 112227 92382
rect 115054 92380 115060 92444
rect 115124 92442 115130 92444
rect 115473 92442 115539 92445
rect 116761 92444 116827 92445
rect 119705 92444 119771 92445
rect 116710 92442 116716 92444
rect 115124 92440 115539 92442
rect 115124 92384 115478 92440
rect 115534 92384 115539 92440
rect 115124 92382 115539 92384
rect 116670 92382 116716 92442
rect 116780 92440 116827 92444
rect 119654 92442 119660 92444
rect 116822 92384 116827 92440
rect 115124 92380 115130 92382
rect 115473 92379 115539 92382
rect 116710 92380 116716 92382
rect 116780 92380 116827 92384
rect 119614 92382 119660 92442
rect 119724 92440 119771 92444
rect 119766 92384 119771 92440
rect 119654 92380 119660 92382
rect 119724 92380 119771 92384
rect 125726 92380 125732 92444
rect 125796 92442 125802 92444
rect 125869 92442 125935 92445
rect 126513 92444 126579 92445
rect 130745 92444 130811 92445
rect 151537 92444 151603 92445
rect 126462 92442 126468 92444
rect 125796 92440 125935 92442
rect 125796 92384 125874 92440
rect 125930 92384 125935 92440
rect 125796 92382 125935 92384
rect 126422 92382 126468 92442
rect 126532 92440 126579 92444
rect 130694 92442 130700 92444
rect 126574 92384 126579 92440
rect 125796 92380 125802 92382
rect 116761 92379 116827 92380
rect 119705 92379 119771 92380
rect 125869 92379 125935 92382
rect 126462 92380 126468 92382
rect 126532 92380 126579 92384
rect 130654 92382 130700 92442
rect 130764 92440 130811 92444
rect 151486 92442 151492 92444
rect 130806 92384 130811 92440
rect 130694 92380 130700 92382
rect 130764 92380 130811 92384
rect 151446 92382 151492 92442
rect 151556 92440 151603 92444
rect 151598 92384 151603 92440
rect 151486 92380 151492 92382
rect 151556 92380 151603 92384
rect 152038 92380 152044 92444
rect 152108 92442 152114 92444
rect 152917 92442 152983 92445
rect 152108 92440 152983 92442
rect 152108 92384 152922 92440
rect 152978 92384 152983 92440
rect 152108 92382 152983 92384
rect 152108 92380 152114 92382
rect 126513 92379 126579 92380
rect 130745 92379 130811 92380
rect 151537 92379 151603 92380
rect 152917 92379 152983 92382
rect 171726 92380 171732 92444
rect 171796 92442 171802 92444
rect 324405 92442 324471 92445
rect 171796 92440 324471 92442
rect 171796 92384 324410 92440
rect 324466 92384 324471 92440
rect 171796 92382 324471 92384
rect 171796 92380 171802 92382
rect 324405 92379 324471 92382
rect 114134 92244 114140 92308
rect 114204 92306 114210 92308
rect 169293 92306 169359 92309
rect 114204 92304 169359 92306
rect 114204 92248 169298 92304
rect 169354 92248 169359 92304
rect 114204 92246 169359 92248
rect 114204 92244 114210 92246
rect 169293 92243 169359 92246
rect 103278 92108 103284 92172
rect 103348 92170 103354 92172
rect 174629 92170 174695 92173
rect 103348 92168 174695 92170
rect 103348 92112 174634 92168
rect 174690 92112 174695 92168
rect 103348 92110 174695 92112
rect 103348 92108 103354 92110
rect 174629 92107 174695 92110
rect 151353 92036 151419 92037
rect 151302 92034 151308 92036
rect 151262 91974 151308 92034
rect 151372 92032 151419 92036
rect 151414 91976 151419 92032
rect 151302 91972 151308 91974
rect 151372 91972 151419 91976
rect 151353 91971 151419 91972
rect 101857 91628 101923 91629
rect 101806 91626 101812 91628
rect 101766 91566 101812 91626
rect 101876 91624 101923 91628
rect 101918 91568 101923 91624
rect 101806 91564 101812 91566
rect 101876 91564 101923 91568
rect 131982 91564 131988 91628
rect 132052 91626 132058 91628
rect 132217 91626 132283 91629
rect 132052 91624 132283 91626
rect 132052 91568 132222 91624
rect 132278 91568 132283 91624
rect 132052 91566 132283 91568
rect 132052 91564 132058 91566
rect 101857 91563 101923 91564
rect 132217 91563 132283 91566
rect 98126 91428 98132 91492
rect 98196 91490 98202 91492
rect 99189 91490 99255 91493
rect 122833 91492 122899 91493
rect 98196 91488 99255 91490
rect 98196 91432 99194 91488
rect 99250 91432 99255 91488
rect 98196 91430 99255 91432
rect 98196 91428 98202 91430
rect 99189 91427 99255 91430
rect 122782 91428 122788 91492
rect 122852 91490 122899 91492
rect 122852 91488 122944 91490
rect 122894 91432 122944 91488
rect 122852 91430 122944 91432
rect 122852 91428 122899 91430
rect 122833 91427 122899 91428
rect 93894 91292 93900 91356
rect 93964 91354 93970 91356
rect 95049 91354 95115 91357
rect 97257 91356 97323 91357
rect 97206 91354 97212 91356
rect 93964 91352 95115 91354
rect 93964 91296 95054 91352
rect 95110 91296 95115 91352
rect 93964 91294 95115 91296
rect 97166 91294 97212 91354
rect 97276 91352 97323 91356
rect 97318 91296 97323 91352
rect 93964 91292 93970 91294
rect 95049 91291 95115 91294
rect 97206 91292 97212 91294
rect 97276 91292 97323 91296
rect 98494 91292 98500 91356
rect 98564 91354 98570 91356
rect 99097 91354 99163 91357
rect 98564 91352 99163 91354
rect 98564 91296 99102 91352
rect 99158 91296 99163 91352
rect 98564 91294 99163 91296
rect 98564 91292 98570 91294
rect 97257 91291 97323 91292
rect 99097 91291 99163 91294
rect 106774 91292 106780 91356
rect 106844 91354 106850 91356
rect 107009 91354 107075 91357
rect 122097 91356 122163 91357
rect 122046 91354 122052 91356
rect 106844 91352 107075 91354
rect 106844 91296 107014 91352
rect 107070 91296 107075 91352
rect 106844 91294 107075 91296
rect 122006 91294 122052 91354
rect 122116 91352 122163 91356
rect 122158 91296 122163 91352
rect 106844 91292 106850 91294
rect 107009 91291 107075 91294
rect 122046 91292 122052 91294
rect 122116 91292 122163 91296
rect 122097 91291 122163 91292
rect 124029 91356 124095 91357
rect 124029 91352 124076 91356
rect 124140 91354 124146 91356
rect 124029 91296 124034 91352
rect 124029 91292 124076 91296
rect 124140 91294 124186 91354
rect 124140 91292 124146 91294
rect 124438 91292 124444 91356
rect 124508 91354 124514 91356
rect 125409 91354 125475 91357
rect 124508 91352 125475 91354
rect 124508 91296 125414 91352
rect 125470 91296 125475 91352
rect 124508 91294 125475 91296
rect 124508 91292 124514 91294
rect 124029 91291 124095 91292
rect 125409 91291 125475 91294
rect 84326 91156 84332 91220
rect 84396 91218 84402 91220
rect 85481 91218 85547 91221
rect 84396 91216 85547 91218
rect 84396 91160 85486 91216
rect 85542 91160 85547 91216
rect 84396 91158 85547 91160
rect 84396 91156 84402 91158
rect 85481 91155 85547 91158
rect 86718 91156 86724 91220
rect 86788 91218 86794 91220
rect 86861 91218 86927 91221
rect 86788 91216 86927 91218
rect 86788 91160 86866 91216
rect 86922 91160 86927 91216
rect 86788 91158 86927 91160
rect 86788 91156 86794 91158
rect 86861 91155 86927 91158
rect 90214 91156 90220 91220
rect 90284 91218 90290 91220
rect 91001 91218 91067 91221
rect 90284 91216 91067 91218
rect 90284 91160 91006 91216
rect 91062 91160 91067 91216
rect 90284 91158 91067 91160
rect 90284 91156 90290 91158
rect 91001 91155 91067 91158
rect 91318 91156 91324 91220
rect 91388 91218 91394 91220
rect 92381 91218 92447 91221
rect 91388 91216 92447 91218
rect 91388 91160 92386 91216
rect 92442 91160 92447 91216
rect 91388 91158 92447 91160
rect 91388 91156 91394 91158
rect 92381 91155 92447 91158
rect 92606 91156 92612 91220
rect 92676 91218 92682 91220
rect 93761 91218 93827 91221
rect 92676 91216 93827 91218
rect 92676 91160 93766 91216
rect 93822 91160 93827 91216
rect 92676 91158 93827 91160
rect 92676 91156 92682 91158
rect 93761 91155 93827 91158
rect 94998 91156 95004 91220
rect 95068 91218 95074 91220
rect 95141 91218 95207 91221
rect 96153 91220 96219 91221
rect 96102 91218 96108 91220
rect 95068 91216 95207 91218
rect 95068 91160 95146 91216
rect 95202 91160 95207 91216
rect 95068 91158 95207 91160
rect 96062 91158 96108 91218
rect 96172 91216 96219 91220
rect 96214 91160 96219 91216
rect 95068 91156 95074 91158
rect 95141 91155 95207 91158
rect 96102 91156 96108 91158
rect 96172 91156 96219 91160
rect 97022 91156 97028 91220
rect 97092 91218 97098 91220
rect 97901 91218 97967 91221
rect 99281 91220 99347 91221
rect 99230 91218 99236 91220
rect 97092 91216 97967 91218
rect 97092 91160 97906 91216
rect 97962 91160 97967 91216
rect 97092 91158 97967 91160
rect 99190 91158 99236 91218
rect 99300 91216 99347 91220
rect 99342 91160 99347 91216
rect 97092 91156 97098 91158
rect 96153 91155 96219 91156
rect 97901 91155 97967 91158
rect 99230 91156 99236 91158
rect 99300 91156 99347 91160
rect 99598 91156 99604 91220
rect 99668 91218 99674 91220
rect 100477 91218 100543 91221
rect 99668 91216 100543 91218
rect 99668 91160 100482 91216
rect 100538 91160 100543 91216
rect 99668 91158 100543 91160
rect 99668 91156 99674 91158
rect 99281 91155 99347 91156
rect 100477 91155 100543 91158
rect 101622 91156 101628 91220
rect 101692 91218 101698 91220
rect 102041 91218 102107 91221
rect 101692 91216 102107 91218
rect 101692 91160 102046 91216
rect 102102 91160 102107 91216
rect 101692 91158 102107 91160
rect 101692 91156 101698 91158
rect 102041 91155 102107 91158
rect 102910 91156 102916 91220
rect 102980 91218 102986 91220
rect 103421 91218 103487 91221
rect 102980 91216 103487 91218
rect 102980 91160 103426 91216
rect 103482 91160 103487 91216
rect 102980 91158 103487 91160
rect 102980 91156 102986 91158
rect 103421 91155 103487 91158
rect 104198 91156 104204 91220
rect 104268 91218 104274 91220
rect 104341 91218 104407 91221
rect 104617 91220 104683 91221
rect 104566 91218 104572 91220
rect 104268 91216 104407 91218
rect 104268 91160 104346 91216
rect 104402 91160 104407 91216
rect 104268 91158 104407 91160
rect 104526 91158 104572 91218
rect 104636 91216 104683 91220
rect 104678 91160 104683 91216
rect 104268 91156 104274 91158
rect 104341 91155 104407 91158
rect 104566 91156 104572 91158
rect 104636 91156 104683 91160
rect 105118 91156 105124 91220
rect 105188 91218 105194 91220
rect 105721 91218 105787 91221
rect 105188 91216 105787 91218
rect 105188 91160 105726 91216
rect 105782 91160 105787 91216
rect 105188 91158 105787 91160
rect 105188 91156 105194 91158
rect 104617 91155 104683 91156
rect 105721 91155 105787 91158
rect 106038 91156 106044 91220
rect 106108 91218 106114 91220
rect 106181 91218 106247 91221
rect 106108 91216 106247 91218
rect 106108 91160 106186 91216
rect 106242 91160 106247 91216
rect 106108 91158 106247 91160
rect 106108 91156 106114 91158
rect 106181 91155 106247 91158
rect 106406 91156 106412 91220
rect 106476 91218 106482 91220
rect 107561 91218 107627 91221
rect 106476 91216 107627 91218
rect 106476 91160 107566 91216
rect 107622 91160 107627 91216
rect 106476 91158 107627 91160
rect 106476 91156 106482 91158
rect 107561 91155 107627 91158
rect 107694 91156 107700 91220
rect 107764 91218 107770 91220
rect 107837 91218 107903 91221
rect 107764 91216 107903 91218
rect 107764 91160 107842 91216
rect 107898 91160 107903 91216
rect 107764 91158 107903 91160
rect 107764 91156 107770 91158
rect 107837 91155 107903 91158
rect 108062 91156 108068 91220
rect 108132 91218 108138 91220
rect 108941 91218 109007 91221
rect 108132 91216 109007 91218
rect 108132 91160 108946 91216
rect 109002 91160 109007 91216
rect 108132 91158 109007 91160
rect 108132 91156 108138 91158
rect 108941 91155 109007 91158
rect 109534 91156 109540 91220
rect 109604 91218 109610 91220
rect 110321 91218 110387 91221
rect 109604 91216 110387 91218
rect 109604 91160 110326 91216
rect 110382 91160 110387 91216
rect 109604 91158 110387 91160
rect 109604 91156 109610 91158
rect 110321 91155 110387 91158
rect 110638 91156 110644 91220
rect 110708 91218 110714 91220
rect 110965 91218 111031 91221
rect 110708 91216 111031 91218
rect 110708 91160 110970 91216
rect 111026 91160 111031 91216
rect 110708 91158 111031 91160
rect 110708 91156 110714 91158
rect 110965 91155 111031 91158
rect 111190 91156 111196 91220
rect 111260 91218 111266 91220
rect 111425 91218 111491 91221
rect 111260 91216 111491 91218
rect 111260 91160 111430 91216
rect 111486 91160 111491 91216
rect 111260 91158 111491 91160
rect 111260 91156 111266 91158
rect 111425 91155 111491 91158
rect 112294 91156 112300 91220
rect 112364 91218 112370 91220
rect 113081 91218 113147 91221
rect 112364 91216 113147 91218
rect 112364 91160 113086 91216
rect 113142 91160 113147 91216
rect 112364 91158 113147 91160
rect 112364 91156 112370 91158
rect 113081 91155 113147 91158
rect 113214 91156 113220 91220
rect 113284 91218 113290 91220
rect 114461 91218 114527 91221
rect 115841 91220 115907 91221
rect 115790 91218 115796 91220
rect 113284 91216 114527 91218
rect 113284 91160 114466 91216
rect 114522 91160 114527 91216
rect 113284 91158 114527 91160
rect 115750 91158 115796 91218
rect 115860 91216 115907 91220
rect 115902 91160 115907 91216
rect 113284 91156 113290 91158
rect 114461 91155 114527 91158
rect 115790 91156 115796 91158
rect 115860 91156 115907 91160
rect 117078 91156 117084 91220
rect 117148 91218 117154 91220
rect 117221 91218 117287 91221
rect 118233 91220 118299 91221
rect 118182 91218 118188 91220
rect 117148 91216 117287 91218
rect 117148 91160 117226 91216
rect 117282 91160 117287 91216
rect 117148 91158 117287 91160
rect 118142 91158 118188 91218
rect 118252 91216 118299 91220
rect 118294 91160 118299 91216
rect 117148 91156 117154 91158
rect 115841 91155 115907 91156
rect 117221 91155 117287 91158
rect 118182 91156 118188 91158
rect 118252 91156 118299 91160
rect 120206 91156 120212 91220
rect 120276 91218 120282 91220
rect 120441 91218 120507 91221
rect 120276 91216 120507 91218
rect 120276 91160 120446 91216
rect 120502 91160 120507 91216
rect 120276 91158 120507 91160
rect 120276 91156 120282 91158
rect 118233 91155 118299 91156
rect 120441 91155 120507 91158
rect 120574 91156 120580 91220
rect 120644 91218 120650 91220
rect 121361 91218 121427 91221
rect 120644 91216 121427 91218
rect 120644 91160 121366 91216
rect 121422 91160 121427 91216
rect 120644 91158 121427 91160
rect 120644 91156 120650 91158
rect 121361 91155 121427 91158
rect 121678 91156 121684 91220
rect 121748 91218 121754 91220
rect 122741 91218 122807 91221
rect 121748 91216 122807 91218
rect 121748 91160 122746 91216
rect 122802 91160 122807 91216
rect 121748 91158 122807 91160
rect 121748 91156 121754 91158
rect 122741 91155 122807 91158
rect 122966 91156 122972 91220
rect 123036 91218 123042 91220
rect 124121 91218 124187 91221
rect 123036 91216 124187 91218
rect 123036 91160 124126 91216
rect 124182 91160 124187 91216
rect 123036 91158 124187 91160
rect 123036 91156 123042 91158
rect 124121 91155 124187 91158
rect 125358 91156 125364 91220
rect 125428 91218 125434 91220
rect 125501 91218 125567 91221
rect 125428 91216 125567 91218
rect 125428 91160 125506 91216
rect 125562 91160 125567 91216
rect 125428 91158 125567 91160
rect 125428 91156 125434 91158
rect 125501 91155 125567 91158
rect 126646 91156 126652 91220
rect 126716 91218 126722 91220
rect 126789 91218 126855 91221
rect 126716 91216 126855 91218
rect 126716 91160 126794 91216
rect 126850 91160 126855 91216
rect 126716 91158 126855 91160
rect 126716 91156 126722 91158
rect 126789 91155 126855 91158
rect 129406 91156 129412 91220
rect 129476 91218 129482 91220
rect 129641 91218 129707 91221
rect 129476 91216 129707 91218
rect 129476 91160 129646 91216
rect 129702 91160 129707 91216
rect 129476 91158 129707 91160
rect 129476 91156 129482 91158
rect 129641 91155 129707 91158
rect 135662 91156 135668 91220
rect 135732 91218 135738 91220
rect 136449 91218 136515 91221
rect 135732 91216 136515 91218
rect 135732 91160 136454 91216
rect 136510 91160 136515 91216
rect 135732 91158 136515 91160
rect 135732 91156 135738 91158
rect 136449 91155 136515 91158
rect 67541 91082 67607 91085
rect 324497 91082 324563 91085
rect 67541 91080 324563 91082
rect 67541 91024 67546 91080
rect 67602 91024 324502 91080
rect 324558 91024 324563 91080
rect 67541 91022 324563 91024
rect 67541 91019 67607 91022
rect 324497 91019 324563 91022
rect 63309 90946 63375 90949
rect 202321 90946 202387 90949
rect 63309 90944 202387 90946
rect 63309 90888 63314 90944
rect 63370 90888 202326 90944
rect 202382 90888 202387 90944
rect 63309 90886 202387 90888
rect 63309 90883 63375 90886
rect 202321 90883 202387 90886
rect 110965 88226 111031 88229
rect 167494 88226 167500 88228
rect 110965 88224 167500 88226
rect 110965 88168 110970 88224
rect 111026 88168 167500 88224
rect 110965 88166 167500 88168
rect 110965 88163 111031 88166
rect 167494 88164 167500 88166
rect 167564 88164 167570 88228
rect 96153 86866 96219 86869
rect 167862 86866 167868 86868
rect 96153 86864 167868 86866
rect 96153 86808 96158 86864
rect 96214 86808 167868 86864
rect 96153 86806 167868 86808
rect 96153 86803 96219 86806
rect 167862 86804 167868 86806
rect 167932 86804 167938 86868
rect 107009 86730 107075 86733
rect 166390 86730 166396 86732
rect 107009 86728 166396 86730
rect 107009 86672 107014 86728
rect 107070 86672 166396 86728
rect 107009 86670 166396 86672
rect 107009 86667 107075 86670
rect 166390 86668 166396 86670
rect 166460 86668 166466 86732
rect 583520 86186 584960 86276
rect 583342 86126 584960 86186
rect 583342 86050 583402 86126
rect 583520 86050 584960 86126
rect 583342 86036 584960 86050
rect 583342 85990 583586 86036
rect 275134 85580 275140 85644
rect 275204 85642 275210 85644
rect 583526 85642 583586 85990
rect 275204 85582 583586 85642
rect 275204 85580 275210 85582
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 106181 84146 106247 84149
rect 169150 84146 169156 84148
rect 106181 84144 169156 84146
rect 106181 84088 106186 84144
rect 106242 84088 169156 84144
rect 106181 84086 169156 84088
rect 106181 84083 106247 84086
rect 169150 84084 169156 84086
rect 169220 84084 169226 84148
rect 285765 80746 285831 80749
rect 292614 80746 292620 80748
rect 285765 80744 292620 80746
rect 285765 80688 285770 80744
rect 285826 80688 292620 80744
rect 285765 80686 292620 80688
rect 285765 80683 285831 80686
rect 292614 80684 292620 80686
rect 292684 80684 292690 80748
rect 64638 78508 64644 78572
rect 64708 78570 64714 78572
rect 324262 78570 324268 78572
rect 64708 78510 324268 78570
rect 64708 78508 64714 78510
rect 324262 78508 324268 78510
rect 324332 78508 324338 78572
rect 99281 78434 99347 78437
rect 166206 78434 166212 78436
rect 99281 78432 166212 78434
rect 99281 78376 99286 78432
rect 99342 78376 166212 78432
rect 99281 78374 166212 78376
rect 99281 78371 99347 78374
rect 166206 78372 166212 78374
rect 166276 78372 166282 78436
rect 297214 73748 297220 73812
rect 297284 73810 297290 73812
rect 321553 73810 321619 73813
rect 297284 73808 321619 73810
rect 297284 73752 321558 73808
rect 321614 73752 321619 73808
rect 297284 73750 321619 73752
rect 297284 73748 297290 73750
rect 321553 73747 321619 73750
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 49693 62794 49759 62797
rect 307150 62794 307156 62796
rect 49693 62792 307156 62794
rect 49693 62736 49698 62792
rect 49754 62736 307156 62792
rect 49693 62734 307156 62736
rect 49693 62731 49759 62734
rect 307150 62732 307156 62734
rect 307220 62732 307226 62796
rect 177062 61372 177068 61436
rect 177132 61434 177138 61436
rect 356697 61434 356763 61437
rect 177132 61432 356763 61434
rect 177132 61376 356702 61432
rect 356758 61376 356763 61432
rect 177132 61374 356763 61376
rect 177132 61372 177138 61374
rect 356697 61371 356763 61374
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 56593 55858 56659 55861
rect 295926 55858 295932 55860
rect 56593 55856 295932 55858
rect 56593 55800 56598 55856
rect 56654 55800 295932 55856
rect 56593 55798 295932 55800
rect 56593 55795 56659 55798
rect 295926 55796 295932 55798
rect 295996 55796 296002 55860
rect 174854 53076 174860 53140
rect 174924 53138 174930 53140
rect 336733 53138 336799 53141
rect 174924 53136 336799 53138
rect 174924 53080 336738 53136
rect 336794 53080 336799 53136
rect 174924 53078 336799 53080
rect 174924 53076 174930 53078
rect 336733 53075 336799 53078
rect 265566 47500 265572 47564
rect 265636 47562 265642 47564
rect 580165 47562 580231 47565
rect 265636 47560 580231 47562
rect 265636 47504 580170 47560
rect 580226 47504 580231 47560
rect 265636 47502 580231 47504
rect 265636 47500 265642 47502
rect 580165 47499 580231 47502
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 9673 46202 9739 46205
rect 300158 46202 300164 46204
rect 9673 46200 300164 46202
rect 9673 46144 9678 46200
rect 9734 46144 300164 46200
rect 9673 46142 300164 46144
rect 9673 46139 9739 46142
rect 300158 46140 300164 46142
rect 300228 46140 300234 46204
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 62113 44842 62179 44845
rect 305494 44842 305500 44844
rect 62113 44840 305500 44842
rect 62113 44784 62118 44840
rect 62174 44784 305500 44840
rect 62113 44782 305500 44784
rect 62113 44779 62179 44782
rect 305494 44780 305500 44782
rect 305564 44780 305570 44844
rect 582465 33146 582531 33149
rect 583520 33146 584960 33236
rect 582465 33144 584960 33146
rect 582465 33088 582470 33144
rect 582526 33088 584960 33144
rect 582465 33086 584960 33088
rect 582465 33083 582531 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 179822 25604 179828 25668
rect 179892 25666 179898 25668
rect 303613 25666 303679 25669
rect 179892 25664 303679 25666
rect 179892 25608 303618 25664
rect 303674 25608 303679 25664
rect 179892 25606 303679 25608
rect 179892 25604 179898 25606
rect 303613 25603 303679 25606
rect 66253 25530 66319 25533
rect 304206 25530 304212 25532
rect 66253 25528 304212 25530
rect 66253 25472 66258 25528
rect 66314 25472 304212 25528
rect 66253 25470 304212 25472
rect 66253 25467 66319 25470
rect 304206 25468 304212 25470
rect 304276 25468 304282 25532
rect 175038 22612 175044 22676
rect 175108 22674 175114 22676
rect 339493 22674 339559 22677
rect 175108 22672 339559 22674
rect 175108 22616 339498 22672
rect 339554 22616 339559 22672
rect 175108 22614 339559 22616
rect 175108 22612 175114 22614
rect 339493 22611 339559 22614
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 176326 18668 176332 18732
rect 176396 18730 176402 18732
rect 313273 18730 313339 18733
rect 176396 18728 313339 18730
rect 176396 18672 313278 18728
rect 313334 18672 313339 18728
rect 176396 18670 313339 18672
rect 176396 18668 176402 18670
rect 313273 18667 313339 18670
rect 12433 18594 12499 18597
rect 282126 18594 282132 18596
rect 12433 18592 282132 18594
rect 12433 18536 12438 18592
rect 12494 18536 282132 18592
rect 12433 18534 282132 18536
rect 12433 18531 12499 18534
rect 282126 18532 282132 18534
rect 282196 18532 282202 18596
rect 22093 17234 22159 17237
rect 306966 17234 306972 17236
rect 22093 17232 306972 17234
rect 22093 17176 22098 17232
rect 22154 17176 306972 17232
rect 22093 17174 306972 17176
rect 22093 17171 22159 17174
rect 306966 17172 306972 17174
rect 307036 17172 307042 17236
rect 176510 12956 176516 13020
rect 176580 13018 176586 13020
rect 331213 13018 331279 13021
rect 176580 13016 331279 13018
rect 176580 12960 331218 13016
rect 331274 12960 331279 13016
rect 176580 12958 331279 12960
rect 176580 12956 176586 12958
rect 331213 12955 331279 12958
rect 582373 6626 582439 6629
rect 583520 6626 584960 6716
rect 582373 6624 584960 6626
rect -960 6490 480 6580
rect 582373 6568 582378 6624
rect 582434 6568 584960 6624
rect 582373 6566 584960 6568
rect 582373 6563 582439 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 305545 6354 305611 6357
rect 331254 6354 331260 6356
rect 305545 6352 331260 6354
rect 305545 6296 305550 6352
rect 305606 6296 331260 6352
rect 305545 6294 331260 6296
rect 305545 6291 305611 6294
rect 331254 6292 331260 6294
rect 331324 6292 331330 6356
rect 303153 6218 303219 6221
rect 332542 6218 332548 6220
rect 303153 6216 332548 6218
rect 303153 6160 303158 6216
rect 303214 6160 332548 6216
rect 303153 6158 332548 6160
rect 303153 6155 303219 6158
rect 332542 6156 332548 6158
rect 332612 6156 332618 6220
rect 52545 4858 52611 4861
rect 299974 4858 299980 4860
rect 52545 4856 299980 4858
rect 52545 4800 52550 4856
rect 52606 4800 299980 4856
rect 52545 4798 299980 4800
rect 52545 4795 52611 4798
rect 299974 4796 299980 4798
rect 300044 4796 300050 4860
rect 301446 3980 301452 4044
rect 301516 4042 301522 4044
rect 309041 4042 309107 4045
rect 301516 4040 309107 4042
rect 301516 3984 309046 4040
rect 309102 3984 309107 4040
rect 301516 3982 309107 3984
rect 301516 3980 301522 3982
rect 309041 3979 309107 3982
rect 251030 3436 251036 3500
rect 251100 3498 251106 3500
rect 255865 3498 255931 3501
rect 251100 3496 255931 3498
rect 251100 3440 255870 3496
rect 255926 3440 255931 3496
rect 251100 3438 255931 3440
rect 251100 3436 251106 3438
rect 255865 3435 255931 3438
rect 292798 3436 292804 3500
rect 292868 3498 292874 3500
rect 293677 3498 293743 3501
rect 292868 3496 293743 3498
rect 292868 3440 293682 3496
rect 293738 3440 293743 3496
rect 292868 3438 293743 3440
rect 292868 3436 292874 3438
rect 293677 3435 293743 3438
rect 296069 3498 296135 3501
rect 309174 3498 309180 3500
rect 296069 3496 309180 3498
rect 296069 3440 296074 3496
rect 296130 3440 309180 3496
rect 296069 3438 309180 3440
rect 296069 3435 296135 3438
rect 309174 3436 309180 3438
rect 309244 3436 309250 3500
rect 342161 3498 342227 3501
rect 342294 3498 342300 3500
rect 342161 3496 342300 3498
rect 342161 3440 342166 3496
rect 342222 3440 342300 3496
rect 342161 3438 342300 3440
rect 342161 3435 342227 3438
rect 342294 3436 342300 3438
rect 342364 3436 342370 3500
rect 170990 3300 170996 3364
rect 171060 3362 171066 3364
rect 242893 3362 242959 3365
rect 171060 3360 242959 3362
rect 171060 3304 242898 3360
rect 242954 3304 242959 3360
rect 171060 3302 242959 3304
rect 171060 3300 171066 3302
rect 242893 3299 242959 3302
rect 264145 3362 264211 3365
rect 271086 3362 271092 3364
rect 264145 3360 271092 3362
rect 264145 3304 264150 3360
rect 264206 3304 271092 3360
rect 264145 3302 271092 3304
rect 264145 3299 264211 3302
rect 271086 3300 271092 3302
rect 271156 3300 271162 3364
rect 307937 3362 308003 3365
rect 336774 3362 336780 3364
rect 307937 3360 336780 3362
rect 307937 3304 307942 3360
rect 307998 3304 336780 3360
rect 307937 3302 336780 3304
rect 307937 3299 308003 3302
rect 336774 3300 336780 3302
rect 336844 3300 336850 3364
<< obsm3 >>
rect 68800 171594 164756 174600
rect 68800 171534 164694 171594
rect 68800 129304 164756 171534
rect 68816 129244 164756 129304
rect 68800 128080 164756 129244
rect 68816 128020 164756 128080
rect 68800 126312 164756 128020
rect 68816 126252 164756 126312
rect 68800 125224 164756 126252
rect 68816 125164 164756 125224
rect 68800 123592 164756 125164
rect 68816 123532 164756 123592
rect 68800 122640 164756 123532
rect 68816 122580 164756 122640
rect 68800 120872 164756 122580
rect 68816 120812 164756 120872
rect 68800 111754 164756 120812
rect 68800 111694 164694 111754
rect 68800 110122 164756 111694
rect 68800 110062 164694 110122
rect 68800 108762 164756 110062
rect 68800 108702 164694 108762
rect 68800 102376 164756 108702
rect 68816 102316 164756 102376
rect 68800 100744 164756 102316
rect 68816 100684 164756 100744
rect 68800 95100 164756 100684
<< via3 >>
rect 179276 702612 179340 702676
rect 180564 702476 180628 702540
rect 120028 514796 120092 514860
rect 299980 484468 300044 484532
rect 342300 363020 342364 363084
rect 332548 361660 332612 361724
rect 293908 358804 293972 358868
rect 152964 357716 153028 357780
rect 170996 357580 171060 357644
rect 297220 357580 297284 357644
rect 292804 356220 292868 356284
rect 301452 356084 301516 356148
rect 70900 354724 70964 354788
rect 179828 351868 179892 351932
rect 175044 350100 175108 350164
rect 295380 349556 295444 349620
rect 292620 346972 292684 347036
rect 293908 345476 293972 345540
rect 156460 345068 156524 345132
rect 177068 339220 177132 339284
rect 174860 330380 174924 330444
rect 176516 327660 176580 327724
rect 176332 323580 176396 323644
rect 170260 296788 170324 296852
rect 171916 295292 171980 295356
rect 119660 294204 119724 294268
rect 119292 292844 119356 292908
rect 64644 288628 64708 288692
rect 119660 289172 119724 289236
rect 119292 288084 119356 288148
rect 179276 283596 179340 283660
rect 293908 281556 293972 281620
rect 57836 278836 57900 278900
rect 59124 271900 59188 271964
rect 70532 267412 70596 267476
rect 153700 263604 153764 263668
rect 157932 258028 157996 258092
rect 64460 257212 64524 257276
rect 120580 256940 120644 257004
rect 160692 255444 160756 255508
rect 178540 255308 178604 255372
rect 119292 254084 119356 254148
rect 161980 251228 162044 251292
rect 61884 248508 61948 248572
rect 120028 247964 120092 248028
rect 299612 247072 299676 247076
rect 299612 247016 299662 247072
rect 299662 247016 299676 247072
rect 299612 247012 299676 247016
rect 63356 245788 63420 245852
rect 120948 245924 121012 245988
rect 179828 242932 179892 242996
rect 120948 242524 121012 242588
rect 63172 241708 63236 241772
rect 291700 241028 291764 241092
rect 119108 239804 119172 239868
rect 178540 238988 178604 239052
rect 161980 238852 162044 238916
rect 293908 238716 293972 238780
rect 57836 238580 57900 238644
rect 171916 238444 171980 238508
rect 299980 238444 300044 238508
rect 171732 238036 171796 238100
rect 265572 238036 265636 238100
rect 328500 237900 328564 237964
rect 156460 237220 156524 237284
rect 160692 237220 160756 237284
rect 120580 237084 120644 237148
rect 64460 236540 64524 236604
rect 61884 235860 61948 235924
rect 295380 235860 295444 235924
rect 322060 233820 322124 233884
rect 63172 233140 63236 233204
rect 59124 231780 59188 231844
rect 153700 231644 153764 231708
rect 63356 230420 63420 230484
rect 299612 230420 299676 230484
rect 269620 229740 269684 229804
rect 271092 228244 271156 228308
rect 157932 227564 157996 227628
rect 273852 226884 273916 226948
rect 291700 226884 291764 226948
rect 251220 225524 251284 225588
rect 336964 221444 337028 221508
rect 260972 215868 261036 215932
rect 327212 214508 327276 214572
rect 265020 213148 265084 213212
rect 335860 211924 335924 211988
rect 335676 211788 335740 211852
rect 346348 210564 346412 210628
rect 269068 210428 269132 210492
rect 328684 210292 328748 210356
rect 263548 206348 263612 206412
rect 255268 206212 255332 206276
rect 331260 204852 331324 204916
rect 340828 200636 340892 200700
rect 270540 199276 270604 199340
rect 327028 197916 327092 197980
rect 152964 193836 153028 193900
rect 259684 192612 259748 192676
rect 329788 192476 329852 192540
rect 259500 190980 259564 191044
rect 260972 189620 261036 189684
rect 306236 189620 306300 189684
rect 254532 188260 254596 188324
rect 320404 186900 320468 186964
rect 256924 185540 256988 185604
rect 266308 184316 266372 184380
rect 332732 182820 332796 182884
rect 255452 181460 255516 181524
rect 256740 180100 256804 180164
rect 249012 179964 249076 180028
rect 334020 178740 334084 178804
rect 249196 177652 249260 177716
rect 99420 177516 99484 177580
rect 101996 177576 102060 177580
rect 101996 177520 102046 177576
rect 102046 177520 102060 177576
rect 101996 177516 102060 177520
rect 106044 177516 106108 177580
rect 106964 177516 107028 177580
rect 112116 177516 112180 177580
rect 114140 177516 114204 177580
rect 116900 177576 116964 177580
rect 116900 177520 116950 177576
rect 116950 177520 116964 177576
rect 116900 177516 116964 177520
rect 118372 177516 118436 177580
rect 127020 177516 127084 177580
rect 129412 177576 129476 177580
rect 129412 177520 129462 177576
rect 129462 177520 129476 177576
rect 129412 177516 129476 177520
rect 133092 177516 133156 177580
rect 331444 177380 331508 177444
rect 257844 177244 257908 177308
rect 336780 177244 336844 177308
rect 110644 177168 110708 177172
rect 110644 177112 110694 177168
rect 110694 177112 110708 177168
rect 110644 177108 110708 177112
rect 113220 177108 113284 177172
rect 103284 176972 103348 177036
rect 97028 176836 97092 176900
rect 100708 176836 100772 176900
rect 166212 176836 166276 176900
rect 108068 176760 108132 176764
rect 108068 176704 108118 176760
rect 108118 176704 108132 176760
rect 108068 176700 108132 176704
rect 109540 176700 109604 176764
rect 119660 176760 119724 176764
rect 119660 176704 119710 176760
rect 119710 176704 119724 176760
rect 119660 176700 119724 176704
rect 121868 176700 121932 176764
rect 122972 176760 123036 176764
rect 122972 176704 123022 176760
rect 123022 176704 123036 176760
rect 122972 176700 123036 176704
rect 124444 176700 124508 176764
rect 125732 176700 125796 176764
rect 131988 176760 132052 176764
rect 131988 176704 132038 176760
rect 132038 176704 132052 176760
rect 131988 176700 132052 176704
rect 134380 176760 134444 176764
rect 134380 176704 134430 176760
rect 134430 176704 134444 176760
rect 134380 176700 134444 176704
rect 135668 176760 135732 176764
rect 135668 176704 135718 176760
rect 135718 176704 135732 176760
rect 135668 176700 135732 176704
rect 148180 176760 148244 176764
rect 148180 176704 148230 176760
rect 148230 176704 148244 176760
rect 148180 176700 148244 176704
rect 158852 176700 158916 176764
rect 264100 176700 264164 176764
rect 320220 176760 320284 176764
rect 320220 176704 320234 176760
rect 320234 176704 320284 176760
rect 320220 176700 320284 176704
rect 128124 176428 128188 176492
rect 321508 176156 321572 176220
rect 252508 176020 252572 176084
rect 98316 175476 98380 175540
rect 104572 175536 104636 175540
rect 104572 175480 104622 175536
rect 104622 175480 104636 175536
rect 104572 175476 104636 175480
rect 120764 175536 120828 175540
rect 120764 175480 120814 175536
rect 120814 175480 120828 175536
rect 120764 175476 120828 175480
rect 130700 175536 130764 175540
rect 130700 175480 130750 175536
rect 130750 175480 130764 175536
rect 130700 175476 130764 175480
rect 115726 174992 115790 174996
rect 115726 174936 115754 174992
rect 115754 174936 115790 174992
rect 115726 174932 115790 174936
rect 214420 174524 214484 174588
rect 249196 174252 249260 174316
rect 249380 173708 249444 173772
rect 321508 172076 321572 172140
rect 321324 171396 321388 171460
rect 321324 170580 321388 170644
rect 214420 168948 214484 169012
rect 256924 168540 256988 168604
rect 251036 166228 251100 166292
rect 269068 163100 269132 163164
rect 266308 162964 266372 163028
rect 265020 162148 265084 162212
rect 275140 162012 275204 162076
rect 260788 161468 260852 161532
rect 256740 161060 256804 161124
rect 166212 160652 166276 160716
rect 255452 158204 255516 158268
rect 307156 157388 307220 157452
rect 306972 154804 307036 154868
rect 257844 152900 257908 152964
rect 251956 149636 252020 149700
rect 307156 148276 307220 148340
rect 252508 147868 252572 147932
rect 254532 146916 254596 146980
rect 335676 145556 335740 145620
rect 327212 145420 327276 145484
rect 263548 144604 263612 144668
rect 322060 144604 322124 144668
rect 306972 144060 307036 144124
rect 259684 142156 259748 142220
rect 253428 141340 253492 141404
rect 260972 141204 261036 141268
rect 251220 140796 251284 140860
rect 270540 139708 270604 139772
rect 255268 139436 255332 139500
rect 273852 138620 273916 138684
rect 259500 138484 259564 138548
rect 334020 138076 334084 138140
rect 167500 134132 167564 134196
rect 331444 134132 331508 134196
rect 332732 133860 332796 133924
rect 166396 132500 166460 132564
rect 169156 131412 169220 131476
rect 251772 131684 251836 131748
rect 295932 131412 295996 131476
rect 307156 130596 307220 130660
rect 166212 128556 166276 128620
rect 300164 126380 300228 126444
rect 328500 125564 328564 125628
rect 329788 123252 329852 123316
rect 327028 121620 327092 121684
rect 304212 119036 304276 119100
rect 305500 118628 305564 118692
rect 299980 117404 300044 117468
rect 340828 114548 340892 114612
rect 306972 114004 307036 114068
rect 282132 113460 282196 113524
rect 251956 111148 252020 111212
rect 335676 110468 335740 110532
rect 167868 109108 167932 109172
rect 336964 109108 337028 109172
rect 328684 106388 328748 106452
rect 214420 104892 214484 104956
rect 346348 102172 346412 102236
rect 253060 101764 253124 101828
rect 306236 99996 306300 100060
rect 309180 99860 309244 99924
rect 324268 98500 324332 98564
rect 264100 97004 264164 97068
rect 251772 96596 251836 96660
rect 170260 95372 170324 95436
rect 101990 94752 102054 94756
rect 101990 94696 102046 94752
rect 102046 94696 102054 94752
rect 101990 94692 102054 94696
rect 113686 94752 113750 94756
rect 113686 94696 113730 94752
rect 113730 94696 113750 94752
rect 113686 94692 113750 94696
rect 115454 94752 115518 94756
rect 115454 94696 115478 94752
rect 115478 94696 115518 94752
rect 115454 94692 115518 94696
rect 119398 94692 119462 94756
rect 119660 94692 119724 94756
rect 133134 94752 133198 94756
rect 133134 94696 133142 94752
rect 133142 94696 133198 94752
rect 133134 94692 133198 94696
rect 151308 94692 151372 94756
rect 151766 94692 151830 94756
rect 269620 94420 269684 94484
rect 214420 93740 214484 93804
rect 134380 93664 134444 93668
rect 134380 93608 134430 93664
rect 134430 93608 134444 93664
rect 134380 93604 134444 93608
rect 151676 93664 151740 93668
rect 151676 93608 151726 93664
rect 151726 93608 151740 93664
rect 151676 93604 151740 93608
rect 110092 93528 110156 93532
rect 110092 93472 110142 93528
rect 110142 93472 110156 93528
rect 110092 93468 110156 93472
rect 118004 93528 118068 93532
rect 118004 93472 118054 93528
rect 118054 93472 118068 93528
rect 118004 93468 118068 93472
rect 119476 93528 119540 93532
rect 119476 93472 119526 93528
rect 119526 93472 119540 93528
rect 119476 93468 119540 93472
rect 128124 93256 128188 93260
rect 128124 93200 128174 93256
rect 128174 93200 128188 93256
rect 128124 93196 128188 93200
rect 74764 92440 74828 92444
rect 74764 92384 74814 92440
rect 74814 92384 74828 92440
rect 74764 92380 74828 92384
rect 85620 92380 85684 92444
rect 88012 92440 88076 92444
rect 88012 92384 88062 92440
rect 88062 92384 88076 92440
rect 88012 92380 88076 92384
rect 88932 92440 88996 92444
rect 88932 92384 88982 92440
rect 88982 92384 88996 92440
rect 88932 92380 88996 92384
rect 100524 92440 100588 92444
rect 100524 92384 100574 92440
rect 100574 92384 100588 92440
rect 100524 92380 100588 92384
rect 109172 92440 109236 92444
rect 109172 92384 109222 92440
rect 109222 92384 109236 92440
rect 109172 92380 109236 92384
rect 111932 92380 111996 92444
rect 115060 92380 115124 92444
rect 116716 92440 116780 92444
rect 116716 92384 116766 92440
rect 116766 92384 116780 92440
rect 116716 92380 116780 92384
rect 119660 92440 119724 92444
rect 119660 92384 119710 92440
rect 119710 92384 119724 92440
rect 119660 92380 119724 92384
rect 125732 92380 125796 92444
rect 126468 92440 126532 92444
rect 126468 92384 126518 92440
rect 126518 92384 126532 92440
rect 126468 92380 126532 92384
rect 130700 92440 130764 92444
rect 130700 92384 130750 92440
rect 130750 92384 130764 92440
rect 130700 92380 130764 92384
rect 151492 92440 151556 92444
rect 151492 92384 151542 92440
rect 151542 92384 151556 92440
rect 151492 92380 151556 92384
rect 152044 92380 152108 92444
rect 171732 92380 171796 92444
rect 114140 92244 114204 92308
rect 103284 92108 103348 92172
rect 151308 92032 151372 92036
rect 151308 91976 151358 92032
rect 151358 91976 151372 92032
rect 151308 91972 151372 91976
rect 101812 91624 101876 91628
rect 101812 91568 101862 91624
rect 101862 91568 101876 91624
rect 101812 91564 101876 91568
rect 131988 91564 132052 91628
rect 98132 91428 98196 91492
rect 122788 91488 122852 91492
rect 122788 91432 122838 91488
rect 122838 91432 122852 91488
rect 122788 91428 122852 91432
rect 93900 91292 93964 91356
rect 97212 91352 97276 91356
rect 97212 91296 97262 91352
rect 97262 91296 97276 91352
rect 97212 91292 97276 91296
rect 98500 91292 98564 91356
rect 106780 91292 106844 91356
rect 122052 91352 122116 91356
rect 122052 91296 122102 91352
rect 122102 91296 122116 91352
rect 122052 91292 122116 91296
rect 124076 91352 124140 91356
rect 124076 91296 124090 91352
rect 124090 91296 124140 91352
rect 124076 91292 124140 91296
rect 124444 91292 124508 91356
rect 84332 91156 84396 91220
rect 86724 91156 86788 91220
rect 90220 91156 90284 91220
rect 91324 91156 91388 91220
rect 92612 91156 92676 91220
rect 95004 91156 95068 91220
rect 96108 91216 96172 91220
rect 96108 91160 96158 91216
rect 96158 91160 96172 91216
rect 96108 91156 96172 91160
rect 97028 91156 97092 91220
rect 99236 91216 99300 91220
rect 99236 91160 99286 91216
rect 99286 91160 99300 91216
rect 99236 91156 99300 91160
rect 99604 91156 99668 91220
rect 101628 91156 101692 91220
rect 102916 91156 102980 91220
rect 104204 91156 104268 91220
rect 104572 91216 104636 91220
rect 104572 91160 104622 91216
rect 104622 91160 104636 91216
rect 104572 91156 104636 91160
rect 105124 91156 105188 91220
rect 106044 91156 106108 91220
rect 106412 91156 106476 91220
rect 107700 91156 107764 91220
rect 108068 91156 108132 91220
rect 109540 91156 109604 91220
rect 110644 91156 110708 91220
rect 111196 91156 111260 91220
rect 112300 91156 112364 91220
rect 113220 91156 113284 91220
rect 115796 91216 115860 91220
rect 115796 91160 115846 91216
rect 115846 91160 115860 91216
rect 115796 91156 115860 91160
rect 117084 91156 117148 91220
rect 118188 91216 118252 91220
rect 118188 91160 118238 91216
rect 118238 91160 118252 91216
rect 118188 91156 118252 91160
rect 120212 91156 120276 91220
rect 120580 91156 120644 91220
rect 121684 91156 121748 91220
rect 122972 91156 123036 91220
rect 125364 91156 125428 91220
rect 126652 91156 126716 91220
rect 129412 91156 129476 91220
rect 135668 91156 135732 91220
rect 167500 88164 167564 88228
rect 167868 86804 167932 86868
rect 166396 86668 166460 86732
rect 275140 85580 275204 85644
rect 169156 84084 169220 84148
rect 292620 80684 292684 80748
rect 64644 78508 64708 78572
rect 324268 78508 324332 78572
rect 166212 78372 166276 78436
rect 297220 73748 297284 73812
rect 307156 62732 307220 62796
rect 177068 61372 177132 61436
rect 295932 55796 295996 55860
rect 174860 53076 174924 53140
rect 265572 47500 265636 47564
rect 300164 46140 300228 46204
rect 305500 44780 305564 44844
rect 179828 25604 179892 25668
rect 304212 25468 304276 25532
rect 175044 22612 175108 22676
rect 176332 18668 176396 18732
rect 282132 18532 282196 18596
rect 306972 17172 307036 17236
rect 176516 12956 176580 13020
rect 331260 6292 331324 6356
rect 332548 6156 332612 6220
rect 299980 4796 300044 4860
rect 301452 3980 301516 4044
rect 251036 3436 251100 3500
rect 292804 3436 292868 3500
rect 309180 3436 309244 3500
rect 342300 3436 342364 3500
rect 170996 3300 171060 3364
rect 271092 3300 271156 3364
rect 336780 3300 336844 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 57835 278900 57901 278901
rect 57835 278836 57836 278900
rect 57900 278836 57901 278900
rect 57835 278835 57901 278836
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 57838 238645 57898 278835
rect 60294 277954 60914 313398
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64643 288692 64709 288693
rect 64643 288628 64644 288692
rect 64708 288628 64709 288692
rect 64643 288627 64709 288628
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 59123 271964 59189 271965
rect 59123 271900 59124 271964
rect 59188 271900 59189 271964
rect 59123 271899 59189 271900
rect 57835 238644 57901 238645
rect 57835 238580 57836 238644
rect 57900 238580 57901 238644
rect 57835 238579 57901 238580
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 59126 231845 59186 271899
rect 60294 241954 60914 277398
rect 64459 257276 64525 257277
rect 64459 257212 64460 257276
rect 64524 257212 64525 257276
rect 64459 257211 64525 257212
rect 61883 248572 61949 248573
rect 61883 248508 61884 248572
rect 61948 248508 61949 248572
rect 61883 248507 61949 248508
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 59123 231844 59189 231845
rect 59123 231780 59124 231844
rect 59188 231780 59189 231844
rect 59123 231779 59189 231780
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 205954 60914 241398
rect 61886 235925 61946 248507
rect 63355 245852 63421 245853
rect 63355 245788 63356 245852
rect 63420 245788 63421 245852
rect 63355 245787 63421 245788
rect 63171 241772 63237 241773
rect 63171 241708 63172 241772
rect 63236 241708 63237 241772
rect 63171 241707 63237 241708
rect 61883 235924 61949 235925
rect 61883 235860 61884 235924
rect 61948 235860 61949 235924
rect 61883 235859 61949 235860
rect 63174 233205 63234 241707
rect 63171 233204 63237 233205
rect 63171 233140 63172 233204
rect 63236 233140 63237 233204
rect 63171 233139 63237 233140
rect 63358 230485 63418 245787
rect 64462 236605 64522 257211
rect 64459 236604 64525 236605
rect 64459 236540 64460 236604
rect 64524 236540 64525 236604
rect 64459 236539 64525 236540
rect 63355 230484 63421 230485
rect 63355 230420 63356 230484
rect 63420 230420 63421 230484
rect 63355 230419 63421 230420
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 64646 78573 64706 288627
rect 64794 282454 65414 317898
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 70899 354788 70965 354789
rect 70899 354724 70900 354788
rect 70964 354724 70965 354788
rect 70899 354723 70965 354724
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 294000 69914 322398
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 70902 267750 70962 354723
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 294000 74414 326898
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 294000 78914 295398
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 294000 83414 299898
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 294000 87914 304398
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 294000 92414 308898
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 294000 96914 313398
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 294000 101414 317898
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 294000 105914 322398
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 294000 110414 326898
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 294000 114914 295398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 120027 514860 120093 514861
rect 120027 514796 120028 514860
rect 120092 514796 120093 514860
rect 120027 514795 120093 514796
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 294000 119414 299898
rect 119659 294268 119725 294269
rect 119659 294204 119660 294268
rect 119724 294204 119725 294268
rect 119659 294203 119725 294204
rect 119291 292908 119357 292909
rect 119291 292844 119292 292908
rect 119356 292844 119357 292908
rect 119291 292843 119357 292844
rect 119294 288149 119354 292843
rect 119662 289237 119722 294203
rect 119659 289236 119725 289237
rect 119659 289172 119660 289236
rect 119724 289172 119725 289236
rect 119659 289171 119725 289172
rect 119291 288148 119357 288149
rect 119291 288084 119292 288148
rect 119356 288084 119357 288148
rect 119291 288083 119357 288084
rect 70534 267690 70962 267750
rect 70534 267477 70594 267690
rect 70531 267476 70597 267477
rect 70531 267412 70532 267476
rect 70596 267412 70597 267476
rect 70531 267411 70597 267412
rect 89568 259954 89888 259986
rect 89568 259718 89610 259954
rect 89846 259718 89888 259954
rect 89568 259634 89888 259718
rect 89568 259398 89610 259634
rect 89846 259398 89888 259634
rect 89568 259366 89888 259398
rect 74208 255454 74528 255486
rect 74208 255218 74250 255454
rect 74486 255218 74528 255454
rect 74208 255134 74528 255218
rect 74208 254898 74250 255134
rect 74486 254898 74528 255134
rect 74208 254866 74528 254898
rect 104928 255454 105248 255486
rect 104928 255218 104970 255454
rect 105206 255218 105248 255454
rect 104928 255134 105248 255218
rect 104928 254898 104970 255134
rect 105206 254898 105248 255134
rect 104928 254866 105248 254898
rect 119291 254148 119357 254149
rect 119291 254084 119292 254148
rect 119356 254084 119357 254148
rect 119291 254083 119357 254084
rect 119294 248430 119354 254083
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 119110 248370 119354 248430
rect 119110 239869 119170 248370
rect 120030 248029 120090 514795
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 120579 257004 120645 257005
rect 120579 256940 120580 257004
rect 120644 256940 120645 257004
rect 120579 256939 120645 256940
rect 120027 248028 120093 248029
rect 120027 247964 120028 248028
rect 120092 247964 120093 248028
rect 120027 247963 120093 247964
rect 119107 239868 119173 239869
rect 119107 239804 119108 239868
rect 119172 239804 119173 239868
rect 119107 239803 119173 239804
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 69294 214954 69914 238000
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 176600 69914 178398
rect 73794 219454 74414 238000
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 176600 74414 182898
rect 78294 223954 78914 238000
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 176600 78914 187398
rect 82794 228454 83414 238000
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 176600 83414 191898
rect 87294 232954 87914 238000
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 176600 87914 196398
rect 91794 237454 92414 238000
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 176600 92414 200898
rect 105294 214954 105914 238000
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 99419 177580 99485 177581
rect 99419 177516 99420 177580
rect 99484 177516 99485 177580
rect 99419 177515 99485 177516
rect 101995 177580 102061 177581
rect 101995 177516 101996 177580
rect 102060 177516 102061 177580
rect 101995 177515 102061 177516
rect 97027 176900 97093 176901
rect 97027 176836 97028 176900
rect 97092 176836 97093 176900
rect 97027 176835 97093 176836
rect 97030 175130 97090 176835
rect 98315 175540 98381 175541
rect 98315 175476 98316 175540
rect 98380 175476 98381 175540
rect 98315 175475 98381 175476
rect 96960 175070 97090 175130
rect 98318 175130 98378 175475
rect 99422 175130 99482 177515
rect 100707 176900 100773 176901
rect 100707 176836 100708 176900
rect 100772 176836 100773 176900
rect 100707 176835 100773 176836
rect 98318 175070 98380 175130
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64643 78572 64709 78573
rect 64643 78508 64644 78572
rect 64708 78508 64709 78572
rect 64643 78507 64709 78508
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 66454 65414 101898
rect 96960 174494 97020 175070
rect 98320 174494 98380 175070
rect 99408 175070 99482 175130
rect 100710 175130 100770 176835
rect 101998 175130 102058 177515
rect 103283 177036 103349 177037
rect 103283 176972 103284 177036
rect 103348 176972 103349 177036
rect 103283 176971 103349 176972
rect 100710 175070 100828 175130
rect 99408 174494 99468 175070
rect 100768 174494 100828 175070
rect 101992 175070 102058 175130
rect 103286 175130 103346 176971
rect 105294 176600 105914 178398
rect 109794 219454 110414 238000
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 106043 177580 106109 177581
rect 106043 177516 106044 177580
rect 106108 177516 106109 177580
rect 106043 177515 106109 177516
rect 106963 177580 107029 177581
rect 106963 177516 106964 177580
rect 107028 177516 107029 177580
rect 106963 177515 107029 177516
rect 104571 175540 104637 175541
rect 104571 175476 104572 175540
rect 104636 175476 104637 175540
rect 104571 175475 104637 175476
rect 104574 175130 104634 175475
rect 106046 175130 106106 177515
rect 103286 175070 103412 175130
rect 104574 175070 104636 175130
rect 101992 174494 102052 175070
rect 103352 174494 103412 175070
rect 104576 174494 104636 175070
rect 105664 175070 106106 175130
rect 106966 175130 107026 177515
rect 108067 176764 108133 176765
rect 108067 176700 108068 176764
rect 108132 176700 108133 176764
rect 108067 176699 108133 176700
rect 109539 176764 109605 176765
rect 109539 176700 109540 176764
rect 109604 176700 109605 176764
rect 109539 176699 109605 176700
rect 108070 175130 108130 176699
rect 109542 175130 109602 176699
rect 109794 176600 110414 182898
rect 114294 223954 114914 238000
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 112115 177580 112181 177581
rect 112115 177516 112116 177580
rect 112180 177516 112181 177580
rect 112115 177515 112181 177516
rect 114139 177580 114205 177581
rect 114139 177516 114140 177580
rect 114204 177516 114205 177580
rect 114139 177515 114205 177516
rect 110643 177172 110709 177173
rect 110643 177108 110644 177172
rect 110708 177108 110709 177172
rect 110643 177107 110709 177108
rect 106966 175070 107084 175130
rect 108070 175070 108172 175130
rect 105664 174494 105724 175070
rect 107024 174494 107084 175070
rect 108112 174494 108172 175070
rect 109472 175070 109602 175130
rect 110646 175130 110706 177107
rect 112118 175130 112178 177515
rect 113219 177172 113285 177173
rect 113219 177108 113220 177172
rect 113284 177108 113285 177172
rect 113219 177107 113285 177108
rect 113222 175130 113282 177107
rect 110646 175070 110756 175130
rect 109472 174494 109532 175070
rect 110696 174494 110756 175070
rect 112056 175070 112178 175130
rect 113144 175070 113282 175130
rect 114142 175130 114202 177515
rect 114294 176600 114914 187398
rect 118794 228454 119414 238000
rect 120582 237149 120642 256939
rect 120947 245988 121013 245989
rect 120947 245924 120948 245988
rect 121012 245924 121013 245988
rect 120947 245923 121013 245924
rect 120950 242589 121010 245923
rect 120947 242588 121013 242589
rect 120947 242524 120948 242588
rect 121012 242524 121013 242588
rect 120947 242523 121013 242524
rect 120579 237148 120645 237149
rect 120579 237084 120580 237148
rect 120644 237084 120645 237148
rect 120579 237083 120645 237084
rect 118794 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 119414 228454
rect 118794 228134 119414 228218
rect 118794 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 119414 228134
rect 118794 192454 119414 227898
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 116899 177580 116965 177581
rect 116899 177516 116900 177580
rect 116964 177516 116965 177580
rect 116899 177515 116965 177516
rect 118371 177580 118437 177581
rect 118371 177516 118372 177580
rect 118436 177516 118437 177580
rect 118371 177515 118437 177516
rect 116902 175130 116962 177515
rect 118374 175130 118434 177515
rect 118794 176600 119414 191898
rect 123294 232954 123914 268398
rect 123294 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 123914 232954
rect 123294 232634 123914 232718
rect 123294 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 123914 232634
rect 123294 196954 123914 232398
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 119659 176764 119725 176765
rect 119659 176700 119660 176764
rect 119724 176700 119725 176764
rect 119659 176699 119725 176700
rect 121867 176764 121933 176765
rect 121867 176700 121868 176764
rect 121932 176700 121933 176764
rect 121867 176699 121933 176700
rect 122971 176764 123037 176765
rect 122971 176700 122972 176764
rect 123036 176700 123037 176764
rect 122971 176699 123037 176700
rect 119662 175130 119722 176699
rect 120763 175540 120829 175541
rect 120763 175476 120764 175540
rect 120828 175476 120829 175540
rect 120763 175475 120829 175476
rect 120766 175130 120826 175475
rect 121870 175130 121930 176699
rect 114142 175070 114428 175130
rect 116902 175070 117012 175130
rect 112056 174494 112116 175070
rect 113144 174494 113204 175070
rect 114368 174494 114428 175070
rect 115725 174996 115791 174997
rect 115725 174932 115726 174996
rect 115790 174932 115791 174996
rect 115725 174931 115791 174932
rect 115728 174494 115788 174931
rect 116952 174494 117012 175070
rect 118312 175070 118434 175130
rect 119400 175070 119722 175130
rect 120760 175070 120826 175130
rect 121848 175070 121930 175130
rect 122974 175130 123034 176699
rect 123294 176600 123914 196398
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127019 177580 127085 177581
rect 127019 177516 127020 177580
rect 127084 177516 127085 177580
rect 127019 177515 127085 177516
rect 124443 176764 124509 176765
rect 124443 176700 124444 176764
rect 124508 176700 124509 176764
rect 124443 176699 124509 176700
rect 125731 176764 125797 176765
rect 125731 176700 125732 176764
rect 125796 176700 125797 176764
rect 125731 176699 125797 176700
rect 124446 175130 124506 176699
rect 125734 175130 125794 176699
rect 127022 175130 127082 177515
rect 127794 176600 128414 200898
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 241954 132914 277398
rect 132294 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 132914 241954
rect 132294 241634 132914 241718
rect 132294 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 132914 241634
rect 132294 205954 132914 241398
rect 132294 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 132914 205954
rect 132294 205634 132914 205718
rect 132294 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 132914 205634
rect 129411 177580 129477 177581
rect 129411 177516 129412 177580
rect 129476 177516 129477 177580
rect 129411 177515 129477 177516
rect 128123 176492 128189 176493
rect 128123 176428 128124 176492
rect 128188 176428 128189 176492
rect 128123 176427 128189 176428
rect 128126 175130 128186 176427
rect 122974 175070 123132 175130
rect 118312 174494 118372 175070
rect 119400 174494 119460 175070
rect 120760 174494 120820 175070
rect 121848 174494 121908 175070
rect 123072 174494 123132 175070
rect 124432 175070 124506 175130
rect 125656 175070 125794 175130
rect 127016 175070 127082 175130
rect 128104 175070 128186 175130
rect 129414 175130 129474 177515
rect 131987 176764 132053 176765
rect 131987 176700 131988 176764
rect 132052 176700 132053 176764
rect 131987 176699 132053 176700
rect 130699 175540 130765 175541
rect 130699 175476 130700 175540
rect 130764 175476 130765 175540
rect 130699 175475 130765 175476
rect 130702 175130 130762 175475
rect 129414 175070 129524 175130
rect 124432 174494 124492 175070
rect 125656 174494 125716 175070
rect 127016 174494 127076 175070
rect 128104 174494 128164 175070
rect 129464 174494 129524 175070
rect 130688 175070 130762 175130
rect 131990 175130 132050 176699
rect 132294 176600 132914 205398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 246454 137414 281898
rect 136794 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 137414 246454
rect 136794 246134 137414 246218
rect 136794 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 137414 246134
rect 136794 210454 137414 245898
rect 136794 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 137414 210454
rect 136794 210134 137414 210218
rect 136794 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 137414 210134
rect 133091 177580 133157 177581
rect 133091 177516 133092 177580
rect 133156 177516 133157 177580
rect 133091 177515 133157 177516
rect 133094 175130 133154 177515
rect 134379 176764 134445 176765
rect 134379 176700 134380 176764
rect 134444 176700 134445 176764
rect 134379 176699 134445 176700
rect 135667 176764 135733 176765
rect 135667 176700 135668 176764
rect 135732 176700 135733 176764
rect 135667 176699 135733 176700
rect 134382 175130 134442 176699
rect 131990 175070 132108 175130
rect 133094 175070 133196 175130
rect 130688 174494 130748 175070
rect 132048 174494 132108 175070
rect 133136 174494 133196 175070
rect 134360 175070 134442 175130
rect 135670 175130 135730 176699
rect 136794 176600 137414 209898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 214954 141914 250398
rect 141294 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 141914 214954
rect 141294 214634 141914 214718
rect 141294 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 141914 214634
rect 141294 178954 141914 214398
rect 141294 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 141914 178954
rect 141294 178634 141914 178718
rect 141294 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 141914 178634
rect 141294 176600 141914 178398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 176600 146414 182898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 152963 357780 153029 357781
rect 152963 357716 152964 357780
rect 153028 357716 153029 357780
rect 152963 357715 153029 357716
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 223954 150914 259398
rect 150294 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 150914 223954
rect 150294 223634 150914 223718
rect 150294 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 150914 223634
rect 150294 187954 150914 223398
rect 152966 193901 153026 357715
rect 154794 336454 155414 371898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 156459 345132 156525 345133
rect 156459 345068 156460 345132
rect 156524 345068 156525 345132
rect 156459 345067 156525 345068
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 153699 263668 153765 263669
rect 153699 263604 153700 263668
rect 153764 263604 153765 263668
rect 153699 263603 153765 263604
rect 153702 231709 153762 263603
rect 153699 231708 153765 231709
rect 153699 231644 153700 231708
rect 153764 231644 153765 231708
rect 153699 231643 153765 231644
rect 154794 228454 155414 263898
rect 156462 237285 156522 345067
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 157931 258092 157997 258093
rect 157931 258028 157932 258092
rect 157996 258028 157997 258092
rect 157931 258027 157997 258028
rect 156459 237284 156525 237285
rect 156459 237220 156460 237284
rect 156524 237220 156525 237284
rect 156459 237219 156525 237220
rect 154794 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 155414 228454
rect 154794 228134 155414 228218
rect 154794 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 155414 228134
rect 152963 193900 153029 193901
rect 152963 193836 152964 193900
rect 153028 193836 153029 193900
rect 152963 193835 153029 193836
rect 150294 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 150914 187954
rect 150294 187634 150914 187718
rect 150294 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 150914 187634
rect 148179 176764 148245 176765
rect 148179 176700 148180 176764
rect 148244 176700 148245 176764
rect 148179 176699 148245 176700
rect 148182 175130 148242 176699
rect 150294 176600 150914 187398
rect 154794 192454 155414 227898
rect 157934 227629 157994 258027
rect 159294 232954 159914 268398
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 160691 255508 160757 255509
rect 160691 255444 160692 255508
rect 160756 255444 160757 255508
rect 160691 255443 160757 255444
rect 160694 237285 160754 255443
rect 161979 251292 162045 251293
rect 161979 251228 161980 251292
rect 162044 251228 162045 251292
rect 161979 251227 162045 251228
rect 161982 238917 162042 251227
rect 161979 238916 162045 238917
rect 161979 238852 161980 238916
rect 162044 238852 162045 238916
rect 161979 238851 162045 238852
rect 163794 237454 164414 272898
rect 160691 237284 160757 237285
rect 160691 237220 160692 237284
rect 160756 237220 160757 237284
rect 160691 237219 160757 237220
rect 159294 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 159914 232954
rect 159294 232634 159914 232718
rect 159294 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 159914 232634
rect 157931 227628 157997 227629
rect 157931 227564 157932 227628
rect 157996 227564 157997 227628
rect 157931 227563 157997 227564
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 154794 176600 155414 191898
rect 159294 196954 159914 232398
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 159294 196634 159914 196718
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 158851 176764 158917 176765
rect 158851 176700 158852 176764
rect 158916 176700 158917 176764
rect 158851 176699 158917 176700
rect 158854 175130 158914 176699
rect 159294 176600 159914 196398
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 176600 164414 200898
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 170995 357644 171061 357645
rect 170995 357580 170996 357644
rect 171060 357580 171061 357644
rect 170995 357579 171061 357580
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 170259 296852 170325 296853
rect 170259 296788 170260 296852
rect 170324 296788 170325 296852
rect 170259 296787 170325 296788
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 241954 168914 277398
rect 168294 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 168914 241954
rect 168294 241634 168914 241718
rect 168294 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 168914 241634
rect 168294 205954 168914 241398
rect 168294 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 168914 205954
rect 168294 205634 168914 205718
rect 168294 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 168914 205634
rect 166211 176900 166277 176901
rect 166211 176836 166212 176900
rect 166276 176836 166277 176900
rect 166211 176835 166277 176836
rect 135670 175070 135780 175130
rect 148182 175070 148292 175130
rect 134360 174494 134420 175070
rect 135720 174494 135780 175070
rect 148232 174494 148292 175070
rect 158840 175070 158914 175130
rect 158840 174494 158900 175070
rect 166214 160717 166274 176835
rect 168294 169954 168914 205398
rect 168294 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 168914 169954
rect 168294 169634 168914 169718
rect 168294 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 168914 169634
rect 166211 160716 166277 160717
rect 166211 160652 166212 160716
rect 166276 160652 166277 160716
rect 166211 160651 166277 160652
rect 69072 151954 69420 151986
rect 69072 151718 69128 151954
rect 69364 151718 69420 151954
rect 69072 151634 69420 151718
rect 69072 151398 69128 151634
rect 69364 151398 69420 151634
rect 69072 151366 69420 151398
rect 164136 151954 164484 151986
rect 164136 151718 164192 151954
rect 164428 151718 164484 151954
rect 164136 151634 164484 151718
rect 164136 151398 164192 151634
rect 164428 151398 164484 151634
rect 164136 151366 164484 151398
rect 69752 147454 70100 147486
rect 69752 147218 69808 147454
rect 70044 147218 70100 147454
rect 69752 147134 70100 147218
rect 69752 146898 69808 147134
rect 70044 146898 70100 147134
rect 69752 146866 70100 146898
rect 163456 147454 163804 147486
rect 163456 147218 163512 147454
rect 163748 147218 163804 147454
rect 163456 147134 163804 147218
rect 163456 146898 163512 147134
rect 163748 146898 163804 147134
rect 163456 146866 163804 146898
rect 167499 134196 167565 134197
rect 167499 134132 167500 134196
rect 167564 134132 167565 134196
rect 167499 134131 167565 134132
rect 166395 132564 166461 132565
rect 166395 132500 166396 132564
rect 166460 132500 166461 132564
rect 166395 132499 166461 132500
rect 166211 128620 166277 128621
rect 166211 128556 166212 128620
rect 166276 128556 166277 128620
rect 166211 128555 166277 128556
rect 69072 115954 69420 115986
rect 69072 115718 69128 115954
rect 69364 115718 69420 115954
rect 69072 115634 69420 115718
rect 69072 115398 69128 115634
rect 69364 115398 69420 115634
rect 69072 115366 69420 115398
rect 164136 115954 164484 115986
rect 164136 115718 164192 115954
rect 164428 115718 164484 115954
rect 164136 115634 164484 115718
rect 164136 115398 164192 115634
rect 164428 115398 164484 115634
rect 164136 115366 164484 115398
rect 69752 111454 70100 111486
rect 69752 111218 69808 111454
rect 70044 111218 70100 111454
rect 69752 111134 70100 111218
rect 69752 110898 69808 111134
rect 70044 110898 70100 111134
rect 69752 110866 70100 110898
rect 163456 111454 163804 111486
rect 163456 111218 163512 111454
rect 163748 111218 163804 111454
rect 163456 111134 163804 111218
rect 163456 110898 163512 111134
rect 163748 110898 163804 111134
rect 163456 110866 163804 110898
rect 74656 94890 74716 95200
rect 84312 94890 84372 95200
rect 85536 94890 85596 95200
rect 86624 94890 86684 95200
rect 87984 94890 88044 95200
rect 88936 94890 88996 95200
rect 74656 94830 74826 94890
rect 84312 94830 84394 94890
rect 85536 94830 85682 94890
rect 86624 94830 86786 94890
rect 87984 94830 88074 94890
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 70954 69914 93100
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 75454 74414 93100
rect 74766 92445 74826 94830
rect 74763 92444 74829 92445
rect 74763 92380 74764 92444
rect 74828 92380 74829 92444
rect 74763 92379 74829 92380
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 79954 78914 93100
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 84454 83414 93100
rect 84334 91221 84394 94830
rect 85622 92445 85682 94830
rect 85619 92444 85685 92445
rect 85619 92380 85620 92444
rect 85684 92380 85685 92444
rect 85619 92379 85685 92380
rect 86726 91221 86786 94830
rect 84331 91220 84397 91221
rect 84331 91156 84332 91220
rect 84396 91156 84397 91220
rect 84331 91155 84397 91156
rect 86723 91220 86789 91221
rect 86723 91156 86724 91220
rect 86788 91156 86789 91220
rect 86723 91155 86789 91156
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 88954 87914 93100
rect 88014 92445 88074 94830
rect 88934 94830 88996 94890
rect 90160 94890 90220 95200
rect 91384 94890 91444 95200
rect 90160 94830 90282 94890
rect 88934 92445 88994 94830
rect 88011 92444 88077 92445
rect 88011 92380 88012 92444
rect 88076 92380 88077 92444
rect 88011 92379 88077 92380
rect 88931 92444 88997 92445
rect 88931 92380 88932 92444
rect 88996 92380 88997 92444
rect 88931 92379 88997 92380
rect 90222 91221 90282 94830
rect 91326 94830 91444 94890
rect 92472 94890 92532 95200
rect 93832 94890 93892 95200
rect 94920 94890 94980 95200
rect 96008 94890 96068 95200
rect 96688 94890 96748 95200
rect 97096 94890 97156 95200
rect 98048 94890 98108 95200
rect 98456 94890 98516 95200
rect 99136 94890 99196 95200
rect 99544 94890 99604 95200
rect 100632 94890 100692 95200
rect 92472 94830 92674 94890
rect 93832 94830 93962 94890
rect 94920 94830 95066 94890
rect 96008 94830 96170 94890
rect 96688 94830 96906 94890
rect 97096 94830 97274 94890
rect 98048 94830 98194 94890
rect 98456 94830 98562 94890
rect 99136 94830 99298 94890
rect 99544 94830 99666 94890
rect 91326 91221 91386 94830
rect 90219 91220 90285 91221
rect 90219 91156 90220 91220
rect 90284 91156 90285 91220
rect 90219 91155 90285 91156
rect 91323 91220 91389 91221
rect 91323 91156 91324 91220
rect 91388 91156 91389 91220
rect 91323 91155 91389 91156
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 57454 92414 93100
rect 92614 91221 92674 94830
rect 93902 91357 93962 94830
rect 93899 91356 93965 91357
rect 93899 91292 93900 91356
rect 93964 91292 93965 91356
rect 93899 91291 93965 91292
rect 95006 91221 95066 94830
rect 96110 91221 96170 94830
rect 96846 93870 96906 94830
rect 96846 93810 97090 93870
rect 92611 91220 92677 91221
rect 92611 91156 92612 91220
rect 92676 91156 92677 91220
rect 92611 91155 92677 91156
rect 95003 91220 95069 91221
rect 95003 91156 95004 91220
rect 95068 91156 95069 91220
rect 95003 91155 95069 91156
rect 96107 91220 96173 91221
rect 96107 91156 96108 91220
rect 96172 91156 96173 91220
rect 96107 91155 96173 91156
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 61954 96914 93100
rect 97030 91221 97090 93810
rect 97214 91357 97274 94830
rect 98134 91493 98194 94830
rect 98131 91492 98197 91493
rect 98131 91428 98132 91492
rect 98196 91428 98197 91492
rect 98131 91427 98197 91428
rect 98502 91357 98562 94830
rect 97211 91356 97277 91357
rect 97211 91292 97212 91356
rect 97276 91292 97277 91356
rect 97211 91291 97277 91292
rect 98499 91356 98565 91357
rect 98499 91292 98500 91356
rect 98564 91292 98565 91356
rect 98499 91291 98565 91292
rect 99238 91221 99298 94830
rect 99606 91221 99666 94830
rect 100526 94830 100692 94890
rect 100768 94890 100828 95200
rect 101856 94890 101916 95200
rect 100768 94830 101690 94890
rect 100526 92445 100586 94830
rect 100523 92444 100589 92445
rect 100523 92380 100524 92444
rect 100588 92380 100589 92444
rect 100523 92379 100589 92380
rect 97027 91220 97093 91221
rect 97027 91156 97028 91220
rect 97092 91156 97093 91220
rect 97027 91155 97093 91156
rect 99235 91220 99301 91221
rect 99235 91156 99236 91220
rect 99300 91156 99301 91220
rect 99235 91155 99301 91156
rect 99603 91220 99669 91221
rect 99603 91156 99604 91220
rect 99668 91156 99669 91220
rect 99603 91155 99669 91156
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 66454 101414 93100
rect 101630 91221 101690 94830
rect 101814 94830 101916 94890
rect 101814 91629 101874 94830
rect 101992 94757 102052 95200
rect 102944 94890 103004 95200
rect 102918 94830 103004 94890
rect 103216 94890 103276 95200
rect 104304 94890 104364 95200
rect 103216 94830 103346 94890
rect 101989 94756 102055 94757
rect 101989 94692 101990 94756
rect 102054 94692 102055 94756
rect 101989 94691 102055 94692
rect 101811 91628 101877 91629
rect 101811 91564 101812 91628
rect 101876 91564 101877 91628
rect 101811 91563 101877 91564
rect 102918 91221 102978 94830
rect 103286 92173 103346 94830
rect 104206 94830 104364 94890
rect 104440 94890 104500 95200
rect 105392 94890 105452 95200
rect 104440 94830 104634 94890
rect 103283 92172 103349 92173
rect 103283 92108 103284 92172
rect 103348 92108 103349 92172
rect 103283 92107 103349 92108
rect 104206 91221 104266 94830
rect 104574 91221 104634 94830
rect 105126 94830 105452 94890
rect 105664 94890 105724 95200
rect 106480 94890 106540 95200
rect 105664 94830 106106 94890
rect 105126 91221 105186 94830
rect 101627 91220 101693 91221
rect 101627 91156 101628 91220
rect 101692 91156 101693 91220
rect 101627 91155 101693 91156
rect 102915 91220 102981 91221
rect 102915 91156 102916 91220
rect 102980 91156 102981 91220
rect 102915 91155 102981 91156
rect 104203 91220 104269 91221
rect 104203 91156 104204 91220
rect 104268 91156 104269 91220
rect 104203 91155 104269 91156
rect 104571 91220 104637 91221
rect 104571 91156 104572 91220
rect 104636 91156 104637 91220
rect 104571 91155 104637 91156
rect 105123 91220 105189 91221
rect 105123 91156 105124 91220
rect 105188 91156 105189 91220
rect 105123 91155 105189 91156
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 70954 105914 93100
rect 106046 91221 106106 94830
rect 106414 94830 106540 94890
rect 106616 94890 106676 95200
rect 107704 94890 107764 95200
rect 108112 94890 108172 95200
rect 106616 94830 106842 94890
rect 106414 91221 106474 94830
rect 106782 91357 106842 94830
rect 107702 94830 107764 94890
rect 108070 94830 108172 94890
rect 109064 94890 109124 95200
rect 109472 94890 109532 95200
rect 110152 94890 110212 95200
rect 110696 94890 110756 95200
rect 111240 94890 111300 95200
rect 109064 94830 109234 94890
rect 109472 94830 109602 94890
rect 106779 91356 106845 91357
rect 106779 91292 106780 91356
rect 106844 91292 106845 91356
rect 106779 91291 106845 91292
rect 107702 91221 107762 94830
rect 108070 91221 108130 94830
rect 109174 92445 109234 94830
rect 109171 92444 109237 92445
rect 109171 92380 109172 92444
rect 109236 92380 109237 92444
rect 109171 92379 109237 92380
rect 109542 91221 109602 94830
rect 110094 94830 110212 94890
rect 110646 94830 110756 94890
rect 111198 94830 111300 94890
rect 111920 94890 111980 95200
rect 112328 94890 112388 95200
rect 111920 94830 111994 94890
rect 110094 93533 110154 94830
rect 110091 93532 110157 93533
rect 110091 93468 110092 93532
rect 110156 93468 110157 93532
rect 110091 93467 110157 93468
rect 106043 91220 106109 91221
rect 106043 91156 106044 91220
rect 106108 91156 106109 91220
rect 106043 91155 106109 91156
rect 106411 91220 106477 91221
rect 106411 91156 106412 91220
rect 106476 91156 106477 91220
rect 106411 91155 106477 91156
rect 107699 91220 107765 91221
rect 107699 91156 107700 91220
rect 107764 91156 107765 91220
rect 107699 91155 107765 91156
rect 108067 91220 108133 91221
rect 108067 91156 108068 91220
rect 108132 91156 108133 91220
rect 108067 91155 108133 91156
rect 109539 91220 109605 91221
rect 109539 91156 109540 91220
rect 109604 91156 109605 91220
rect 109539 91155 109605 91156
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 75454 110414 93100
rect 110646 91221 110706 94830
rect 111198 91221 111258 94830
rect 111934 92445 111994 94830
rect 112302 94830 112388 94890
rect 113144 94890 113204 95200
rect 113144 94830 113282 94890
rect 111931 92444 111997 92445
rect 111931 92380 111932 92444
rect 111996 92380 111997 92444
rect 111931 92379 111997 92380
rect 112302 91221 112362 94830
rect 113222 91221 113282 94830
rect 113688 94757 113748 95200
rect 114368 94890 114428 95200
rect 114142 94830 114428 94890
rect 114776 94890 114836 95200
rect 114776 94830 115122 94890
rect 113685 94756 113751 94757
rect 113685 94692 113686 94756
rect 113750 94692 113751 94756
rect 113685 94691 113751 94692
rect 114142 92309 114202 94830
rect 114139 92308 114205 92309
rect 114139 92244 114140 92308
rect 114204 92244 114205 92308
rect 114139 92243 114205 92244
rect 110643 91220 110709 91221
rect 110643 91156 110644 91220
rect 110708 91156 110709 91220
rect 110643 91155 110709 91156
rect 111195 91220 111261 91221
rect 111195 91156 111196 91220
rect 111260 91156 111261 91220
rect 111195 91155 111261 91156
rect 112299 91220 112365 91221
rect 112299 91156 112300 91220
rect 112364 91156 112365 91220
rect 112299 91155 112365 91156
rect 113219 91220 113285 91221
rect 113219 91156 113220 91220
rect 113284 91156 113285 91220
rect 113219 91155 113285 91156
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 79954 114914 93100
rect 115062 92445 115122 94830
rect 115456 94757 115516 95200
rect 115864 94890 115924 95200
rect 115798 94830 115924 94890
rect 116680 94890 116740 95200
rect 117088 94890 117148 95200
rect 116680 94830 116778 94890
rect 115453 94756 115519 94757
rect 115453 94692 115454 94756
rect 115518 94692 115519 94756
rect 115453 94691 115519 94692
rect 115059 92444 115125 92445
rect 115059 92380 115060 92444
rect 115124 92380 115125 92444
rect 115059 92379 115125 92380
rect 115798 91221 115858 94830
rect 116718 92445 116778 94830
rect 117086 94830 117148 94890
rect 117904 94890 117964 95200
rect 118176 94890 118236 95200
rect 117904 94830 118066 94890
rect 118176 94830 118250 94890
rect 116715 92444 116781 92445
rect 116715 92380 116716 92444
rect 116780 92380 116781 92444
rect 116715 92379 116781 92380
rect 117086 91221 117146 94830
rect 118006 93533 118066 94830
rect 118003 93532 118069 93533
rect 118003 93468 118004 93532
rect 118068 93468 118069 93532
rect 118003 93467 118069 93468
rect 118190 91221 118250 94830
rect 119400 94757 119460 95200
rect 119397 94756 119463 94757
rect 119397 94692 119398 94756
rect 119462 94692 119463 94756
rect 119397 94691 119463 94692
rect 119536 94210 119596 95200
rect 120216 94890 120276 95200
rect 120624 94890 120684 95200
rect 121712 94890 121772 95200
rect 120214 94830 120276 94890
rect 120582 94830 120684 94890
rect 121686 94830 121772 94890
rect 121984 94890 122044 95200
rect 121984 94830 122114 94890
rect 119659 94756 119725 94757
rect 119659 94692 119660 94756
rect 119724 94692 119725 94756
rect 119659 94691 119725 94692
rect 119478 94150 119596 94210
rect 119478 93533 119538 94150
rect 119475 93532 119541 93533
rect 119475 93468 119476 93532
rect 119540 93468 119541 93532
rect 119475 93467 119541 93468
rect 115795 91220 115861 91221
rect 115795 91156 115796 91220
rect 115860 91156 115861 91220
rect 115795 91155 115861 91156
rect 117083 91220 117149 91221
rect 117083 91156 117084 91220
rect 117148 91156 117149 91220
rect 117083 91155 117149 91156
rect 118187 91220 118253 91221
rect 118187 91156 118188 91220
rect 118252 91156 118253 91220
rect 118187 91155 118253 91156
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114294 43954 114914 79398
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 84454 119414 93100
rect 119662 92445 119722 94691
rect 119659 92444 119725 92445
rect 119659 92380 119660 92444
rect 119724 92380 119725 92444
rect 119659 92379 119725 92380
rect 120214 91221 120274 94830
rect 120582 91221 120642 94830
rect 121686 91221 121746 94830
rect 122054 91357 122114 94830
rect 122800 93870 122860 95200
rect 123208 94890 123268 95200
rect 122606 93810 122860 93870
rect 122974 94830 123268 94890
rect 124024 94890 124084 95200
rect 124432 94890 124492 95200
rect 125384 94890 125444 95200
rect 124024 94830 124138 94890
rect 124432 94830 124506 94890
rect 122606 91490 122666 93810
rect 122787 91492 122853 91493
rect 122787 91490 122788 91492
rect 122606 91430 122788 91490
rect 122787 91428 122788 91430
rect 122852 91428 122853 91492
rect 122787 91427 122853 91428
rect 122051 91356 122117 91357
rect 122051 91292 122052 91356
rect 122116 91292 122117 91356
rect 122051 91291 122117 91292
rect 122974 91221 123034 94830
rect 120211 91220 120277 91221
rect 120211 91156 120212 91220
rect 120276 91156 120277 91220
rect 120211 91155 120277 91156
rect 120579 91220 120645 91221
rect 120579 91156 120580 91220
rect 120644 91156 120645 91220
rect 120579 91155 120645 91156
rect 121683 91220 121749 91221
rect 121683 91156 121684 91220
rect 121748 91156 121749 91220
rect 121683 91155 121749 91156
rect 122971 91220 123037 91221
rect 122971 91156 122972 91220
rect 123036 91156 123037 91220
rect 122971 91155 123037 91156
rect 118794 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 119414 84454
rect 118794 84134 119414 84218
rect 118794 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 119414 84134
rect 118794 48454 119414 83898
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 88954 123914 93100
rect 124078 91357 124138 94830
rect 124446 91357 124506 94830
rect 125366 94830 125444 94890
rect 125656 94890 125716 95200
rect 126472 94890 126532 95200
rect 125656 94830 125794 94890
rect 124075 91356 124141 91357
rect 124075 91292 124076 91356
rect 124140 91292 124141 91356
rect 124075 91291 124141 91292
rect 124443 91356 124509 91357
rect 124443 91292 124444 91356
rect 124508 91292 124509 91356
rect 124443 91291 124509 91292
rect 125366 91221 125426 94830
rect 125734 92445 125794 94830
rect 126470 94830 126532 94890
rect 126608 94890 126668 95200
rect 128104 94890 128164 95200
rect 129328 94890 129388 95200
rect 130688 94890 130748 95200
rect 131912 94890 131972 95200
rect 126608 94830 126714 94890
rect 128104 94830 128186 94890
rect 129328 94830 129474 94890
rect 130688 94830 130762 94890
rect 131912 94830 132050 94890
rect 126470 92445 126530 94830
rect 125731 92444 125797 92445
rect 125731 92380 125732 92444
rect 125796 92380 125797 92444
rect 125731 92379 125797 92380
rect 126467 92444 126533 92445
rect 126467 92380 126468 92444
rect 126532 92380 126533 92444
rect 126467 92379 126533 92380
rect 126654 91221 126714 94830
rect 128126 93261 128186 94830
rect 128123 93260 128189 93261
rect 128123 93196 128124 93260
rect 128188 93196 128189 93260
rect 128123 93195 128189 93196
rect 125363 91220 125429 91221
rect 125363 91156 125364 91220
rect 125428 91156 125429 91220
rect 125363 91155 125429 91156
rect 126651 91220 126717 91221
rect 126651 91156 126652 91220
rect 126716 91156 126717 91220
rect 126651 91155 126717 91156
rect 123294 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 123914 88954
rect 123294 88634 123914 88718
rect 123294 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 123914 88634
rect 123294 52954 123914 88398
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 57454 128414 93100
rect 129414 91221 129474 94830
rect 130702 92445 130762 94830
rect 130699 92444 130765 92445
rect 130699 92380 130700 92444
rect 130764 92380 130765 92444
rect 130699 92379 130765 92380
rect 131990 91629 132050 94830
rect 133136 94757 133196 95200
rect 134360 94890 134420 95200
rect 135584 94890 135644 95200
rect 151496 94890 151556 95200
rect 134360 94830 134442 94890
rect 135584 94830 135730 94890
rect 133133 94756 133199 94757
rect 133133 94692 133134 94756
rect 133198 94692 133199 94756
rect 133133 94691 133199 94692
rect 134382 93669 134442 94830
rect 134379 93668 134445 93669
rect 134379 93604 134380 93668
rect 134444 93604 134445 93668
rect 134379 93603 134445 93604
rect 131987 91628 132053 91629
rect 131987 91564 131988 91628
rect 132052 91564 132053 91628
rect 131987 91563 132053 91564
rect 129411 91220 129477 91221
rect 129411 91156 129412 91220
rect 129476 91156 129477 91220
rect 129411 91155 129477 91156
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 61954 132914 93100
rect 135670 91221 135730 94830
rect 151494 94830 151556 94890
rect 151307 94756 151373 94757
rect 151307 94692 151308 94756
rect 151372 94692 151373 94756
rect 151307 94691 151373 94692
rect 135667 91220 135733 91221
rect 135667 91156 135668 91220
rect 135732 91156 135733 91220
rect 135667 91155 135733 91156
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5146 132914 25398
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 66454 137414 93100
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6106 137414 29898
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 70954 141914 93100
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7066 141914 34398
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 75454 146414 93100
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 79954 150914 93100
rect 151310 92037 151370 94691
rect 151494 92445 151554 94830
rect 151632 94210 151692 95200
rect 151768 94757 151828 95200
rect 151904 94890 151964 95200
rect 151904 94830 152106 94890
rect 151765 94756 151831 94757
rect 151765 94692 151766 94756
rect 151830 94692 151831 94756
rect 151765 94691 151831 94692
rect 151632 94150 151738 94210
rect 151678 93669 151738 94150
rect 151675 93668 151741 93669
rect 151675 93604 151676 93668
rect 151740 93604 151741 93668
rect 151675 93603 151741 93604
rect 152046 92445 152106 94830
rect 151491 92444 151557 92445
rect 151491 92380 151492 92444
rect 151556 92380 151557 92444
rect 151491 92379 151557 92380
rect 152043 92444 152109 92445
rect 152043 92380 152044 92444
rect 152108 92380 152109 92444
rect 152043 92379 152109 92380
rect 151307 92036 151373 92037
rect 151307 91972 151308 92036
rect 151372 91972 151373 92036
rect 151307 91971 151373 91972
rect 150294 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 150914 79954
rect 150294 79634 150914 79718
rect 150294 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 150914 79634
rect 150294 43954 150914 79398
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 84454 155414 93100
rect 154794 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 155414 84454
rect 154794 84134 155414 84218
rect 154794 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 155414 84134
rect 154794 48454 155414 83898
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 88954 159914 93100
rect 159294 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 159914 88954
rect 159294 88634 159914 88718
rect 159294 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 159914 88634
rect 159294 52954 159914 88398
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 57454 164414 93100
rect 166214 78437 166274 128555
rect 166398 86733 166458 132499
rect 167502 88229 167562 134131
rect 168294 133954 168914 169398
rect 168294 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 168914 133954
rect 168294 133634 168914 133718
rect 168294 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 168914 133634
rect 167867 109172 167933 109173
rect 167867 109108 167868 109172
rect 167932 109108 167933 109172
rect 167867 109107 167933 109108
rect 167499 88228 167565 88229
rect 167499 88164 167500 88228
rect 167564 88164 167565 88228
rect 167499 88163 167565 88164
rect 167870 86869 167930 109107
rect 168294 97954 168914 133398
rect 169155 131476 169221 131477
rect 169155 131412 169156 131476
rect 169220 131412 169221 131476
rect 169155 131411 169221 131412
rect 168294 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 168914 97954
rect 168294 97634 168914 97718
rect 168294 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 168914 97634
rect 167867 86868 167933 86869
rect 167867 86804 167868 86868
rect 167932 86804 167933 86868
rect 167867 86803 167933 86804
rect 166395 86732 166461 86733
rect 166395 86668 166396 86732
rect 166460 86668 166461 86732
rect 166395 86667 166461 86668
rect 166211 78436 166277 78437
rect 166211 78372 166212 78436
rect 166276 78372 166277 78436
rect 166211 78371 166277 78372
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 61954 168914 97398
rect 169158 84149 169218 131411
rect 170262 95437 170322 296787
rect 170259 95436 170325 95437
rect 170259 95372 170260 95436
rect 170324 95372 170325 95436
rect 170259 95371 170325 95372
rect 169155 84148 169221 84149
rect 169155 84084 169156 84148
rect 169220 84084 169221 84148
rect 169155 84083 169221 84084
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5146 168914 25398
rect 170998 3365 171058 357579
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 179275 702676 179341 702677
rect 179275 702612 179276 702676
rect 179340 702612 179341 702676
rect 179275 702611 179341 702612
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 175043 350164 175109 350165
rect 175043 350100 175044 350164
rect 175108 350100 175109 350164
rect 175043 350099 175109 350100
rect 174859 330444 174925 330445
rect 174859 330380 174860 330444
rect 174924 330380 174925 330444
rect 174859 330379 174925 330380
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 171915 295356 171981 295357
rect 171915 295292 171916 295356
rect 171980 295292 171981 295356
rect 171915 295291 171981 295292
rect 171918 238509 171978 295291
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 246454 173414 281898
rect 172794 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 173414 246454
rect 172794 246134 173414 246218
rect 172794 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 173414 246134
rect 171915 238508 171981 238509
rect 171915 238444 171916 238508
rect 171980 238444 171981 238508
rect 171915 238443 171981 238444
rect 171731 238100 171797 238101
rect 171731 238036 171732 238100
rect 171796 238036 171797 238100
rect 171731 238035 171797 238036
rect 171734 92445 171794 238035
rect 172794 210454 173414 245898
rect 172794 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 173414 210454
rect 172794 210134 173414 210218
rect 172794 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 173414 210134
rect 172794 174454 173414 209898
rect 172794 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 173414 174454
rect 172794 174134 173414 174218
rect 172794 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 173414 174134
rect 172794 138454 173414 173898
rect 172794 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 173414 138454
rect 172794 138134 173414 138218
rect 172794 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 173414 138134
rect 172794 102454 173414 137898
rect 172794 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 173414 102454
rect 172794 102134 173414 102218
rect 172794 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 173414 102134
rect 171731 92444 171797 92445
rect 171731 92380 171732 92444
rect 171796 92380 171797 92444
rect 171731 92379 171797 92380
rect 172794 66454 173414 101898
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 30454 173414 65898
rect 174862 53141 174922 330379
rect 174859 53140 174925 53141
rect 174859 53076 174860 53140
rect 174924 53076 174925 53140
rect 174859 53075 174925 53076
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 170995 3364 171061 3365
rect 170995 3300 170996 3364
rect 171060 3300 171061 3364
rect 170995 3299 171061 3300
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 -6106 173414 29898
rect 175046 22677 175106 350099
rect 177067 339284 177133 339285
rect 177067 339220 177068 339284
rect 177132 339220 177133 339284
rect 177067 339219 177133 339220
rect 176515 327724 176581 327725
rect 176515 327660 176516 327724
rect 176580 327660 176581 327724
rect 176515 327659 176581 327660
rect 176331 323644 176397 323645
rect 176331 323580 176332 323644
rect 176396 323580 176397 323644
rect 176331 323579 176397 323580
rect 175043 22676 175109 22677
rect 175043 22612 175044 22676
rect 175108 22612 175109 22676
rect 175043 22611 175109 22612
rect 176334 18733 176394 323579
rect 176331 18732 176397 18733
rect 176331 18668 176332 18732
rect 176396 18668 176397 18732
rect 176331 18667 176397 18668
rect 176518 13021 176578 327659
rect 177070 61437 177130 339219
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 250954 177914 286398
rect 179278 283661 179338 702611
rect 180563 702540 180629 702541
rect 180563 702476 180564 702540
rect 180628 702476 180629 702540
rect 180563 702475 180629 702476
rect 180566 354690 180626 702475
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 357154 182414 362898
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 357154 186914 367398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 357154 191414 371898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 357154 195914 376398
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 357154 200414 380898
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 357154 204914 385398
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 357154 209414 389898
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 357154 213914 358398
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 357154 218414 362898
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 547954 222914 583398
rect 222294 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 222914 547954
rect 222294 547634 222914 547718
rect 222294 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 222914 547634
rect 222294 511954 222914 547398
rect 222294 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 222914 511954
rect 222294 511634 222914 511718
rect 222294 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 222914 511634
rect 222294 475954 222914 511398
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 357154 222914 367398
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 552454 227414 587898
rect 226794 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 227414 552454
rect 226794 552134 227414 552218
rect 226794 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 227414 552134
rect 226794 516454 227414 551898
rect 226794 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 227414 516454
rect 226794 516134 227414 516218
rect 226794 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 227414 516134
rect 226794 480454 227414 515898
rect 226794 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 227414 480454
rect 226794 480134 227414 480218
rect 226794 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 227414 480134
rect 226794 444454 227414 479898
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 357154 227414 371898
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 556954 231914 592398
rect 231294 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 231914 556954
rect 231294 556634 231914 556718
rect 231294 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 231914 556634
rect 231294 520954 231914 556398
rect 231294 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 231914 520954
rect 231294 520634 231914 520718
rect 231294 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 231914 520634
rect 231294 484954 231914 520398
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 231294 412954 231914 448398
rect 231294 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 231914 412954
rect 231294 412634 231914 412718
rect 231294 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 231914 412634
rect 231294 376954 231914 412398
rect 231294 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 231914 376954
rect 231294 376634 231914 376718
rect 231294 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 231914 376634
rect 231294 357154 231914 376398
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 357154 236414 380898
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 529954 240914 565398
rect 240294 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 240914 529954
rect 240294 529634 240914 529718
rect 240294 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 240914 529634
rect 240294 493954 240914 529398
rect 240294 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 240914 493954
rect 240294 493634 240914 493718
rect 240294 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 240914 493634
rect 240294 457954 240914 493398
rect 240294 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 240914 457954
rect 240294 457634 240914 457718
rect 240294 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 240914 457634
rect 240294 421954 240914 457398
rect 240294 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 240914 421954
rect 240294 421634 240914 421718
rect 240294 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 240914 421634
rect 240294 385954 240914 421398
rect 240294 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 240914 385954
rect 240294 385634 240914 385718
rect 240294 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 240914 385634
rect 240294 357154 240914 385398
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 534454 245414 569898
rect 244794 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 245414 534454
rect 244794 534134 245414 534218
rect 244794 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 245414 534134
rect 244794 498454 245414 533898
rect 244794 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 245414 498454
rect 244794 498134 245414 498218
rect 244794 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 245414 498134
rect 244794 462454 245414 497898
rect 244794 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 245414 462454
rect 244794 462134 245414 462218
rect 244794 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 245414 462134
rect 244794 426454 245414 461898
rect 244794 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 245414 426454
rect 244794 426134 245414 426218
rect 244794 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 245414 426134
rect 244794 390454 245414 425898
rect 244794 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 245414 390454
rect 244794 390134 245414 390218
rect 244794 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 245414 390134
rect 244794 357154 245414 389898
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 538954 249914 574398
rect 249294 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 249914 538954
rect 249294 538634 249914 538718
rect 249294 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 249914 538634
rect 249294 502954 249914 538398
rect 249294 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 249914 502954
rect 249294 502634 249914 502718
rect 249294 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 249914 502634
rect 249294 466954 249914 502398
rect 249294 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 249914 466954
rect 249294 466634 249914 466718
rect 249294 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 249914 466634
rect 249294 430954 249914 466398
rect 249294 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 249914 430954
rect 249294 430634 249914 430718
rect 249294 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 249914 430634
rect 249294 394954 249914 430398
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 249294 358954 249914 394398
rect 249294 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 249914 358954
rect 249294 358634 249914 358718
rect 249294 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 249914 358634
rect 249294 357154 249914 358398
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 357154 254414 362898
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 258294 367954 258914 403398
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 258294 357154 258914 367398
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 372454 263414 407898
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 357154 263414 371898
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 376954 267914 412398
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 357154 267914 376398
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 357154 272414 380898
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 529954 276914 565398
rect 276294 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 276914 529954
rect 276294 529634 276914 529718
rect 276294 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 276914 529634
rect 276294 493954 276914 529398
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 357154 276914 385398
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 534454 281414 569898
rect 280794 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 281414 534454
rect 280794 534134 281414 534218
rect 280794 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 281414 534134
rect 280794 498454 281414 533898
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 462454 281414 497898
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 357154 281414 389898
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 357154 285914 358398
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 357154 290414 362898
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 293907 358868 293973 358869
rect 293907 358804 293908 358868
rect 293972 358804 293973 358868
rect 293907 358803 293973 358804
rect 292803 356284 292869 356285
rect 292803 356220 292804 356284
rect 292868 356220 292869 356284
rect 292803 356219 292869 356220
rect 179830 354630 180626 354690
rect 179830 351933 179890 354630
rect 179827 351932 179893 351933
rect 179827 351868 179828 351932
rect 179892 351868 179893 351932
rect 179827 351867 179893 351868
rect 292619 347036 292685 347037
rect 292619 346972 292620 347036
rect 292684 346972 292685 347036
rect 292619 346971 292685 346972
rect 199568 331954 199888 331986
rect 199568 331718 199610 331954
rect 199846 331718 199888 331954
rect 199568 331634 199888 331718
rect 199568 331398 199610 331634
rect 199846 331398 199888 331634
rect 199568 331366 199888 331398
rect 230288 331954 230608 331986
rect 230288 331718 230330 331954
rect 230566 331718 230608 331954
rect 230288 331634 230608 331718
rect 230288 331398 230330 331634
rect 230566 331398 230608 331634
rect 230288 331366 230608 331398
rect 261008 331954 261328 331986
rect 261008 331718 261050 331954
rect 261286 331718 261328 331954
rect 261008 331634 261328 331718
rect 261008 331398 261050 331634
rect 261286 331398 261328 331634
rect 261008 331366 261328 331398
rect 184208 327454 184528 327486
rect 184208 327218 184250 327454
rect 184486 327218 184528 327454
rect 184208 327134 184528 327218
rect 184208 326898 184250 327134
rect 184486 326898 184528 327134
rect 184208 326866 184528 326898
rect 214928 327454 215248 327486
rect 214928 327218 214970 327454
rect 215206 327218 215248 327454
rect 214928 327134 215248 327218
rect 214928 326898 214970 327134
rect 215206 326898 215248 327134
rect 214928 326866 215248 326898
rect 245648 327454 245968 327486
rect 245648 327218 245690 327454
rect 245926 327218 245968 327454
rect 245648 327134 245968 327218
rect 245648 326898 245690 327134
rect 245926 326898 245968 327134
rect 245648 326866 245968 326898
rect 276368 327454 276688 327486
rect 276368 327218 276410 327454
rect 276646 327218 276688 327454
rect 276368 327134 276688 327218
rect 276368 326898 276410 327134
rect 276646 326898 276688 327134
rect 276368 326866 276688 326898
rect 199568 295954 199888 295986
rect 199568 295718 199610 295954
rect 199846 295718 199888 295954
rect 199568 295634 199888 295718
rect 199568 295398 199610 295634
rect 199846 295398 199888 295634
rect 199568 295366 199888 295398
rect 230288 295954 230608 295986
rect 230288 295718 230330 295954
rect 230566 295718 230608 295954
rect 230288 295634 230608 295718
rect 230288 295398 230330 295634
rect 230566 295398 230608 295634
rect 230288 295366 230608 295398
rect 261008 295954 261328 295986
rect 261008 295718 261050 295954
rect 261286 295718 261328 295954
rect 261008 295634 261328 295718
rect 261008 295398 261050 295634
rect 261286 295398 261328 295634
rect 261008 295366 261328 295398
rect 184208 291454 184528 291486
rect 184208 291218 184250 291454
rect 184486 291218 184528 291454
rect 184208 291134 184528 291218
rect 184208 290898 184250 291134
rect 184486 290898 184528 291134
rect 184208 290866 184528 290898
rect 214928 291454 215248 291486
rect 214928 291218 214970 291454
rect 215206 291218 215248 291454
rect 214928 291134 215248 291218
rect 214928 290898 214970 291134
rect 215206 290898 215248 291134
rect 214928 290866 215248 290898
rect 245648 291454 245968 291486
rect 245648 291218 245690 291454
rect 245926 291218 245968 291454
rect 245648 291134 245968 291218
rect 245648 290898 245690 291134
rect 245926 290898 245968 291134
rect 245648 290866 245968 290898
rect 276368 291454 276688 291486
rect 276368 291218 276410 291454
rect 276646 291218 276688 291454
rect 276368 291134 276688 291218
rect 276368 290898 276410 291134
rect 276646 290898 276688 291134
rect 276368 290866 276688 290898
rect 179275 283660 179341 283661
rect 179275 283596 179276 283660
rect 179340 283596 179341 283660
rect 179275 283595 179341 283596
rect 199568 259954 199888 259986
rect 199568 259718 199610 259954
rect 199846 259718 199888 259954
rect 199568 259634 199888 259718
rect 199568 259398 199610 259634
rect 199846 259398 199888 259634
rect 199568 259366 199888 259398
rect 230288 259954 230608 259986
rect 230288 259718 230330 259954
rect 230566 259718 230608 259954
rect 230288 259634 230608 259718
rect 230288 259398 230330 259634
rect 230566 259398 230608 259634
rect 230288 259366 230608 259398
rect 261008 259954 261328 259986
rect 261008 259718 261050 259954
rect 261286 259718 261328 259954
rect 261008 259634 261328 259718
rect 261008 259398 261050 259634
rect 261286 259398 261328 259634
rect 261008 259366 261328 259398
rect 184208 255454 184528 255486
rect 178539 255372 178605 255373
rect 178539 255308 178540 255372
rect 178604 255308 178605 255372
rect 178539 255307 178605 255308
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 214954 177914 250398
rect 178542 239053 178602 255307
rect 184208 255218 184250 255454
rect 184486 255218 184528 255454
rect 184208 255134 184528 255218
rect 184208 254898 184250 255134
rect 184486 254898 184528 255134
rect 184208 254866 184528 254898
rect 214928 255454 215248 255486
rect 214928 255218 214970 255454
rect 215206 255218 215248 255454
rect 214928 255134 215248 255218
rect 214928 254898 214970 255134
rect 215206 254898 215248 255134
rect 214928 254866 215248 254898
rect 245648 255454 245968 255486
rect 245648 255218 245690 255454
rect 245926 255218 245968 255454
rect 245648 255134 245968 255218
rect 245648 254898 245690 255134
rect 245926 254898 245968 255134
rect 245648 254866 245968 254898
rect 276368 255454 276688 255486
rect 276368 255218 276410 255454
rect 276646 255218 276688 255454
rect 276368 255134 276688 255218
rect 276368 254898 276410 255134
rect 276646 254898 276688 255134
rect 276368 254866 276688 254898
rect 179827 242996 179893 242997
rect 179827 242932 179828 242996
rect 179892 242932 179893 242996
rect 179827 242931 179893 242932
rect 178539 239052 178605 239053
rect 178539 238988 178540 239052
rect 178604 238988 178605 239052
rect 178539 238987 178605 238988
rect 177294 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 177914 214954
rect 177294 214634 177914 214718
rect 177294 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 177914 214634
rect 177294 178954 177914 214398
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 106954 177914 142398
rect 177294 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 177914 106954
rect 177294 106634 177914 106718
rect 177294 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 177914 106634
rect 177294 70954 177914 106398
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177067 61436 177133 61437
rect 177067 61372 177068 61436
rect 177132 61372 177133 61436
rect 177067 61371 177133 61372
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 176515 13020 176581 13021
rect 176515 12956 176516 13020
rect 176580 12956 176581 13020
rect 176515 12955 176581 12956
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 -7066 177914 34398
rect 179830 25669 179890 242931
rect 291699 241092 291765 241093
rect 291699 241028 291700 241092
rect 291764 241028 291765 241092
rect 291699 241027 291765 241028
rect 265571 238100 265637 238101
rect 265571 238036 265572 238100
rect 265636 238036 265637 238100
rect 265571 238035 265637 238036
rect 181794 219454 182414 238000
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 179827 25668 179893 25669
rect 179827 25604 179828 25668
rect 179892 25604 179893 25668
rect 179827 25603 179893 25604
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 223954 186914 238000
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 187954 186914 223398
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 115954 186914 151398
rect 186294 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 186914 115954
rect 186294 115634 186914 115718
rect 186294 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 186914 115634
rect 186294 79954 186914 115398
rect 186294 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 186914 79954
rect 186294 79634 186914 79718
rect 186294 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 186914 79634
rect 186294 43954 186914 79398
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 228454 191414 238000
rect 190794 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 191414 228454
rect 190794 228134 191414 228218
rect 190794 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 191414 228134
rect 190794 192454 191414 227898
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 120454 191414 155898
rect 190794 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 191414 120454
rect 190794 120134 191414 120218
rect 190794 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 191414 120134
rect 190794 84454 191414 119898
rect 190794 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 191414 84454
rect 190794 84134 191414 84218
rect 190794 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 191414 84134
rect 190794 48454 191414 83898
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 232954 195914 238000
rect 195294 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 195914 232954
rect 195294 232634 195914 232718
rect 195294 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 195914 232634
rect 195294 196954 195914 232398
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 237454 200414 238000
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 205954 204914 238000
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 210454 209414 238000
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 214954 213914 238000
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 217794 219454 218414 238000
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 178000 218414 182898
rect 222294 223954 222914 238000
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 178000 222914 187398
rect 226794 228454 227414 238000
rect 226794 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 227414 228454
rect 226794 228134 227414 228218
rect 226794 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 227414 228134
rect 226794 192454 227414 227898
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 178000 227414 191898
rect 231294 232954 231914 238000
rect 231294 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 231914 232954
rect 231294 232634 231914 232718
rect 231294 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 231914 232634
rect 231294 196954 231914 232398
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 178000 231914 196398
rect 235794 237454 236414 238000
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 178000 236414 200898
rect 249294 214954 249914 238000
rect 251219 225588 251285 225589
rect 251219 225524 251220 225588
rect 251284 225524 251285 225588
rect 251219 225523 251285 225524
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249011 180028 249077 180029
rect 249011 179964 249012 180028
rect 249076 179964 249077 180028
rect 249011 179963 249077 179964
rect 249014 177850 249074 179963
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 178000 249914 178398
rect 249014 177790 249442 177850
rect 249195 177716 249261 177717
rect 249195 177652 249196 177716
rect 249260 177652 249261 177716
rect 249195 177651 249261 177652
rect 214419 174588 214485 174589
rect 214419 174524 214420 174588
rect 214484 174524 214485 174588
rect 214419 174523 214485 174524
rect 214422 169013 214482 174523
rect 249198 174317 249258 177651
rect 249195 174316 249261 174317
rect 249195 174252 249196 174316
rect 249260 174252 249261 174316
rect 249195 174251 249261 174252
rect 249382 173773 249442 177790
rect 249379 173772 249445 173773
rect 249379 173708 249380 173772
rect 249444 173708 249445 173772
rect 249379 173707 249445 173708
rect 214419 169012 214485 169013
rect 214419 168948 214420 169012
rect 214484 168948 214485 169012
rect 214419 168947 214485 168948
rect 251035 166292 251101 166293
rect 251035 166228 251036 166292
rect 251100 166228 251101 166292
rect 251035 166227 251101 166228
rect 227874 151954 228194 151986
rect 227874 151718 227916 151954
rect 228152 151718 228194 151954
rect 227874 151634 228194 151718
rect 227874 151398 227916 151634
rect 228152 151398 228194 151634
rect 227874 151366 228194 151398
rect 237805 151954 238125 151986
rect 237805 151718 237847 151954
rect 238083 151718 238125 151954
rect 237805 151634 238125 151718
rect 237805 151398 237847 151634
rect 238083 151398 238125 151634
rect 237805 151366 238125 151398
rect 222910 147454 223230 147486
rect 222910 147218 222952 147454
rect 223188 147218 223230 147454
rect 222910 147134 223230 147218
rect 222910 146898 222952 147134
rect 223188 146898 223230 147134
rect 222910 146866 223230 146898
rect 232840 147454 233160 147486
rect 232840 147218 232882 147454
rect 233118 147218 233160 147454
rect 232840 147134 233160 147218
rect 232840 146898 232882 147134
rect 233118 146898 233160 147134
rect 232840 146866 233160 146898
rect 242771 147454 243091 147486
rect 242771 147218 242813 147454
rect 243049 147218 243091 147454
rect 242771 147134 243091 147218
rect 242771 146898 242813 147134
rect 243049 146898 243091 147134
rect 242771 146866 243091 146898
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 227874 115954 228194 115986
rect 227874 115718 227916 115954
rect 228152 115718 228194 115954
rect 227874 115634 228194 115718
rect 227874 115398 227916 115634
rect 228152 115398 228194 115634
rect 227874 115366 228194 115398
rect 237805 115954 238125 115986
rect 237805 115718 237847 115954
rect 238083 115718 238125 115954
rect 237805 115634 238125 115718
rect 237805 115398 237847 115634
rect 238083 115398 238125 115634
rect 237805 115366 238125 115398
rect 222910 111454 223230 111486
rect 222910 111218 222952 111454
rect 223188 111218 223230 111454
rect 222910 111134 223230 111218
rect 222910 110898 222952 111134
rect 223188 110898 223230 111134
rect 222910 110866 223230 110898
rect 232840 111454 233160 111486
rect 232840 111218 232882 111454
rect 233118 111218 233160 111454
rect 232840 111134 233160 111218
rect 232840 110898 232882 111134
rect 233118 110898 233160 111134
rect 232840 110866 233160 110898
rect 242771 111454 243091 111486
rect 242771 111218 242813 111454
rect 243049 111218 243091 111454
rect 242771 111134 243091 111218
rect 242771 110898 242813 111134
rect 243049 110898 243091 111134
rect 242771 110866 243091 110898
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 214419 104956 214485 104957
rect 214419 104892 214420 104956
rect 214484 104892 214485 104956
rect 214419 104891 214485 104892
rect 214422 93805 214482 104891
rect 214419 93804 214485 93805
rect 214419 93740 214420 93804
rect 214484 93740 214485 93804
rect 214419 93739 214485 93740
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 75454 218414 94000
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 79954 222914 94000
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 84454 227414 94000
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 88954 231914 94000
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 93454 236414 94000
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 61954 240914 94000
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 66454 245414 94000
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 70954 249914 94000
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 251038 3501 251098 166227
rect 251222 140861 251282 225523
rect 253794 219454 254414 238000
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 258294 223954 258914 238000
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 255267 206276 255333 206277
rect 255267 206212 255268 206276
rect 255332 206212 255333 206276
rect 255267 206211 255333 206212
rect 254531 188324 254597 188325
rect 254531 188260 254532 188324
rect 254596 188260 254597 188324
rect 254531 188259 254597 188260
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 252507 176084 252573 176085
rect 252507 176020 252508 176084
rect 252572 176020 252573 176084
rect 252507 176019 252573 176020
rect 251955 149700 252021 149701
rect 251955 149636 251956 149700
rect 252020 149636 252021 149700
rect 251955 149635 252021 149636
rect 251219 140860 251285 140861
rect 251219 140796 251220 140860
rect 251284 140796 251285 140860
rect 251219 140795 251285 140796
rect 251771 131748 251837 131749
rect 251771 131684 251772 131748
rect 251836 131684 251837 131748
rect 251771 131683 251837 131684
rect 251774 96661 251834 131683
rect 251958 111213 252018 149635
rect 252510 147933 252570 176019
rect 252507 147932 252573 147933
rect 252507 147868 252508 147932
rect 252572 147868 252573 147932
rect 252507 147867 252573 147868
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 254534 146981 254594 188259
rect 254531 146980 254597 146981
rect 254531 146916 254532 146980
rect 254596 146916 254597 146980
rect 254531 146915 254597 146916
rect 253427 141404 253493 141405
rect 253427 141340 253428 141404
rect 253492 141340 253493 141404
rect 253427 141339 253493 141340
rect 253430 122850 253490 141339
rect 253062 122790 253490 122850
rect 251955 111212 252021 111213
rect 251955 111148 251956 111212
rect 252020 111148 252021 111212
rect 251955 111147 252021 111148
rect 253062 101829 253122 122790
rect 253794 111454 254414 146898
rect 255270 139501 255330 206211
rect 258294 187954 258914 223398
rect 262794 228454 263414 238000
rect 262794 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 263414 228454
rect 262794 228134 263414 228218
rect 262794 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 263414 228134
rect 260971 215932 261037 215933
rect 260971 215868 260972 215932
rect 261036 215868 261037 215932
rect 260971 215867 261037 215868
rect 259683 192676 259749 192677
rect 259683 192612 259684 192676
rect 259748 192612 259749 192676
rect 259683 192611 259749 192612
rect 259499 191044 259565 191045
rect 259499 190980 259500 191044
rect 259564 190980 259565 191044
rect 259499 190979 259565 190980
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 256923 185604 256989 185605
rect 256923 185540 256924 185604
rect 256988 185540 256989 185604
rect 256923 185539 256989 185540
rect 255451 181524 255517 181525
rect 255451 181460 255452 181524
rect 255516 181460 255517 181524
rect 255451 181459 255517 181460
rect 255454 158269 255514 181459
rect 256739 180164 256805 180165
rect 256739 180100 256740 180164
rect 256804 180100 256805 180164
rect 256739 180099 256805 180100
rect 256742 161125 256802 180099
rect 256926 168605 256986 185539
rect 257843 177308 257909 177309
rect 257843 177244 257844 177308
rect 257908 177244 257909 177308
rect 257843 177243 257909 177244
rect 256923 168604 256989 168605
rect 256923 168540 256924 168604
rect 256988 168540 256989 168604
rect 256923 168539 256989 168540
rect 256739 161124 256805 161125
rect 256739 161060 256740 161124
rect 256804 161060 256805 161124
rect 256739 161059 256805 161060
rect 255451 158268 255517 158269
rect 255451 158204 255452 158268
rect 255516 158204 255517 158268
rect 255451 158203 255517 158204
rect 257846 152965 257906 177243
rect 257843 152964 257909 152965
rect 257843 152900 257844 152964
rect 257908 152900 257909 152964
rect 257843 152899 257909 152900
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 255267 139500 255333 139501
rect 255267 139436 255268 139500
rect 255332 139436 255333 139500
rect 255267 139435 255333 139436
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253059 101828 253125 101829
rect 253059 101764 253060 101828
rect 253124 101764 253125 101828
rect 253059 101763 253125 101764
rect 251771 96660 251837 96661
rect 251771 96596 251772 96660
rect 251836 96596 251837 96660
rect 251771 96595 251837 96596
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 251035 3500 251101 3501
rect 251035 3436 251036 3500
rect 251100 3436 251101 3500
rect 251035 3435 251101 3436
rect 253794 3454 254414 38898
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 115954 258914 151398
rect 259502 138549 259562 190979
rect 259686 142221 259746 192611
rect 260974 190470 261034 215867
rect 260790 190410 261034 190470
rect 262794 192454 263414 227898
rect 265019 213212 265085 213213
rect 265019 213148 265020 213212
rect 265084 213148 265085 213212
rect 265019 213147 265085 213148
rect 263547 206412 263613 206413
rect 263547 206348 263548 206412
rect 263612 206348 263613 206412
rect 263547 206347 263613 206348
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 260790 161533 260850 190410
rect 260971 189684 261037 189685
rect 260971 189620 260972 189684
rect 261036 189620 261037 189684
rect 260971 189619 261037 189620
rect 260787 161532 260853 161533
rect 260787 161468 260788 161532
rect 260852 161468 260853 161532
rect 260787 161467 260853 161468
rect 259683 142220 259749 142221
rect 259683 142156 259684 142220
rect 259748 142156 259749 142220
rect 259683 142155 259749 142156
rect 260974 141269 261034 189619
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 260971 141268 261037 141269
rect 260971 141204 260972 141268
rect 261036 141204 261037 141268
rect 260971 141203 261037 141204
rect 259499 138548 259565 138549
rect 259499 138484 259500 138548
rect 259564 138484 259565 138548
rect 259499 138483 259565 138484
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 120454 263414 155898
rect 263550 144669 263610 206347
rect 264099 176764 264165 176765
rect 264099 176700 264100 176764
rect 264164 176700 264165 176764
rect 264099 176699 264165 176700
rect 263547 144668 263613 144669
rect 263547 144604 263548 144668
rect 263612 144604 263613 144668
rect 263547 144603 263613 144604
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 264102 97069 264162 176699
rect 265022 162213 265082 213147
rect 265019 162212 265085 162213
rect 265019 162148 265020 162212
rect 265084 162148 265085 162212
rect 265019 162147 265085 162148
rect 264099 97068 264165 97069
rect 264099 97004 264100 97068
rect 264164 97004 264165 97068
rect 264099 97003 264165 97004
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 265574 47565 265634 238035
rect 267294 232954 267914 238000
rect 267294 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 267914 232954
rect 267294 232634 267914 232718
rect 267294 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 267914 232634
rect 267294 196954 267914 232398
rect 271794 237454 272414 238000
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 269619 229804 269685 229805
rect 269619 229740 269620 229804
rect 269684 229740 269685 229804
rect 269619 229739 269685 229740
rect 269067 210492 269133 210493
rect 269067 210428 269068 210492
rect 269132 210428 269133 210492
rect 269067 210427 269133 210428
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 266307 184380 266373 184381
rect 266307 184316 266308 184380
rect 266372 184316 266373 184380
rect 266307 184315 266373 184316
rect 266310 163029 266370 184315
rect 266307 163028 266373 163029
rect 266307 162964 266308 163028
rect 266372 162964 266373 163028
rect 266307 162963 266373 162964
rect 267294 160954 267914 196398
rect 269070 163165 269130 210427
rect 269067 163164 269133 163165
rect 269067 163100 269068 163164
rect 269132 163100 269133 163164
rect 269067 163099 269133 163100
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 269622 94485 269682 229739
rect 271091 228308 271157 228309
rect 271091 228244 271092 228308
rect 271156 228244 271157 228308
rect 271091 228243 271157 228244
rect 270539 199340 270605 199341
rect 270539 199276 270540 199340
rect 270604 199276 270605 199340
rect 270539 199275 270605 199276
rect 270542 139773 270602 199275
rect 270539 139772 270605 139773
rect 270539 139708 270540 139772
rect 270604 139708 270605 139772
rect 270539 139707 270605 139708
rect 269619 94484 269685 94485
rect 269619 94420 269620 94484
rect 269684 94420 269685 94484
rect 269619 94419 269685 94420
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 265571 47564 265637 47565
rect 265571 47500 265572 47564
rect 265636 47500 265637 47564
rect 265571 47499 265637 47500
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 271094 3365 271154 228243
rect 271794 201454 272414 236898
rect 273851 226948 273917 226949
rect 273851 226884 273852 226948
rect 273916 226884 273917 226948
rect 273851 226883 273917 226884
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 273854 138685 273914 226883
rect 276294 205954 276914 238000
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 275139 162076 275205 162077
rect 275139 162012 275140 162076
rect 275204 162012 275205 162076
rect 275139 162011 275205 162012
rect 273851 138684 273917 138685
rect 273851 138620 273852 138684
rect 273916 138620 273917 138684
rect 273851 138619 273917 138620
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 275142 85645 275202 162011
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 275139 85644 275205 85645
rect 275139 85580 275140 85644
rect 275204 85580 275205 85644
rect 275139 85579 275205 85580
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271091 3364 271157 3365
rect 271091 3300 271092 3364
rect 271156 3300 271157 3364
rect 271091 3299 271157 3300
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 210454 281414 238000
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 285294 214954 285914 238000
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 282131 113524 282197 113525
rect 282131 113460 282132 113524
rect 282196 113460 282197 113524
rect 282131 113459 282197 113460
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 282134 18597 282194 113459
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 282131 18596 282197 18597
rect 282131 18532 282132 18596
rect 282196 18532 282197 18596
rect 282131 18531 282197 18532
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 219454 290414 238000
rect 291702 226949 291762 241027
rect 291699 226948 291765 226949
rect 291699 226884 291700 226948
rect 291764 226884 291765 226948
rect 291699 226883 291765 226884
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 292622 80749 292682 346971
rect 292619 80748 292685 80749
rect 292619 80684 292620 80748
rect 292684 80684 292685 80748
rect 292619 80683 292685 80684
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 292806 3501 292866 356219
rect 293910 345541 293970 358803
rect 294294 357154 294914 367398
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 552454 299414 587898
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 298794 516454 299414 551898
rect 298794 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 299414 516454
rect 298794 516134 299414 516218
rect 298794 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 299414 516134
rect 298794 480454 299414 515898
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 556954 303914 592398
rect 303294 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 303914 556954
rect 303294 556634 303914 556718
rect 303294 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 303914 556634
rect 303294 520954 303914 556398
rect 303294 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 303914 520954
rect 303294 520634 303914 520718
rect 303294 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 303914 520634
rect 303294 484954 303914 520398
rect 303294 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 303914 484954
rect 303294 484634 303914 484718
rect 299979 484532 300045 484533
rect 299979 484468 299980 484532
rect 300044 484468 300045 484532
rect 299979 484467 300045 484468
rect 298794 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 299414 480454
rect 298794 480134 299414 480218
rect 298794 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 299414 480134
rect 298794 444454 299414 479898
rect 298794 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 299414 444454
rect 298794 444134 299414 444218
rect 298794 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 299414 444134
rect 298794 408454 299414 443898
rect 298794 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 299414 408454
rect 298794 408134 299414 408218
rect 298794 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 299414 408134
rect 298794 372454 299414 407898
rect 298794 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 299414 372454
rect 298794 372134 299414 372218
rect 298794 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 299414 372134
rect 297219 357644 297285 357645
rect 297219 357580 297220 357644
rect 297284 357580 297285 357644
rect 297219 357579 297285 357580
rect 295379 349620 295445 349621
rect 295379 349556 295380 349620
rect 295444 349556 295445 349620
rect 295379 349555 295445 349556
rect 293907 345540 293973 345541
rect 293907 345476 293908 345540
rect 293972 345476 293973 345540
rect 293907 345475 293973 345476
rect 293907 281620 293973 281621
rect 293907 281556 293908 281620
rect 293972 281556 293973 281620
rect 293907 281555 293973 281556
rect 293910 238781 293970 281555
rect 293907 238780 293973 238781
rect 293907 238716 293908 238780
rect 293972 238716 293973 238780
rect 293907 238715 293973 238716
rect 294294 223954 294914 238000
rect 295382 235925 295442 349555
rect 295379 235924 295445 235925
rect 295379 235860 295380 235924
rect 295444 235860 295445 235924
rect 295379 235859 295445 235860
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 295931 131476 295997 131477
rect 295931 131412 295932 131476
rect 295996 131412 295997 131476
rect 295931 131411 295997 131412
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 295934 55861 295994 131411
rect 297222 73813 297282 357579
rect 298794 336454 299414 371898
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 298794 300454 299414 335898
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 228454 299414 263898
rect 299611 247076 299677 247077
rect 299611 247012 299612 247076
rect 299676 247012 299677 247076
rect 299611 247011 299677 247012
rect 299614 230485 299674 247011
rect 299982 238509 300042 484467
rect 303294 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 303914 484634
rect 303294 448954 303914 484398
rect 303294 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 303914 448954
rect 303294 448634 303914 448718
rect 303294 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 303914 448634
rect 303294 412954 303914 448398
rect 303294 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 303914 412954
rect 303294 412634 303914 412718
rect 303294 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 303914 412634
rect 303294 376954 303914 412398
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 301451 356148 301517 356149
rect 301451 356084 301452 356148
rect 301516 356084 301517 356148
rect 301451 356083 301517 356084
rect 299979 238508 300045 238509
rect 299979 238444 299980 238508
rect 300044 238444 300045 238508
rect 299979 238443 300045 238444
rect 299611 230484 299677 230485
rect 299611 230420 299612 230484
rect 299676 230420 299677 230484
rect 299611 230419 299677 230420
rect 298794 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 299414 228454
rect 298794 228134 299414 228218
rect 298794 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 299414 228134
rect 298794 192454 299414 227898
rect 298794 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 299414 192454
rect 298794 192134 299414 192218
rect 298794 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 299414 192134
rect 298794 156454 299414 191898
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 300163 126444 300229 126445
rect 300163 126380 300164 126444
rect 300228 126380 300229 126444
rect 300163 126379 300229 126380
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 299979 117468 300045 117469
rect 299979 117404 299980 117468
rect 300044 117404 300045 117468
rect 299979 117403 300045 117404
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 297219 73812 297285 73813
rect 297219 73748 297220 73812
rect 297284 73748 297285 73812
rect 297219 73747 297285 73748
rect 295931 55860 295997 55861
rect 295931 55796 295932 55860
rect 295996 55796 295997 55860
rect 295931 55795 295997 55796
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 292803 3500 292869 3501
rect 292803 3436 292804 3500
rect 292868 3436 292869 3500
rect 292803 3435 292869 3436
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 299982 4861 300042 117403
rect 300166 46205 300226 126379
rect 300163 46204 300229 46205
rect 300163 46140 300164 46204
rect 300228 46140 300229 46204
rect 300163 46139 300229 46140
rect 299979 4860 300045 4861
rect 299979 4796 299980 4860
rect 300044 4796 300045 4860
rect 299979 4795 300045 4796
rect 301454 4045 301514 356083
rect 303294 340954 303914 376398
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 303294 304954 303914 340398
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 232954 303914 268398
rect 303294 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 303914 232954
rect 303294 232634 303914 232718
rect 303294 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 303914 232634
rect 303294 196954 303914 232398
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 306235 189684 306301 189685
rect 306235 189620 306236 189684
rect 306300 189620 306301 189684
rect 306235 189619 306301 189620
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 303294 124954 303914 160398
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 304211 119100 304277 119101
rect 304211 119036 304212 119100
rect 304276 119036 304277 119100
rect 304211 119035 304277 119036
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 304214 25533 304274 119035
rect 305499 118692 305565 118693
rect 305499 118628 305500 118692
rect 305564 118628 305565 118692
rect 305499 118627 305565 118628
rect 305502 44845 305562 118627
rect 306238 100061 306298 189619
rect 307794 178000 308414 200898
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 529954 312914 565398
rect 312294 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 312914 529954
rect 312294 529634 312914 529718
rect 312294 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 312914 529634
rect 312294 493954 312914 529398
rect 312294 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 312914 493954
rect 312294 493634 312914 493718
rect 312294 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 312914 493634
rect 312294 457954 312914 493398
rect 312294 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 312914 457954
rect 312294 457634 312914 457718
rect 312294 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 312914 457634
rect 312294 421954 312914 457398
rect 312294 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 312914 421954
rect 312294 421634 312914 421718
rect 312294 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 312914 421634
rect 312294 385954 312914 421398
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 313954 312914 349398
rect 312294 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 312914 313954
rect 312294 313634 312914 313718
rect 312294 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 312914 313634
rect 312294 277954 312914 313398
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 241954 312914 277398
rect 312294 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 312914 241954
rect 312294 241634 312914 241718
rect 312294 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 312914 241634
rect 312294 205954 312914 241398
rect 312294 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 312914 205954
rect 312294 205634 312914 205718
rect 312294 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 312914 205634
rect 312294 178000 312914 205398
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 534454 317414 569898
rect 316794 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 317414 534454
rect 316794 534134 317414 534218
rect 316794 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 317414 534134
rect 316794 498454 317414 533898
rect 316794 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 317414 498454
rect 316794 498134 317414 498218
rect 316794 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 317414 498134
rect 316794 462454 317414 497898
rect 316794 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 317414 462454
rect 316794 462134 317414 462218
rect 316794 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 317414 462134
rect 316794 426454 317414 461898
rect 316794 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 317414 426454
rect 316794 426134 317414 426218
rect 316794 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 317414 426134
rect 316794 390454 317414 425898
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 318454 317414 353898
rect 316794 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 317414 318454
rect 316794 318134 317414 318218
rect 316794 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 317414 318134
rect 316794 282454 317414 317898
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 246454 317414 281898
rect 316794 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 317414 246454
rect 316794 246134 317414 246218
rect 316794 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 317414 246134
rect 316794 210454 317414 245898
rect 316794 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 317414 210454
rect 316794 210134 317414 210218
rect 316794 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 317414 210134
rect 316794 178000 317414 209898
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 538954 321914 574398
rect 321294 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 321914 538954
rect 321294 538634 321914 538718
rect 321294 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 321914 538634
rect 321294 502954 321914 538398
rect 321294 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 321914 502954
rect 321294 502634 321914 502718
rect 321294 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 321914 502634
rect 321294 466954 321914 502398
rect 321294 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 321914 466954
rect 321294 466634 321914 466718
rect 321294 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 321914 466634
rect 321294 430954 321914 466398
rect 321294 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 321914 430954
rect 321294 430634 321914 430718
rect 321294 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 321914 430634
rect 321294 394954 321914 430398
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 322954 321914 358398
rect 321294 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 321914 322954
rect 321294 322634 321914 322718
rect 321294 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 321914 322634
rect 321294 286954 321914 322398
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 214954 321914 250398
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 322059 233884 322125 233885
rect 322059 233820 322060 233884
rect 322124 233820 322125 233884
rect 322059 233819 322125 233820
rect 321294 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 321914 214954
rect 321294 214634 321914 214718
rect 321294 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 321914 214634
rect 320403 186964 320469 186965
rect 320403 186900 320404 186964
rect 320468 186900 320469 186964
rect 320403 186899 320469 186900
rect 320219 176764 320285 176765
rect 320219 176700 320220 176764
rect 320284 176700 320285 176764
rect 320219 176699 320285 176700
rect 320222 171150 320282 176699
rect 320406 175810 320466 186899
rect 321294 178954 321914 214398
rect 321294 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 321914 178954
rect 321294 178634 321914 178718
rect 321294 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 321914 178634
rect 321294 178000 321914 178398
rect 321507 176220 321573 176221
rect 321507 176156 321508 176220
rect 321572 176156 321573 176220
rect 321507 176155 321573 176156
rect 320406 175750 321386 175810
rect 321326 171461 321386 175750
rect 321510 172141 321570 176155
rect 321507 172140 321573 172141
rect 321507 172076 321508 172140
rect 321572 172076 321573 172140
rect 321507 172075 321573 172076
rect 321323 171460 321389 171461
rect 321323 171396 321324 171460
rect 321388 171396 321389 171460
rect 321323 171395 321389 171396
rect 320222 171090 321386 171150
rect 321326 170645 321386 171090
rect 321323 170644 321389 170645
rect 321323 170580 321324 170644
rect 321388 170580 321389 170644
rect 321323 170579 321389 170580
rect 307155 157452 307221 157453
rect 307155 157388 307156 157452
rect 307220 157388 307221 157452
rect 307155 157387 307221 157388
rect 306971 154868 307037 154869
rect 306971 154804 306972 154868
rect 307036 154804 307037 154868
rect 306971 154803 307037 154804
rect 306974 144125 307034 154803
rect 307158 148341 307218 157387
rect 314208 151954 314528 151986
rect 314208 151718 314250 151954
rect 314486 151718 314528 151954
rect 314208 151634 314528 151718
rect 314208 151398 314250 151634
rect 314486 151398 314528 151634
rect 314208 151366 314528 151398
rect 317472 151954 317792 151986
rect 317472 151718 317514 151954
rect 317750 151718 317792 151954
rect 317472 151634 317792 151718
rect 317472 151398 317514 151634
rect 317750 151398 317792 151634
rect 317472 151366 317792 151398
rect 307155 148340 307221 148341
rect 307155 148276 307156 148340
rect 307220 148276 307221 148340
rect 307155 148275 307221 148276
rect 312576 147454 312896 147486
rect 312576 147218 312618 147454
rect 312854 147218 312896 147454
rect 312576 147134 312896 147218
rect 312576 146898 312618 147134
rect 312854 146898 312896 147134
rect 312576 146866 312896 146898
rect 315840 147454 316160 147486
rect 315840 147218 315882 147454
rect 316118 147218 316160 147454
rect 315840 147134 316160 147218
rect 315840 146898 315882 147134
rect 316118 146898 316160 147134
rect 315840 146866 316160 146898
rect 319104 147454 319424 147486
rect 319104 147218 319146 147454
rect 319382 147218 319424 147454
rect 319104 147134 319424 147218
rect 319104 146898 319146 147134
rect 319382 146898 319424 147134
rect 319104 146866 319424 146898
rect 322062 144669 322122 233819
rect 325794 219454 326414 254898
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 511954 330914 547398
rect 330294 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 330914 511954
rect 330294 511634 330914 511718
rect 330294 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 330914 511634
rect 330294 475954 330914 511398
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 330294 439954 330914 475398
rect 330294 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 330914 439954
rect 330294 439634 330914 439718
rect 330294 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 330914 439634
rect 330294 403954 330914 439398
rect 330294 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 330914 403954
rect 330294 403634 330914 403718
rect 330294 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 330914 403634
rect 330294 367954 330914 403398
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 331954 330914 367398
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 552454 335414 587898
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 516454 335414 551898
rect 334794 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 335414 516454
rect 334794 516134 335414 516218
rect 334794 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 335414 516134
rect 334794 480454 335414 515898
rect 334794 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 335414 480454
rect 334794 480134 335414 480218
rect 334794 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 335414 480134
rect 334794 444454 335414 479898
rect 334794 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 335414 444454
rect 334794 444134 335414 444218
rect 334794 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 335414 444134
rect 334794 408454 335414 443898
rect 334794 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 335414 408454
rect 334794 408134 335414 408218
rect 334794 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 335414 408134
rect 334794 372454 335414 407898
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 332547 361724 332613 361725
rect 332547 361660 332548 361724
rect 332612 361660 332613 361724
rect 332547 361659 332613 361660
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 328499 237964 328565 237965
rect 328499 237900 328500 237964
rect 328564 237900 328565 237964
rect 328499 237899 328565 237900
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 327211 214572 327277 214573
rect 327211 214508 327212 214572
rect 327276 214508 327277 214572
rect 327211 214507 327277 214508
rect 327027 197980 327093 197981
rect 327027 197916 327028 197980
rect 327092 197916 327093 197980
rect 327027 197915 327093 197916
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 322059 144668 322125 144669
rect 322059 144604 322060 144668
rect 322124 144604 322125 144668
rect 322059 144603 322125 144604
rect 306971 144124 307037 144125
rect 306971 144060 306972 144124
rect 307036 144060 307037 144124
rect 306971 144059 307037 144060
rect 307155 130660 307221 130661
rect 307155 130596 307156 130660
rect 307220 130596 307221 130660
rect 307155 130595 307221 130596
rect 306971 114068 307037 114069
rect 306971 114004 306972 114068
rect 307036 114004 307037 114068
rect 306971 114003 307037 114004
rect 306235 100060 306301 100061
rect 306235 99996 306236 100060
rect 306300 99996 306301 100060
rect 306235 99995 306301 99996
rect 305499 44844 305565 44845
rect 305499 44780 305500 44844
rect 305564 44780 305565 44844
rect 305499 44779 305565 44780
rect 304211 25532 304277 25533
rect 304211 25468 304212 25532
rect 304276 25468 304277 25532
rect 304211 25467 304277 25468
rect 306974 17237 307034 114003
rect 307158 62797 307218 130595
rect 314208 115954 314528 115986
rect 314208 115718 314250 115954
rect 314486 115718 314528 115954
rect 314208 115634 314528 115718
rect 314208 115398 314250 115634
rect 314486 115398 314528 115634
rect 314208 115366 314528 115398
rect 317472 115954 317792 115986
rect 317472 115718 317514 115954
rect 317750 115718 317792 115954
rect 317472 115634 317792 115718
rect 317472 115398 317514 115634
rect 317750 115398 317792 115634
rect 317472 115366 317792 115398
rect 312576 111454 312896 111486
rect 312576 111218 312618 111454
rect 312854 111218 312896 111454
rect 312576 111134 312896 111218
rect 312576 110898 312618 111134
rect 312854 110898 312896 111134
rect 312576 110866 312896 110898
rect 315840 111454 316160 111486
rect 315840 111218 315882 111454
rect 316118 111218 316160 111454
rect 315840 111134 316160 111218
rect 315840 110898 315882 111134
rect 316118 110898 316160 111134
rect 315840 110866 316160 110898
rect 319104 111454 319424 111486
rect 319104 111218 319146 111454
rect 319382 111218 319424 111454
rect 319104 111134 319424 111218
rect 319104 110898 319146 111134
rect 319382 110898 319424 111134
rect 319104 110866 319424 110898
rect 325794 111454 326414 146898
rect 327030 121685 327090 197915
rect 327214 145485 327274 214507
rect 327211 145484 327277 145485
rect 327211 145420 327212 145484
rect 327276 145420 327277 145484
rect 327211 145419 327277 145420
rect 328502 125629 328562 237899
rect 330294 223954 330914 259398
rect 330294 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 330914 223954
rect 330294 223634 330914 223718
rect 330294 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 330914 223634
rect 328683 210356 328749 210357
rect 328683 210292 328684 210356
rect 328748 210292 328749 210356
rect 328683 210291 328749 210292
rect 328499 125628 328565 125629
rect 328499 125564 328500 125628
rect 328564 125564 328565 125628
rect 328499 125563 328565 125564
rect 327027 121684 327093 121685
rect 327027 121620 327028 121684
rect 327092 121620 327093 121684
rect 327027 121619 327093 121620
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 309179 99924 309245 99925
rect 309179 99860 309180 99924
rect 309244 99860 309245 99924
rect 309179 99859 309245 99860
rect 307794 93454 308414 94000
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307155 62796 307221 62797
rect 307155 62732 307156 62796
rect 307220 62732 307221 62796
rect 307155 62731 307221 62732
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 306971 17236 307037 17237
rect 306971 17172 306972 17236
rect 307036 17172 307037 17236
rect 306971 17171 307037 17172
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 301451 4044 301517 4045
rect 301451 3980 301452 4044
rect 301516 3980 301517 4044
rect 301451 3979 301517 3980
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 -4186 308414 20898
rect 309182 3501 309242 99859
rect 324267 98564 324333 98565
rect 324267 98500 324268 98564
rect 324332 98500 324333 98564
rect 324267 98499 324333 98500
rect 312294 61954 312914 94000
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 309179 3500 309245 3501
rect 309179 3436 309180 3500
rect 309244 3436 309245 3500
rect 309179 3435 309245 3436
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 66454 317414 94000
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 70954 321914 94000
rect 324270 78573 324330 98499
rect 324267 78572 324333 78573
rect 324267 78508 324268 78572
rect 324332 78508 324333 78572
rect 324267 78507 324333 78508
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 75454 326414 110898
rect 328686 106453 328746 210291
rect 329787 192540 329853 192541
rect 329787 192476 329788 192540
rect 329852 192476 329853 192540
rect 329787 192475 329853 192476
rect 329790 123317 329850 192475
rect 330294 187954 330914 223398
rect 331259 204916 331325 204917
rect 331259 204852 331260 204916
rect 331324 204852 331325 204916
rect 331259 204851 331325 204852
rect 330294 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 330914 187954
rect 330294 187634 330914 187718
rect 330294 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 330914 187634
rect 330294 151954 330914 187398
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 329787 123316 329853 123317
rect 329787 123252 329788 123316
rect 329852 123252 329853 123316
rect 329787 123251 329853 123252
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 328683 106452 328749 106453
rect 328683 106388 328684 106452
rect 328748 106388 328749 106452
rect 328683 106387 328749 106388
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 331262 6357 331322 204851
rect 331443 177444 331509 177445
rect 331443 177380 331444 177444
rect 331508 177380 331509 177444
rect 331443 177379 331509 177380
rect 331446 134197 331506 177379
rect 331443 134196 331509 134197
rect 331443 134132 331444 134196
rect 331508 134132 331509 134196
rect 331443 134131 331509 134132
rect 331259 6356 331325 6357
rect 331259 6292 331260 6356
rect 331324 6292 331325 6356
rect 331259 6291 331325 6292
rect 332550 6221 332610 361659
rect 334794 336454 335414 371898
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 300454 335414 335898
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 228454 335414 263898
rect 334794 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 335414 228454
rect 334794 228134 335414 228218
rect 334794 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 335414 228134
rect 334794 192454 335414 227898
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 556954 339914 592398
rect 339294 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 339914 556954
rect 339294 556634 339914 556718
rect 339294 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 339914 556634
rect 339294 520954 339914 556398
rect 339294 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 339914 520954
rect 339294 520634 339914 520718
rect 339294 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 339914 520634
rect 339294 484954 339914 520398
rect 339294 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 339914 484954
rect 339294 484634 339914 484718
rect 339294 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 339914 484634
rect 339294 448954 339914 484398
rect 339294 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 339914 448954
rect 339294 448634 339914 448718
rect 339294 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 339914 448634
rect 339294 412954 339914 448398
rect 339294 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 339914 412954
rect 339294 412634 339914 412718
rect 339294 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 339914 412634
rect 339294 376954 339914 412398
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 339294 340954 339914 376398
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 342299 363084 342365 363085
rect 342299 363020 342300 363084
rect 342364 363020 342365 363084
rect 342299 363019 342365 363020
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 304954 339914 340398
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 232954 339914 268398
rect 339294 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 339914 232954
rect 339294 232634 339914 232718
rect 339294 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 339914 232634
rect 336963 221508 337029 221509
rect 336963 221444 336964 221508
rect 337028 221444 337029 221508
rect 336963 221443 337029 221444
rect 335859 211988 335925 211989
rect 335859 211924 335860 211988
rect 335924 211924 335925 211988
rect 335859 211923 335925 211924
rect 335675 211852 335741 211853
rect 335675 211850 335676 211852
rect 334794 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 335414 192454
rect 334794 192134 335414 192218
rect 334794 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 335414 192134
rect 332731 182884 332797 182885
rect 332731 182820 332732 182884
rect 332796 182820 332797 182884
rect 332731 182819 332797 182820
rect 332734 133925 332794 182819
rect 334019 178804 334085 178805
rect 334019 178740 334020 178804
rect 334084 178740 334085 178804
rect 334019 178739 334085 178740
rect 334022 138141 334082 178739
rect 334794 156454 335414 191898
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334019 138140 334085 138141
rect 334019 138076 334020 138140
rect 334084 138076 334085 138140
rect 334019 138075 334085 138076
rect 332731 133924 332797 133925
rect 332731 133860 332732 133924
rect 332796 133860 332797 133924
rect 332731 133859 332797 133860
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 335494 211790 335676 211850
rect 335494 110530 335554 211790
rect 335675 211788 335676 211790
rect 335740 211788 335741 211852
rect 335675 211787 335741 211788
rect 335862 200130 335922 211923
rect 335678 200070 335922 200130
rect 335678 145621 335738 200070
rect 336779 177308 336845 177309
rect 336779 177244 336780 177308
rect 336844 177244 336845 177308
rect 336779 177243 336845 177244
rect 335675 145620 335741 145621
rect 335675 145556 335676 145620
rect 335740 145556 335741 145620
rect 335675 145555 335741 145556
rect 335675 110532 335741 110533
rect 335675 110530 335676 110532
rect 335494 110470 335676 110530
rect 335675 110468 335676 110470
rect 335740 110468 335741 110532
rect 335675 110467 335741 110468
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 332547 6220 332613 6221
rect 332547 6156 332548 6220
rect 332612 6156 332613 6220
rect 332547 6155 332613 6156
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 -2266 335414 11898
rect 336782 3365 336842 177243
rect 336966 109173 337026 221443
rect 339294 196954 339914 232398
rect 340827 200700 340893 200701
rect 340827 200636 340828 200700
rect 340892 200636 340893 200700
rect 340827 200635 340893 200636
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 339294 160954 339914 196398
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 339294 124954 339914 160398
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 336963 109172 337029 109173
rect 336963 109108 336964 109172
rect 337028 109108 337029 109172
rect 336963 109107 337029 109108
rect 339294 88954 339914 124398
rect 340830 114613 340890 200635
rect 340827 114612 340893 114613
rect 340827 114548 340828 114612
rect 340892 114548 340893 114612
rect 340827 114547 340893 114548
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 336779 3364 336845 3365
rect 336779 3300 336780 3364
rect 336844 3300 336845 3364
rect 336779 3299 336845 3300
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 -3226 339914 16398
rect 342302 3501 342362 363019
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 529954 348914 565398
rect 348294 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 348914 529954
rect 348294 529634 348914 529718
rect 348294 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 348914 529634
rect 348294 493954 348914 529398
rect 348294 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 348914 493954
rect 348294 493634 348914 493718
rect 348294 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 348914 493634
rect 348294 457954 348914 493398
rect 348294 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 348914 457954
rect 348294 457634 348914 457718
rect 348294 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 348914 457634
rect 348294 421954 348914 457398
rect 348294 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 348914 421954
rect 348294 421634 348914 421718
rect 348294 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 348914 421634
rect 348294 385954 348914 421398
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 313954 348914 349398
rect 348294 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 348914 313954
rect 348294 313634 348914 313718
rect 348294 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 348914 313634
rect 348294 277954 348914 313398
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 241954 348914 277398
rect 348294 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 348914 241954
rect 348294 241634 348914 241718
rect 348294 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 348914 241634
rect 346347 210628 346413 210629
rect 346347 210564 346348 210628
rect 346412 210564 346413 210628
rect 346347 210563 346413 210564
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 346350 102237 346410 210563
rect 348294 205954 348914 241398
rect 348294 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 348914 205954
rect 348294 205634 348914 205718
rect 348294 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 348914 205634
rect 348294 169954 348914 205398
rect 348294 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 348914 169954
rect 348294 169634 348914 169718
rect 348294 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 348914 169634
rect 348294 133954 348914 169398
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 346347 102236 346413 102237
rect 346347 102172 346348 102236
rect 346412 102172 346413 102236
rect 346347 102171 346413 102172
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 342299 3500 342365 3501
rect 342299 3436 342300 3500
rect 342364 3436 342365 3500
rect 342299 3435 342365 3436
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 534454 353414 569898
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 352794 498454 353414 533898
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 426454 353414 461898
rect 352794 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 353414 426454
rect 352794 426134 353414 426218
rect 352794 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 353414 426134
rect 352794 390454 353414 425898
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 210454 353414 245898
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 138454 353414 173898
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 538954 357914 574398
rect 357294 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 357914 538954
rect 357294 538634 357914 538718
rect 357294 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 357914 538634
rect 357294 502954 357914 538398
rect 357294 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 357914 502954
rect 357294 502634 357914 502718
rect 357294 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 357914 502634
rect 357294 466954 357914 502398
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 430954 357914 466398
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 357294 430634 357914 430718
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 214954 357914 250398
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 241954 384914 277398
rect 384294 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 384914 241954
rect 384294 241634 384914 241718
rect 384294 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 384914 241634
rect 384294 205954 384914 241398
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 210454 389414 245898
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 214954 393914 250398
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< obsm4 >>
rect 68800 174494 96960 174600
rect 97020 174494 98320 174600
rect 98380 174494 99408 174600
rect 99468 174494 100768 174600
rect 100828 174494 101992 174600
rect 102052 174494 103352 174600
rect 103412 174494 104576 174600
rect 104636 174494 105664 174600
rect 105724 174494 107024 174600
rect 107084 174494 108112 174600
rect 108172 174494 109472 174600
rect 109532 174494 110696 174600
rect 110756 174494 112056 174600
rect 112116 174494 113144 174600
rect 113204 174494 114368 174600
rect 114428 174494 115728 174600
rect 115788 174494 116952 174600
rect 117012 174494 118312 174600
rect 118372 174494 119400 174600
rect 119460 174494 120760 174600
rect 120820 174494 121848 174600
rect 121908 174494 123072 174600
rect 123132 174494 124432 174600
rect 124492 174494 125656 174600
rect 125716 174494 127016 174600
rect 127076 174494 128104 174600
rect 128164 174494 129464 174600
rect 129524 174494 130688 174600
rect 130748 174494 132048 174600
rect 132108 174494 133136 174600
rect 133196 174494 134360 174600
rect 134420 174494 135720 174600
rect 135780 174494 148232 174600
rect 148292 174494 158840 174600
rect 158900 174494 164756 174600
rect 68800 151986 164756 174494
rect 68800 151366 69072 151986
rect 69420 151366 164136 151986
rect 164484 151366 164756 151986
rect 68800 147486 164756 151366
rect 68800 146866 69752 147486
rect 70100 146866 163456 147486
rect 163804 146866 164756 147486
rect 68800 115986 164756 146866
rect 68800 115366 69072 115986
rect 69420 115366 164136 115986
rect 164484 115366 164756 115986
rect 68800 111486 164756 115366
rect 68800 110866 69752 111486
rect 70100 110866 163456 111486
rect 163804 110866 164756 111486
rect 68800 95200 164756 110866
rect 68800 95100 74656 95200
rect 74716 95100 84312 95200
rect 84372 95100 85536 95200
rect 85596 95100 86624 95200
rect 86684 95100 87984 95200
rect 88044 95100 88936 95200
rect 88996 95100 90160 95200
rect 90220 95100 91384 95200
rect 91444 95100 92472 95200
rect 92532 95100 93832 95200
rect 93892 95100 94920 95200
rect 94980 95100 96008 95200
rect 96068 95100 96688 95200
rect 96748 95100 97096 95200
rect 97156 95100 98048 95200
rect 98108 95100 98456 95200
rect 98516 95100 99136 95200
rect 99196 95100 99544 95200
rect 99604 95100 100632 95200
rect 100692 95100 100768 95200
rect 100828 95100 101856 95200
rect 101916 95100 101992 95200
rect 102052 95100 102944 95200
rect 103004 95100 103216 95200
rect 103276 95100 104304 95200
rect 104364 95100 104440 95200
rect 104500 95100 105392 95200
rect 105452 95100 105664 95200
rect 105724 95100 106480 95200
rect 106540 95100 106616 95200
rect 106676 95100 107704 95200
rect 107764 95100 108112 95200
rect 108172 95100 109064 95200
rect 109124 95100 109472 95200
rect 109532 95100 110152 95200
rect 110212 95100 110696 95200
rect 110756 95100 111240 95200
rect 111300 95100 111920 95200
rect 111980 95100 112328 95200
rect 112388 95100 113144 95200
rect 113204 95100 113688 95200
rect 113748 95100 114368 95200
rect 114428 95100 114776 95200
rect 114836 95100 115456 95200
rect 115516 95100 115864 95200
rect 115924 95100 116680 95200
rect 116740 95100 117088 95200
rect 117148 95100 117904 95200
rect 117964 95100 118176 95200
rect 118236 95100 119400 95200
rect 119460 95100 119536 95200
rect 119596 95100 120216 95200
rect 120276 95100 120624 95200
rect 120684 95100 121712 95200
rect 121772 95100 121984 95200
rect 122044 95100 122800 95200
rect 122860 95100 123208 95200
rect 123268 95100 124024 95200
rect 124084 95100 124432 95200
rect 124492 95100 125384 95200
rect 125444 95100 125656 95200
rect 125716 95100 126472 95200
rect 126532 95100 126608 95200
rect 126668 95100 128104 95200
rect 128164 95100 129328 95200
rect 129388 95100 130688 95200
rect 130748 95100 131912 95200
rect 131972 95100 133136 95200
rect 133196 95100 134360 95200
rect 134420 95100 135584 95200
rect 135644 95100 151496 95200
rect 151556 95100 151632 95200
rect 151692 95100 151768 95200
rect 151828 95100 151904 95200
rect 151964 95100 164756 95200
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 89610 259718 89846 259954
rect 89610 259398 89846 259634
rect 74250 255218 74486 255454
rect 74250 254898 74486 255134
rect 104970 255218 105206 255454
rect 104970 254898 105206 255134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 118826 228218 119062 228454
rect 119146 228218 119382 228454
rect 118826 227898 119062 228134
rect 119146 227898 119382 228134
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 123326 232718 123562 232954
rect 123646 232718 123882 232954
rect 123326 232398 123562 232634
rect 123646 232398 123882 232634
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 132326 241718 132562 241954
rect 132646 241718 132882 241954
rect 132326 241398 132562 241634
rect 132646 241398 132882 241634
rect 132326 205718 132562 205954
rect 132646 205718 132882 205954
rect 132326 205398 132562 205634
rect 132646 205398 132882 205634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 136826 246218 137062 246454
rect 137146 246218 137382 246454
rect 136826 245898 137062 246134
rect 137146 245898 137382 246134
rect 136826 210218 137062 210454
rect 137146 210218 137382 210454
rect 136826 209898 137062 210134
rect 137146 209898 137382 210134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 141326 214718 141562 214954
rect 141646 214718 141882 214954
rect 141326 214398 141562 214634
rect 141646 214398 141882 214634
rect 141326 178718 141562 178954
rect 141646 178718 141882 178954
rect 141326 178398 141562 178634
rect 141646 178398 141882 178634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 150326 223718 150562 223954
rect 150646 223718 150882 223954
rect 150326 223398 150562 223634
rect 150646 223398 150882 223634
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 154826 228218 155062 228454
rect 155146 228218 155382 228454
rect 154826 227898 155062 228134
rect 155146 227898 155382 228134
rect 150326 187718 150562 187954
rect 150646 187718 150882 187954
rect 150326 187398 150562 187634
rect 150646 187398 150882 187634
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 159326 232718 159562 232954
rect 159646 232718 159882 232954
rect 159326 232398 159562 232634
rect 159646 232398 159882 232634
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 168326 241718 168562 241954
rect 168646 241718 168882 241954
rect 168326 241398 168562 241634
rect 168646 241398 168882 241634
rect 168326 205718 168562 205954
rect 168646 205718 168882 205954
rect 168326 205398 168562 205634
rect 168646 205398 168882 205634
rect 168326 169718 168562 169954
rect 168646 169718 168882 169954
rect 168326 169398 168562 169634
rect 168646 169398 168882 169634
rect 69128 151718 69364 151954
rect 69128 151398 69364 151634
rect 164192 151718 164428 151954
rect 164192 151398 164428 151634
rect 69808 147218 70044 147454
rect 69808 146898 70044 147134
rect 163512 147218 163748 147454
rect 163512 146898 163748 147134
rect 69128 115718 69364 115954
rect 69128 115398 69364 115634
rect 164192 115718 164428 115954
rect 164192 115398 164428 115634
rect 69808 111218 70044 111454
rect 69808 110898 70044 111134
rect 163512 111218 163748 111454
rect 163512 110898 163748 111134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 84218 119062 84454
rect 119146 84218 119382 84454
rect 118826 83898 119062 84134
rect 119146 83898 119382 84134
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 88718 123562 88954
rect 123646 88718 123882 88954
rect 123326 88398 123562 88634
rect 123646 88398 123882 88634
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 79718 150562 79954
rect 150646 79718 150882 79954
rect 150326 79398 150562 79634
rect 150646 79398 150882 79634
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 154826 84218 155062 84454
rect 155146 84218 155382 84454
rect 154826 83898 155062 84134
rect 155146 83898 155382 84134
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 159326 88718 159562 88954
rect 159646 88718 159882 88954
rect 159326 88398 159562 88634
rect 159646 88398 159882 88634
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 168326 133718 168562 133954
rect 168646 133718 168882 133954
rect 168326 133398 168562 133634
rect 168646 133398 168882 133634
rect 168326 97718 168562 97954
rect 168646 97718 168882 97954
rect 168326 97398 168562 97634
rect 168646 97398 168882 97634
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 172826 246218 173062 246454
rect 173146 246218 173382 246454
rect 172826 245898 173062 246134
rect 173146 245898 173382 246134
rect 172826 210218 173062 210454
rect 173146 210218 173382 210454
rect 172826 209898 173062 210134
rect 173146 209898 173382 210134
rect 172826 174218 173062 174454
rect 173146 174218 173382 174454
rect 172826 173898 173062 174134
rect 173146 173898 173382 174134
rect 172826 138218 173062 138454
rect 173146 138218 173382 138454
rect 172826 137898 173062 138134
rect 173146 137898 173382 138134
rect 172826 102218 173062 102454
rect 173146 102218 173382 102454
rect 172826 101898 173062 102134
rect 173146 101898 173382 102134
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 222326 547718 222562 547954
rect 222646 547718 222882 547954
rect 222326 547398 222562 547634
rect 222646 547398 222882 547634
rect 222326 511718 222562 511954
rect 222646 511718 222882 511954
rect 222326 511398 222562 511634
rect 222646 511398 222882 511634
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 226826 552218 227062 552454
rect 227146 552218 227382 552454
rect 226826 551898 227062 552134
rect 227146 551898 227382 552134
rect 226826 516218 227062 516454
rect 227146 516218 227382 516454
rect 226826 515898 227062 516134
rect 227146 515898 227382 516134
rect 226826 480218 227062 480454
rect 227146 480218 227382 480454
rect 226826 479898 227062 480134
rect 227146 479898 227382 480134
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 231326 556718 231562 556954
rect 231646 556718 231882 556954
rect 231326 556398 231562 556634
rect 231646 556398 231882 556634
rect 231326 520718 231562 520954
rect 231646 520718 231882 520954
rect 231326 520398 231562 520634
rect 231646 520398 231882 520634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 231326 412718 231562 412954
rect 231646 412718 231882 412954
rect 231326 412398 231562 412634
rect 231646 412398 231882 412634
rect 231326 376718 231562 376954
rect 231646 376718 231882 376954
rect 231326 376398 231562 376634
rect 231646 376398 231882 376634
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 240326 529718 240562 529954
rect 240646 529718 240882 529954
rect 240326 529398 240562 529634
rect 240646 529398 240882 529634
rect 240326 493718 240562 493954
rect 240646 493718 240882 493954
rect 240326 493398 240562 493634
rect 240646 493398 240882 493634
rect 240326 457718 240562 457954
rect 240646 457718 240882 457954
rect 240326 457398 240562 457634
rect 240646 457398 240882 457634
rect 240326 421718 240562 421954
rect 240646 421718 240882 421954
rect 240326 421398 240562 421634
rect 240646 421398 240882 421634
rect 240326 385718 240562 385954
rect 240646 385718 240882 385954
rect 240326 385398 240562 385634
rect 240646 385398 240882 385634
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 244826 534218 245062 534454
rect 245146 534218 245382 534454
rect 244826 533898 245062 534134
rect 245146 533898 245382 534134
rect 244826 498218 245062 498454
rect 245146 498218 245382 498454
rect 244826 497898 245062 498134
rect 245146 497898 245382 498134
rect 244826 462218 245062 462454
rect 245146 462218 245382 462454
rect 244826 461898 245062 462134
rect 245146 461898 245382 462134
rect 244826 426218 245062 426454
rect 245146 426218 245382 426454
rect 244826 425898 245062 426134
rect 245146 425898 245382 426134
rect 244826 390218 245062 390454
rect 245146 390218 245382 390454
rect 244826 389898 245062 390134
rect 245146 389898 245382 390134
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 249326 538718 249562 538954
rect 249646 538718 249882 538954
rect 249326 538398 249562 538634
rect 249646 538398 249882 538634
rect 249326 502718 249562 502954
rect 249646 502718 249882 502954
rect 249326 502398 249562 502634
rect 249646 502398 249882 502634
rect 249326 466718 249562 466954
rect 249646 466718 249882 466954
rect 249326 466398 249562 466634
rect 249646 466398 249882 466634
rect 249326 430718 249562 430954
rect 249646 430718 249882 430954
rect 249326 430398 249562 430634
rect 249646 430398 249882 430634
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 249326 358718 249562 358954
rect 249646 358718 249882 358954
rect 249326 358398 249562 358634
rect 249646 358398 249882 358634
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 276326 529718 276562 529954
rect 276646 529718 276882 529954
rect 276326 529398 276562 529634
rect 276646 529398 276882 529634
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 280826 534218 281062 534454
rect 281146 534218 281382 534454
rect 280826 533898 281062 534134
rect 281146 533898 281382 534134
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 199610 331718 199846 331954
rect 199610 331398 199846 331634
rect 230330 331718 230566 331954
rect 230330 331398 230566 331634
rect 261050 331718 261286 331954
rect 261050 331398 261286 331634
rect 184250 327218 184486 327454
rect 184250 326898 184486 327134
rect 214970 327218 215206 327454
rect 214970 326898 215206 327134
rect 245690 327218 245926 327454
rect 245690 326898 245926 327134
rect 276410 327218 276646 327454
rect 276410 326898 276646 327134
rect 199610 295718 199846 295954
rect 199610 295398 199846 295634
rect 230330 295718 230566 295954
rect 230330 295398 230566 295634
rect 261050 295718 261286 295954
rect 261050 295398 261286 295634
rect 184250 291218 184486 291454
rect 184250 290898 184486 291134
rect 214970 291218 215206 291454
rect 214970 290898 215206 291134
rect 245690 291218 245926 291454
rect 245690 290898 245926 291134
rect 276410 291218 276646 291454
rect 276410 290898 276646 291134
rect 199610 259718 199846 259954
rect 199610 259398 199846 259634
rect 230330 259718 230566 259954
rect 230330 259398 230566 259634
rect 261050 259718 261286 259954
rect 261050 259398 261286 259634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 184250 255218 184486 255454
rect 184250 254898 184486 255134
rect 214970 255218 215206 255454
rect 214970 254898 215206 255134
rect 245690 255218 245926 255454
rect 245690 254898 245926 255134
rect 276410 255218 276646 255454
rect 276410 254898 276646 255134
rect 177326 214718 177562 214954
rect 177646 214718 177882 214954
rect 177326 214398 177562 214634
rect 177646 214398 177882 214634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 177326 106718 177562 106954
rect 177646 106718 177882 106954
rect 177326 106398 177562 106634
rect 177646 106398 177882 106634
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 186326 115718 186562 115954
rect 186646 115718 186882 115954
rect 186326 115398 186562 115634
rect 186646 115398 186882 115634
rect 186326 79718 186562 79954
rect 186646 79718 186882 79954
rect 186326 79398 186562 79634
rect 186646 79398 186882 79634
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 228218 191062 228454
rect 191146 228218 191382 228454
rect 190826 227898 191062 228134
rect 191146 227898 191382 228134
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 190826 120218 191062 120454
rect 191146 120218 191382 120454
rect 190826 119898 191062 120134
rect 191146 119898 191382 120134
rect 190826 84218 191062 84454
rect 191146 84218 191382 84454
rect 190826 83898 191062 84134
rect 191146 83898 191382 84134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 232718 195562 232954
rect 195646 232718 195882 232954
rect 195326 232398 195562 232634
rect 195646 232398 195882 232634
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 226826 228218 227062 228454
rect 227146 228218 227382 228454
rect 226826 227898 227062 228134
rect 227146 227898 227382 228134
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 231326 232718 231562 232954
rect 231646 232718 231882 232954
rect 231326 232398 231562 232634
rect 231646 232398 231882 232634
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 227916 151718 228152 151954
rect 227916 151398 228152 151634
rect 237847 151718 238083 151954
rect 237847 151398 238083 151634
rect 222952 147218 223188 147454
rect 222952 146898 223188 147134
rect 232882 147218 233118 147454
rect 232882 146898 233118 147134
rect 242813 147218 243049 147454
rect 242813 146898 243049 147134
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 227916 115718 228152 115954
rect 227916 115398 228152 115634
rect 237847 115718 238083 115954
rect 237847 115398 238083 115634
rect 222952 111218 223188 111454
rect 222952 110898 223188 111134
rect 232882 111218 233118 111454
rect 232882 110898 233118 111134
rect 242813 111218 243049 111454
rect 242813 110898 243049 111134
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 262826 228218 263062 228454
rect 263146 228218 263382 228454
rect 262826 227898 263062 228134
rect 263146 227898 263382 228134
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 267326 232718 267562 232954
rect 267646 232718 267882 232954
rect 267326 232398 267562 232634
rect 267646 232398 267882 232634
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 298826 516218 299062 516454
rect 299146 516218 299382 516454
rect 298826 515898 299062 516134
rect 299146 515898 299382 516134
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 303326 556718 303562 556954
rect 303646 556718 303882 556954
rect 303326 556398 303562 556634
rect 303646 556398 303882 556634
rect 303326 520718 303562 520954
rect 303646 520718 303882 520954
rect 303326 520398 303562 520634
rect 303646 520398 303882 520634
rect 303326 484718 303562 484954
rect 303646 484718 303882 484954
rect 298826 480218 299062 480454
rect 299146 480218 299382 480454
rect 298826 479898 299062 480134
rect 299146 479898 299382 480134
rect 298826 444218 299062 444454
rect 299146 444218 299382 444454
rect 298826 443898 299062 444134
rect 299146 443898 299382 444134
rect 298826 408218 299062 408454
rect 299146 408218 299382 408454
rect 298826 407898 299062 408134
rect 299146 407898 299382 408134
rect 298826 372218 299062 372454
rect 299146 372218 299382 372454
rect 298826 371898 299062 372134
rect 299146 371898 299382 372134
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 303326 484398 303562 484634
rect 303646 484398 303882 484634
rect 303326 448718 303562 448954
rect 303646 448718 303882 448954
rect 303326 448398 303562 448634
rect 303646 448398 303882 448634
rect 303326 412718 303562 412954
rect 303646 412718 303882 412954
rect 303326 412398 303562 412634
rect 303646 412398 303882 412634
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 298826 228218 299062 228454
rect 299146 228218 299382 228454
rect 298826 227898 299062 228134
rect 299146 227898 299382 228134
rect 298826 192218 299062 192454
rect 299146 192218 299382 192454
rect 298826 191898 299062 192134
rect 299146 191898 299382 192134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 303326 232718 303562 232954
rect 303646 232718 303882 232954
rect 303326 232398 303562 232634
rect 303646 232398 303882 232634
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 312326 529718 312562 529954
rect 312646 529718 312882 529954
rect 312326 529398 312562 529634
rect 312646 529398 312882 529634
rect 312326 493718 312562 493954
rect 312646 493718 312882 493954
rect 312326 493398 312562 493634
rect 312646 493398 312882 493634
rect 312326 457718 312562 457954
rect 312646 457718 312882 457954
rect 312326 457398 312562 457634
rect 312646 457398 312882 457634
rect 312326 421718 312562 421954
rect 312646 421718 312882 421954
rect 312326 421398 312562 421634
rect 312646 421398 312882 421634
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 312326 313718 312562 313954
rect 312646 313718 312882 313954
rect 312326 313398 312562 313634
rect 312646 313398 312882 313634
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 312326 241718 312562 241954
rect 312646 241718 312882 241954
rect 312326 241398 312562 241634
rect 312646 241398 312882 241634
rect 312326 205718 312562 205954
rect 312646 205718 312882 205954
rect 312326 205398 312562 205634
rect 312646 205398 312882 205634
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 316826 534218 317062 534454
rect 317146 534218 317382 534454
rect 316826 533898 317062 534134
rect 317146 533898 317382 534134
rect 316826 498218 317062 498454
rect 317146 498218 317382 498454
rect 316826 497898 317062 498134
rect 317146 497898 317382 498134
rect 316826 462218 317062 462454
rect 317146 462218 317382 462454
rect 316826 461898 317062 462134
rect 317146 461898 317382 462134
rect 316826 426218 317062 426454
rect 317146 426218 317382 426454
rect 316826 425898 317062 426134
rect 317146 425898 317382 426134
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 316826 318218 317062 318454
rect 317146 318218 317382 318454
rect 316826 317898 317062 318134
rect 317146 317898 317382 318134
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 316826 246218 317062 246454
rect 317146 246218 317382 246454
rect 316826 245898 317062 246134
rect 317146 245898 317382 246134
rect 316826 210218 317062 210454
rect 317146 210218 317382 210454
rect 316826 209898 317062 210134
rect 317146 209898 317382 210134
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 321326 538718 321562 538954
rect 321646 538718 321882 538954
rect 321326 538398 321562 538634
rect 321646 538398 321882 538634
rect 321326 502718 321562 502954
rect 321646 502718 321882 502954
rect 321326 502398 321562 502634
rect 321646 502398 321882 502634
rect 321326 466718 321562 466954
rect 321646 466718 321882 466954
rect 321326 466398 321562 466634
rect 321646 466398 321882 466634
rect 321326 430718 321562 430954
rect 321646 430718 321882 430954
rect 321326 430398 321562 430634
rect 321646 430398 321882 430634
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 321326 322718 321562 322954
rect 321646 322718 321882 322954
rect 321326 322398 321562 322634
rect 321646 322398 321882 322634
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 321326 214718 321562 214954
rect 321646 214718 321882 214954
rect 321326 214398 321562 214634
rect 321646 214398 321882 214634
rect 321326 178718 321562 178954
rect 321646 178718 321882 178954
rect 321326 178398 321562 178634
rect 321646 178398 321882 178634
rect 314250 151718 314486 151954
rect 314250 151398 314486 151634
rect 317514 151718 317750 151954
rect 317514 151398 317750 151634
rect 312618 147218 312854 147454
rect 312618 146898 312854 147134
rect 315882 147218 316118 147454
rect 315882 146898 316118 147134
rect 319146 147218 319382 147454
rect 319146 146898 319382 147134
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 330326 511718 330562 511954
rect 330646 511718 330882 511954
rect 330326 511398 330562 511634
rect 330646 511398 330882 511634
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 330326 439718 330562 439954
rect 330646 439718 330882 439954
rect 330326 439398 330562 439634
rect 330646 439398 330882 439634
rect 330326 403718 330562 403954
rect 330646 403718 330882 403954
rect 330326 403398 330562 403634
rect 330646 403398 330882 403634
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 334826 516218 335062 516454
rect 335146 516218 335382 516454
rect 334826 515898 335062 516134
rect 335146 515898 335382 516134
rect 334826 480218 335062 480454
rect 335146 480218 335382 480454
rect 334826 479898 335062 480134
rect 335146 479898 335382 480134
rect 334826 444218 335062 444454
rect 335146 444218 335382 444454
rect 334826 443898 335062 444134
rect 335146 443898 335382 444134
rect 334826 408218 335062 408454
rect 335146 408218 335382 408454
rect 334826 407898 335062 408134
rect 335146 407898 335382 408134
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 314250 115718 314486 115954
rect 314250 115398 314486 115634
rect 317514 115718 317750 115954
rect 317514 115398 317750 115634
rect 312618 111218 312854 111454
rect 312618 110898 312854 111134
rect 315882 111218 316118 111454
rect 315882 110898 316118 111134
rect 319146 111218 319382 111454
rect 319146 110898 319382 111134
rect 330326 223718 330562 223954
rect 330646 223718 330882 223954
rect 330326 223398 330562 223634
rect 330646 223398 330882 223634
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 330326 187718 330562 187954
rect 330646 187718 330882 187954
rect 330326 187398 330562 187634
rect 330646 187398 330882 187634
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 334826 228218 335062 228454
rect 335146 228218 335382 228454
rect 334826 227898 335062 228134
rect 335146 227898 335382 228134
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 339326 556718 339562 556954
rect 339646 556718 339882 556954
rect 339326 556398 339562 556634
rect 339646 556398 339882 556634
rect 339326 520718 339562 520954
rect 339646 520718 339882 520954
rect 339326 520398 339562 520634
rect 339646 520398 339882 520634
rect 339326 484718 339562 484954
rect 339646 484718 339882 484954
rect 339326 484398 339562 484634
rect 339646 484398 339882 484634
rect 339326 448718 339562 448954
rect 339646 448718 339882 448954
rect 339326 448398 339562 448634
rect 339646 448398 339882 448634
rect 339326 412718 339562 412954
rect 339646 412718 339882 412954
rect 339326 412398 339562 412634
rect 339646 412398 339882 412634
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 339326 232718 339562 232954
rect 339646 232718 339882 232954
rect 339326 232398 339562 232634
rect 339646 232398 339882 232634
rect 334826 192218 335062 192454
rect 335146 192218 335382 192454
rect 334826 191898 335062 192134
rect 335146 191898 335382 192134
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 348326 529718 348562 529954
rect 348646 529718 348882 529954
rect 348326 529398 348562 529634
rect 348646 529398 348882 529634
rect 348326 493718 348562 493954
rect 348646 493718 348882 493954
rect 348326 493398 348562 493634
rect 348646 493398 348882 493634
rect 348326 457718 348562 457954
rect 348646 457718 348882 457954
rect 348326 457398 348562 457634
rect 348646 457398 348882 457634
rect 348326 421718 348562 421954
rect 348646 421718 348882 421954
rect 348326 421398 348562 421634
rect 348646 421398 348882 421634
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 348326 313718 348562 313954
rect 348646 313718 348882 313954
rect 348326 313398 348562 313634
rect 348646 313398 348882 313634
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 348326 241718 348562 241954
rect 348646 241718 348882 241954
rect 348326 241398 348562 241634
rect 348646 241398 348882 241634
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 348326 205718 348562 205954
rect 348646 205718 348882 205954
rect 348326 205398 348562 205634
rect 348646 205398 348882 205634
rect 348326 169718 348562 169954
rect 348646 169718 348882 169954
rect 348326 169398 348562 169634
rect 348646 169398 348882 169634
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 352826 426218 353062 426454
rect 353146 426218 353382 426454
rect 352826 425898 353062 426134
rect 353146 425898 353382 426134
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 357326 538718 357562 538954
rect 357646 538718 357882 538954
rect 357326 538398 357562 538634
rect 357646 538398 357882 538634
rect 357326 502718 357562 502954
rect 357646 502718 357882 502954
rect 357326 502398 357562 502634
rect 357646 502398 357882 502634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 384326 241718 384562 241954
rect 384646 241718 384882 241954
rect 384326 241398 384562 241634
rect 384646 241398 384882 241634
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 199610 331954
rect 199846 331718 230330 331954
rect 230566 331718 261050 331954
rect 261286 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 199610 331634
rect 199846 331398 230330 331634
rect 230566 331398 261050 331634
rect 261286 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 184250 327454
rect 184486 327218 214970 327454
rect 215206 327218 245690 327454
rect 245926 327218 276410 327454
rect 276646 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 184250 327134
rect 184486 326898 214970 327134
rect 215206 326898 245690 327134
rect 245926 326898 276410 327134
rect 276646 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 199610 295954
rect 199846 295718 230330 295954
rect 230566 295718 261050 295954
rect 261286 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 199610 295634
rect 199846 295398 230330 295634
rect 230566 295398 261050 295634
rect 261286 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 184250 291454
rect 184486 291218 214970 291454
rect 215206 291218 245690 291454
rect 245926 291218 276410 291454
rect 276646 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 184250 291134
rect 184486 290898 214970 291134
rect 215206 290898 245690 291134
rect 245926 290898 276410 291134
rect 276646 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 89610 259954
rect 89846 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 199610 259954
rect 199846 259718 230330 259954
rect 230566 259718 261050 259954
rect 261286 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 89610 259634
rect 89846 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 199610 259634
rect 199846 259398 230330 259634
rect 230566 259398 261050 259634
rect 261286 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 74250 255454
rect 74486 255218 104970 255454
rect 105206 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 184250 255454
rect 184486 255218 214970 255454
rect 215206 255218 245690 255454
rect 245926 255218 276410 255454
rect 276646 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 74250 255134
rect 74486 254898 104970 255134
rect 105206 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 184250 255134
rect 184486 254898 214970 255134
rect 215206 254898 245690 255134
rect 245926 254898 276410 255134
rect 276646 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 69128 151954
rect 69364 151718 164192 151954
rect 164428 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 227916 151954
rect 228152 151718 237847 151954
rect 238083 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 314250 151954
rect 314486 151718 317514 151954
rect 317750 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 69128 151634
rect 69364 151398 164192 151634
rect 164428 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 227916 151634
rect 228152 151398 237847 151634
rect 238083 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 314250 151634
rect 314486 151398 317514 151634
rect 317750 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 69808 147454
rect 70044 147218 163512 147454
rect 163748 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 222952 147454
rect 223188 147218 232882 147454
rect 233118 147218 242813 147454
rect 243049 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 312618 147454
rect 312854 147218 315882 147454
rect 316118 147218 319146 147454
rect 319382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 69808 147134
rect 70044 146898 163512 147134
rect 163748 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 222952 147134
rect 223188 146898 232882 147134
rect 233118 146898 242813 147134
rect 243049 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 312618 147134
rect 312854 146898 315882 147134
rect 316118 146898 319146 147134
rect 319382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 69128 115954
rect 69364 115718 164192 115954
rect 164428 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 227916 115954
rect 228152 115718 237847 115954
rect 238083 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 314250 115954
rect 314486 115718 317514 115954
rect 317750 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 69128 115634
rect 69364 115398 164192 115634
rect 164428 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 227916 115634
rect 228152 115398 237847 115634
rect 238083 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 314250 115634
rect 314486 115398 317514 115634
rect 317750 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 69808 111454
rect 70044 111218 163512 111454
rect 163748 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 222952 111454
rect 223188 111218 232882 111454
rect 233118 111218 242813 111454
rect 243049 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 312618 111454
rect 312854 111218 315882 111454
rect 316118 111218 319146 111454
rect 319382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 69808 111134
rect 70044 110898 163512 111134
rect 163748 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 222952 111134
rect 223188 110898 232882 111134
rect 233118 110898 242813 111134
rect 243049 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 312618 111134
rect 312854 110898 315882 111134
rect 316118 110898 319146 111134
rect 319382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use sky130_sram_1kbyte_1rw1r_32x256_8  openram_1kB
timestamp 0
transform 1 0 68800 0 1 95100
box 0 0 95956 79500
use wb_bridge_2way  wb_bridge_2way
timestamp 0
transform 1 0 310000 0 1 96000
box 0 144 12000 80000
use wb_openram_wrapper  wb_openram_wrapper
timestamp 0
transform 1 0 217000 0 1 96000
box 0 144 32000 79688
use wrapped_function_generator  wrapped_function_generator_0
timestamp 0
transform 1 0 70000 0 1 240000
box 0 0 50000 52000
use wrapped_ibnalhaytham  wrapped_ibnalhaytham_1
timestamp 0
transform 1 0 180000 0 1 240000
box 0 0 113010 115154
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 93100 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 176600 74414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 294000 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 93100 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 176600 110414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 294000 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 93100 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 176600 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 357154 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 94000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 178000 218414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 357154 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 357154 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 357154 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 93100 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 176600 83414 238000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 294000 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 93100 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 176600 119414 238000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 294000 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 93100 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 176600 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 238000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 357154 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 94000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 178000 227414 238000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 357154 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 238000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 357154 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 93100 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 176600 92414 238000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 294000 92414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 93100 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 176600 128414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 93100 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 176600 164414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 238000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 357154 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 94000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 178000 236414 238000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 357154 236414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 238000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 357154 272414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 94000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 178000 308414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 -7654 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 -7654 101414 93100 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 294000 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 93100 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 176600 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 -7654 209414 238000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 357154 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 -7654 245414 94000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 357154 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 -7654 281414 238000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 357154 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 -7654 317414 94000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 178000 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 -7654 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 -7654 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 93100 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 294000 96914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 93100 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 176600 132914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 238000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 357154 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 94000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 357154 240914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 238000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 357154 276914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 94000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 178000 312914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 93100 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 176600 69914 238000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 294000 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 93100 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 176600 105914 238000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 294000 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 93100 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 176600 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 238000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 357154 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 94000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 178000 249914 238000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 357154 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 238000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 357154 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 94000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 178000 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 93100 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 176600 78914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 294000 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 93100 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 176600 114914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 294000 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 93100 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 176600 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 357154 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 94000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 178000 222914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 357154 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 357154 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 357154 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 93100 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 176600 87914 238000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 294000 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 93100 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 176600 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 93100 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 176600 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 238000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 357154 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 94000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 178000 231914 238000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 357154 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 238000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 357154 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
