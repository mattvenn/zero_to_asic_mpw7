magic
tech sky130B
magscale 1 2
timestamp 1657720573
<< obsli1 >>
rect 0 0 584000 704000
<< metal1 >>
rect 201494 703060 201500 703112
rect 201552 703100 201558 703112
rect 202782 703100 202788 703112
rect 201552 703072 202788 703100
rect 201552 703060 201558 703072
rect 202782 703060 202788 703072
rect 202840 703060 202846 703112
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 84286 702992 84292 703044
rect 84344 703032 84350 703044
rect 348786 703032 348792 703044
rect 84344 703004 348792 703032
rect 84344 702992 84350 703004
rect 348786 702992 348792 703004
rect 348844 702992 348850 703044
rect 107654 702924 107660 702976
rect 107712 702964 107718 702976
rect 413646 702964 413652 702976
rect 107712 702936 413652 702964
rect 107712 702924 107718 702936
rect 413646 702924 413652 702936
rect 413704 702924 413710 702976
rect 128998 702856 129004 702908
rect 129056 702896 129062 702908
rect 462314 702896 462320 702908
rect 129056 702868 462320 702896
rect 129056 702856 129062 702868
rect 462314 702856 462320 702868
rect 462372 702856 462378 702908
rect 49602 702788 49608 702840
rect 49660 702828 49666 702840
rect 397454 702828 397460 702840
rect 49660 702800 397460 702828
rect 49660 702788 49666 702800
rect 397454 702788 397460 702800
rect 397512 702788 397518 702840
rect 63402 702720 63408 702772
rect 63460 702760 63466 702772
rect 429838 702760 429844 702772
rect 63460 702732 429844 702760
rect 63460 702720 63466 702732
rect 429838 702720 429844 702732
rect 429896 702720 429902 702772
rect 106274 702652 106280 702704
rect 106332 702692 106338 702704
rect 478506 702692 478512 702704
rect 106332 702664 478512 702692
rect 106332 702652 106338 702664
rect 478506 702652 478512 702664
rect 478564 702652 478570 702704
rect 124858 702584 124864 702636
rect 124916 702624 124922 702636
rect 527174 702624 527180 702636
rect 124916 702596 527180 702624
rect 124916 702584 124922 702596
rect 527174 702584 527180 702596
rect 527232 702584 527238 702636
rect 134518 702516 134524 702568
rect 134576 702556 134582 702568
rect 559650 702556 559656 702568
rect 134576 702528 559656 702556
rect 134576 702516 134582 702528
rect 559650 702516 559656 702528
rect 559708 702516 559714 702568
rect 80698 702448 80704 702500
rect 80756 702488 80762 702500
rect 580902 702488 580908 702500
rect 80756 702460 580908 702488
rect 80756 702448 80762 702460
rect 580902 702448 580908 702460
rect 580960 702448 580966 702500
rect 55122 700408 55128 700460
rect 55180 700448 55186 700460
rect 105446 700448 105452 700460
rect 55180 700420 105452 700448
rect 55180 700408 55186 700420
rect 105446 700408 105452 700420
rect 105504 700408 105510 700460
rect 149698 700408 149704 700460
rect 149756 700448 149762 700460
rect 235166 700448 235172 700460
rect 149756 700420 235172 700448
rect 149756 700408 149762 700420
rect 235166 700408 235172 700420
rect 235224 700408 235230 700460
rect 57882 700340 57888 700392
rect 57940 700380 57946 700392
rect 170306 700380 170312 700392
rect 57940 700352 170312 700380
rect 57940 700340 57946 700352
rect 170306 700340 170312 700352
rect 170364 700340 170370 700392
rect 269758 700340 269764 700392
rect 269816 700380 269822 700392
rect 332502 700380 332508 700392
rect 269816 700352 332508 700380
rect 269816 700340 269822 700352
rect 332502 700340 332508 700352
rect 332560 700340 332566 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 8938 700312 8944 700324
rect 8168 700284 8944 700312
rect 8168 700272 8174 700284
rect 8938 700272 8944 700284
rect 8996 700272 9002 700324
rect 24302 700272 24308 700324
rect 24360 700312 24366 700324
rect 82078 700312 82084 700324
rect 24360 700284 82084 700312
rect 24360 700272 24366 700284
rect 82078 700272 82084 700284
rect 82136 700272 82142 700324
rect 135898 700272 135904 700324
rect 135956 700312 135962 700324
rect 364978 700312 364984 700324
rect 135956 700284 364984 700312
rect 135956 700272 135962 700284
rect 364978 700272 364984 700284
rect 365036 700272 365042 700324
rect 214558 699660 214564 699712
rect 214616 699700 214622 699712
rect 218974 699700 218980 699712
rect 214616 699672 218980 699700
rect 214616 699660 214622 699672
rect 218974 699660 218980 699672
rect 219032 699660 219038 699712
rect 264238 699660 264244 699712
rect 264296 699700 264302 699712
rect 267642 699700 267648 699712
rect 264296 699672 267648 699700
rect 264296 699660 264302 699672
rect 267642 699660 267648 699672
rect 267700 699660 267706 699712
rect 59262 697552 59268 697604
rect 59320 697592 59326 697604
rect 137830 697592 137836 697604
rect 59320 697564 137836 697592
rect 59320 697552 59326 697564
rect 137830 697552 137836 697564
rect 137888 697552 137894 697604
rect 53742 696192 53748 696244
rect 53800 696232 53806 696244
rect 300118 696232 300124 696244
rect 53800 696204 300124 696232
rect 53800 696192 53806 696204
rect 300118 696192 300124 696204
rect 300176 696192 300182 696244
rect 144178 683136 144184 683188
rect 144236 683176 144242 683188
rect 580166 683176 580172 683188
rect 144236 683148 580172 683176
rect 144236 683136 144242 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 26878 670732 26884 670744
rect 3568 670704 26884 670732
rect 3568 670692 3574 670704
rect 26878 670692 26884 670704
rect 26936 670692 26942 670744
rect 148318 670692 148324 670744
rect 148376 670732 148382 670744
rect 580166 670732 580172 670744
rect 148376 670704 580172 670732
rect 148376 670692 148382 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3510 656888 3516 656940
rect 3568 656928 3574 656940
rect 39298 656928 39304 656940
rect 3568 656900 39304 656928
rect 3568 656888 3574 656900
rect 39298 656888 39304 656900
rect 39356 656888 39362 656940
rect 3510 632068 3516 632120
rect 3568 632108 3574 632120
rect 21358 632108 21364 632120
rect 3568 632080 21364 632108
rect 3568 632068 3574 632080
rect 21358 632068 21364 632080
rect 21416 632068 21422 632120
rect 126238 630640 126244 630692
rect 126296 630680 126302 630692
rect 580166 630680 580172 630692
rect 126296 630652 580172 630680
rect 126296 630640 126302 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3510 618264 3516 618316
rect 3568 618304 3574 618316
rect 46198 618304 46204 618316
rect 3568 618276 46204 618304
rect 3568 618264 3574 618276
rect 46198 618264 46204 618276
rect 46256 618264 46262 618316
rect 130378 616836 130384 616888
rect 130436 616876 130442 616888
rect 580166 616876 580172 616888
rect 130436 616848 580172 616876
rect 130436 616836 130442 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 2774 605888 2780 605940
rect 2832 605928 2838 605940
rect 4798 605928 4804 605940
rect 2832 605900 4804 605928
rect 2832 605888 2838 605900
rect 4798 605888 4804 605900
rect 4856 605888 4862 605940
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 116578 579680 116584 579692
rect 3384 579652 116584 579680
rect 3384 579640 3390 579652
rect 116578 579640 116584 579652
rect 116636 579640 116642 579692
rect 142798 576852 142804 576904
rect 142856 576892 142862 576904
rect 580166 576892 580172 576904
rect 142856 576864 580172 576892
rect 142856 576852 142862 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3234 565836 3240 565888
rect 3292 565876 3298 565888
rect 64138 565876 64144 565888
rect 3292 565848 64144 565876
rect 3292 565836 3298 565848
rect 64138 565836 64144 565848
rect 64196 565836 64202 565888
rect 102778 563048 102784 563100
rect 102836 563088 102842 563100
rect 579798 563088 579804 563100
rect 102836 563060 579804 563088
rect 102836 563048 102842 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 3326 553392 3332 553444
rect 3384 553432 3390 553444
rect 18598 553432 18604 553444
rect 3384 553404 18604 553432
rect 3384 553392 3390 553404
rect 18598 553392 18604 553404
rect 18656 553392 18662 553444
rect 2958 527144 2964 527196
rect 3016 527184 3022 527196
rect 36538 527184 36544 527196
rect 3016 527156 36544 527184
rect 3016 527144 3022 527156
rect 36538 527144 36544 527156
rect 36596 527144 36602 527196
rect 140038 524424 140044 524476
rect 140096 524464 140102 524476
rect 580166 524464 580172 524476
rect 140096 524436 580172 524464
rect 140096 524424 140102 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3326 500964 3332 501016
rect 3384 501004 3390 501016
rect 100018 501004 100024 501016
rect 3384 500976 100024 501004
rect 3384 500964 3390 500976
rect 100018 500964 100024 500976
rect 100076 500964 100082 501016
rect 129090 484372 129096 484424
rect 129148 484412 129154 484424
rect 580166 484412 580172 484424
rect 129148 484384 580172 484412
rect 129148 484372 129154 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 3050 474716 3056 474768
rect 3108 474756 3114 474768
rect 111058 474756 111064 474768
rect 3108 474728 111064 474756
rect 3108 474716 3114 474728
rect 111058 474716 111064 474728
rect 111116 474716 111122 474768
rect 138658 470568 138664 470620
rect 138716 470608 138722 470620
rect 580166 470608 580172 470620
rect 138716 470580 580172 470608
rect 138716 470568 138722 470580
rect 580166 470568 580172 470580
rect 580224 470568 580230 470620
rect 3326 462340 3332 462392
rect 3384 462380 3390 462392
rect 31018 462380 31024 462392
rect 3384 462352 31024 462380
rect 3384 462340 3390 462352
rect 31018 462340 31024 462352
rect 31076 462340 31082 462392
rect 59170 456764 59176 456816
rect 59228 456804 59234 456816
rect 580166 456804 580172 456816
rect 59228 456776 580172 456804
rect 59228 456764 59234 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 3326 448536 3332 448588
rect 3384 448576 3390 448588
rect 25498 448576 25504 448588
rect 3384 448548 25504 448576
rect 3384 448536 3390 448548
rect 25498 448536 25504 448548
rect 25556 448536 25562 448588
rect 123478 430584 123484 430636
rect 123536 430624 123542 430636
rect 579890 430624 579896 430636
rect 123536 430596 579896 430624
rect 123536 430584 123542 430596
rect 579890 430584 579896 430596
rect 579948 430584 579954 430636
rect 3326 423308 3332 423360
rect 3384 423348 3390 423360
rect 7558 423348 7564 423360
rect 3384 423320 7564 423348
rect 3384 423308 3390 423320
rect 7558 423308 7564 423320
rect 7616 423308 7622 423360
rect 93118 418140 93124 418192
rect 93176 418180 93182 418192
rect 580166 418180 580172 418192
rect 93176 418152 580172 418180
rect 93176 418140 93182 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 3326 409844 3332 409896
rect 3384 409884 3390 409896
rect 17218 409884 17224 409896
rect 3384 409856 17224 409884
rect 3384 409844 3390 409856
rect 17218 409844 17224 409856
rect 17276 409844 17282 409896
rect 67542 404336 67548 404388
rect 67600 404376 67606 404388
rect 580166 404376 580172 404388
rect 67600 404348 580172 404376
rect 67600 404336 67606 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3326 397468 3332 397520
rect 3384 397508 3390 397520
rect 43438 397508 43444 397520
rect 3384 397480 43444 397508
rect 3384 397468 3390 397480
rect 43438 397468 43444 397480
rect 43496 397468 43502 397520
rect 124950 378156 124956 378208
rect 125008 378196 125014 378208
rect 580166 378196 580172 378208
rect 125008 378168 580172 378196
rect 125008 378156 125014 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 3326 371220 3332 371272
rect 3384 371260 3390 371272
rect 50338 371260 50344 371272
rect 3384 371232 50344 371260
rect 3384 371220 3390 371232
rect 50338 371220 50344 371232
rect 50396 371220 50402 371272
rect 130470 364352 130476 364404
rect 130528 364392 130534 364404
rect 579614 364392 579620 364404
rect 130528 364364 579620 364392
rect 130528 364352 130534 364364
rect 579614 364352 579620 364364
rect 579672 364352 579678 364404
rect 3326 357416 3332 357468
rect 3384 357456 3390 357468
rect 13078 357456 13084 357468
rect 3384 357428 13084 357456
rect 3384 357416 3390 357428
rect 13078 357416 13084 357428
rect 13136 357416 13142 357468
rect 80790 351908 80796 351960
rect 80848 351948 80854 351960
rect 580166 351948 580172 351960
rect 80848 351920 580172 351948
rect 80848 351908 80854 351920
rect 580166 351908 580172 351920
rect 580224 351908 580230 351960
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 117958 345080 117964 345092
rect 3384 345052 117964 345080
rect 3384 345040 3390 345052
rect 117958 345040 117964 345052
rect 118016 345040 118022 345092
rect 13078 338716 13084 338768
rect 13136 338756 13142 338768
rect 97994 338756 98000 338768
rect 13136 338728 98000 338756
rect 13136 338716 13142 338728
rect 97994 338716 98000 338728
rect 98052 338716 98058 338768
rect 88334 334568 88340 334620
rect 88392 334608 88398 334620
rect 103790 334608 103796 334620
rect 88392 334580 103796 334608
rect 88392 334568 88398 334580
rect 103790 334568 103796 334580
rect 103848 334568 103854 334620
rect 3418 326340 3424 326392
rect 3476 326380 3482 326392
rect 120166 326380 120172 326392
rect 3476 326352 120172 326380
rect 3476 326340 3482 326352
rect 120166 326340 120172 326352
rect 120224 326340 120230 326392
rect 123570 324300 123576 324352
rect 123628 324340 123634 324352
rect 580166 324340 580172 324352
rect 123628 324312 580172 324340
rect 123628 324300 123634 324312
rect 580166 324300 580172 324312
rect 580224 324300 580230 324352
rect 68922 323552 68928 323604
rect 68980 323592 68986 323604
rect 269758 323592 269764 323604
rect 68980 323564 269764 323592
rect 68980 323552 68986 323564
rect 269758 323552 269764 323564
rect 269816 323552 269822 323604
rect 111058 322192 111064 322244
rect 111116 322232 111122 322244
rect 121454 322232 121460 322244
rect 111116 322204 121460 322232
rect 111116 322192 111122 322204
rect 121454 322192 121460 322204
rect 121512 322192 121518 322244
rect 91094 319404 91100 319456
rect 91152 319444 91158 319456
rect 148318 319444 148324 319456
rect 91152 319416 148324 319444
rect 91152 319404 91158 319416
rect 148318 319404 148324 319416
rect 148376 319404 148382 319456
rect 3326 318792 3332 318844
rect 3384 318832 3390 318844
rect 22094 318832 22100 318844
rect 3384 318804 22100 318832
rect 3384 318792 3390 318804
rect 22094 318792 22100 318804
rect 22152 318792 22158 318844
rect 22094 318044 22100 318096
rect 22152 318084 22158 318096
rect 115934 318084 115940 318096
rect 22152 318056 115940 318084
rect 22152 318044 22158 318056
rect 115934 318044 115940 318056
rect 115992 318044 115998 318096
rect 93946 317500 93952 317552
rect 94004 317540 94010 317552
rect 102778 317540 102784 317552
rect 94004 317512 102784 317540
rect 94004 317500 94010 317512
rect 102778 317500 102784 317512
rect 102836 317500 102842 317552
rect 77294 315256 77300 315308
rect 77352 315296 77358 315308
rect 93118 315296 93124 315308
rect 77352 315268 93124 315296
rect 77352 315256 77358 315268
rect 93118 315256 93124 315268
rect 93176 315256 93182 315308
rect 3510 313896 3516 313948
rect 3568 313936 3574 313948
rect 120074 313936 120080 313948
rect 3568 313908 120080 313936
rect 3568 313896 3574 313908
rect 120074 313896 120080 313908
rect 120132 313896 120138 313948
rect 125134 313896 125140 313948
rect 125192 313936 125198 313948
rect 282914 313936 282920 313948
rect 125192 313908 282920 313936
rect 125192 313896 125198 313908
rect 282914 313896 282920 313908
rect 282972 313896 282978 313948
rect 4798 312536 4804 312588
rect 4856 312576 4862 312588
rect 94130 312576 94136 312588
rect 4856 312548 94136 312576
rect 4856 312536 4862 312548
rect 94130 312536 94136 312548
rect 94188 312536 94194 312588
rect 100018 312536 100024 312588
rect 100076 312576 100082 312588
rect 121546 312576 121552 312588
rect 100076 312548 121552 312576
rect 100076 312536 100082 312548
rect 121546 312536 121552 312548
rect 121604 312536 121610 312588
rect 126330 311856 126336 311908
rect 126388 311896 126394 311908
rect 580166 311896 580172 311908
rect 126388 311868 580172 311896
rect 126388 311856 126394 311868
rect 580166 311856 580172 311868
rect 580224 311856 580230 311908
rect 69106 311108 69112 311160
rect 69164 311148 69170 311160
rect 153194 311148 153200 311160
rect 69164 311120 153200 311148
rect 69164 311108 69170 311120
rect 153194 311108 153200 311120
rect 153252 311108 153258 311160
rect 39298 309748 39304 309800
rect 39356 309788 39362 309800
rect 121638 309788 121644 309800
rect 39356 309760 121644 309788
rect 39356 309748 39362 309760
rect 121638 309748 121644 309760
rect 121696 309748 121702 309800
rect 71774 308388 71780 308440
rect 71832 308428 71838 308440
rect 114554 308428 114560 308440
rect 71832 308400 114560 308428
rect 71832 308388 71838 308400
rect 114554 308388 114560 308400
rect 114612 308388 114618 308440
rect 98086 307776 98092 307828
rect 98144 307816 98150 307828
rect 283558 307816 283564 307828
rect 98144 307788 283564 307816
rect 98144 307776 98150 307788
rect 283558 307776 283564 307788
rect 283616 307776 283622 307828
rect 69014 307028 69020 307080
rect 69072 307068 69078 307080
rect 580258 307068 580264 307080
rect 69072 307040 580264 307068
rect 69072 307028 69078 307040
rect 580258 307028 580264 307040
rect 580316 307028 580322 307080
rect 75914 306348 75920 306400
rect 75972 306388 75978 306400
rect 342254 306388 342260 306400
rect 75972 306360 342260 306388
rect 75972 306348 75978 306360
rect 342254 306348 342260 306360
rect 342312 306348 342318 306400
rect 123662 305600 123668 305652
rect 123720 305640 123726 305652
rect 201494 305640 201500 305652
rect 123720 305612 201500 305640
rect 123720 305600 123726 305612
rect 201494 305600 201500 305612
rect 201552 305600 201558 305652
rect 3418 305056 3424 305108
rect 3476 305096 3482 305108
rect 119798 305096 119804 305108
rect 3476 305068 119804 305096
rect 3476 305056 3482 305068
rect 119798 305056 119804 305068
rect 119856 305056 119862 305108
rect 112438 304988 112444 305040
rect 112496 305028 112502 305040
rect 281534 305028 281540 305040
rect 112496 305000 281540 305028
rect 112496 304988 112502 305000
rect 281534 304988 281540 305000
rect 281592 304988 281598 305040
rect 102134 303764 102140 303816
rect 102192 303804 102198 303816
rect 185578 303804 185584 303816
rect 102192 303776 185584 303804
rect 102192 303764 102198 303776
rect 185578 303764 185584 303776
rect 185636 303764 185642 303816
rect 102410 303696 102416 303748
rect 102468 303736 102474 303748
rect 224218 303736 224224 303748
rect 102468 303708 224224 303736
rect 102468 303696 102474 303708
rect 224218 303696 224224 303708
rect 224276 303696 224282 303748
rect 90266 303628 90272 303680
rect 90324 303668 90330 303680
rect 278774 303668 278780 303680
rect 90324 303640 278780 303668
rect 90324 303628 90330 303640
rect 278774 303628 278780 303640
rect 278832 303628 278838 303680
rect 82078 303560 82084 303612
rect 82136 303600 82142 303612
rect 84470 303600 84476 303612
rect 82136 303572 84476 303600
rect 82136 303560 82142 303572
rect 84470 303560 84476 303572
rect 84528 303560 84534 303612
rect 79226 302268 79232 302320
rect 79284 302308 79290 302320
rect 189718 302308 189724 302320
rect 79284 302280 189724 302308
rect 79284 302268 79290 302280
rect 189718 302268 189724 302280
rect 189776 302268 189782 302320
rect 112162 302200 112168 302252
rect 112220 302240 112226 302252
rect 273254 302240 273260 302252
rect 112220 302212 273260 302240
rect 112220 302200 112226 302212
rect 273254 302200 273260 302212
rect 273312 302200 273318 302252
rect 117958 301520 117964 301572
rect 118016 301560 118022 301572
rect 119154 301560 119160 301572
rect 118016 301532 119160 301560
rect 118016 301520 118022 301532
rect 119154 301520 119160 301532
rect 119212 301520 119218 301572
rect 25498 301452 25504 301504
rect 25556 301492 25562 301504
rect 70946 301492 70952 301504
rect 25556 301464 70952 301492
rect 25556 301452 25562 301464
rect 70946 301452 70952 301464
rect 71004 301452 71010 301504
rect 73522 301452 73528 301504
rect 73580 301492 73586 301504
rect 80790 301492 80796 301504
rect 73580 301464 80796 301492
rect 73580 301452 73586 301464
rect 80790 301452 80796 301464
rect 80848 301452 80854 301504
rect 67450 300908 67456 300960
rect 67508 300948 67514 300960
rect 152458 300948 152464 300960
rect 67508 300920 152464 300948
rect 67508 300908 67514 300920
rect 152458 300908 152464 300920
rect 152516 300908 152522 300960
rect 86402 300840 86408 300892
rect 86460 300880 86466 300892
rect 319438 300880 319444 300892
rect 86460 300852 319444 300880
rect 86460 300840 86466 300852
rect 319438 300840 319444 300852
rect 319496 300840 319502 300892
rect 110414 299684 110420 299736
rect 110472 299724 110478 299736
rect 184198 299724 184204 299736
rect 110472 299696 184204 299724
rect 110472 299684 110478 299696
rect 184198 299684 184204 299696
rect 184256 299684 184262 299736
rect 87690 299616 87696 299668
rect 87748 299656 87754 299668
rect 225598 299656 225604 299668
rect 87748 299628 225604 299656
rect 87748 299616 87754 299628
rect 225598 299616 225604 299628
rect 225656 299616 225662 299668
rect 68738 299548 68744 299600
rect 68796 299588 68802 299600
rect 308398 299588 308404 299600
rect 68796 299560 308404 299588
rect 68796 299548 68802 299560
rect 308398 299548 308404 299560
rect 308456 299548 308462 299600
rect 71774 299480 71780 299532
rect 71832 299520 71838 299532
rect 343634 299520 343640 299532
rect 71832 299492 343640 299520
rect 71832 299480 71838 299492
rect 343634 299480 343640 299492
rect 343692 299480 343698 299532
rect 7558 298732 7564 298784
rect 7616 298772 7622 298784
rect 72602 298772 72608 298784
rect 7616 298744 72608 298772
rect 7616 298732 7622 298744
rect 72602 298732 72608 298744
rect 72660 298732 72666 298784
rect 89990 298460 89996 298512
rect 90048 298500 90054 298512
rect 166258 298500 166264 298512
rect 90048 298472 166264 298500
rect 90048 298460 90054 298472
rect 166258 298460 166264 298472
rect 166316 298460 166322 298512
rect 93210 298392 93216 298444
rect 93268 298432 93274 298444
rect 174538 298432 174544 298444
rect 93268 298404 174544 298432
rect 93268 298392 93274 298404
rect 174538 298392 174544 298404
rect 174596 298392 174602 298444
rect 74534 298324 74540 298376
rect 74592 298364 74598 298376
rect 192478 298364 192484 298376
rect 74592 298336 192484 298364
rect 74592 298324 74598 298336
rect 192478 298324 192484 298336
rect 192536 298324 192542 298376
rect 75178 298256 75184 298308
rect 75236 298296 75242 298308
rect 274634 298296 274640 298308
rect 75236 298268 274640 298296
rect 75236 298256 75242 298268
rect 274634 298256 274640 298268
rect 274692 298256 274698 298308
rect 81618 298188 81624 298240
rect 81676 298228 81682 298240
rect 333974 298228 333980 298240
rect 81676 298200 333980 298228
rect 81676 298188 81682 298200
rect 333974 298188 333980 298200
rect 334032 298188 334038 298240
rect 106090 298120 106096 298172
rect 106148 298160 106154 298172
rect 582558 298160 582564 298172
rect 106148 298132 582564 298160
rect 106148 298120 106154 298132
rect 582558 298120 582564 298132
rect 582616 298120 582622 298172
rect 114462 297032 114468 297084
rect 114520 297072 114526 297084
rect 160738 297072 160744 297084
rect 114520 297044 160744 297072
rect 114520 297032 114526 297044
rect 160738 297032 160744 297044
rect 160796 297032 160802 297084
rect 86126 296964 86132 297016
rect 86184 297004 86190 297016
rect 210418 297004 210424 297016
rect 86184 296976 210424 297004
rect 86184 296964 86190 296976
rect 210418 296964 210424 296976
rect 210476 296964 210482 297016
rect 70026 296896 70032 296948
rect 70084 296936 70090 296948
rect 248414 296936 248420 296948
rect 70084 296908 248420 296936
rect 70084 296896 70090 296908
rect 248414 296896 248420 296908
rect 248472 296896 248478 296948
rect 89346 296828 89352 296880
rect 89404 296868 89410 296880
rect 339494 296868 339500 296880
rect 89404 296840 339500 296868
rect 89404 296828 89410 296840
rect 339494 296828 339500 296840
rect 339552 296828 339558 296880
rect 88702 296760 88708 296812
rect 88760 296800 88766 296812
rect 340874 296800 340880 296812
rect 88760 296772 340880 296800
rect 88760 296760 88766 296772
rect 340874 296760 340880 296772
rect 340932 296760 340938 296812
rect 70670 296692 70676 296744
rect 70728 296732 70734 296744
rect 325786 296732 325792 296744
rect 70728 296704 325792 296732
rect 70728 296692 70734 296704
rect 325786 296692 325792 296704
rect 325844 296692 325850 296744
rect 111242 295672 111248 295724
rect 111300 295712 111306 295724
rect 157978 295712 157984 295724
rect 111300 295684 157984 295712
rect 111300 295672 111306 295684
rect 157978 295672 157984 295684
rect 158036 295672 158042 295724
rect 77110 295604 77116 295656
rect 77168 295644 77174 295656
rect 126422 295644 126428 295656
rect 77168 295616 126428 295644
rect 77168 295604 77174 295616
rect 126422 295604 126428 295616
rect 126480 295604 126486 295656
rect 82262 295536 82268 295588
rect 82320 295576 82326 295588
rect 178678 295576 178684 295588
rect 82320 295548 178684 295576
rect 82320 295536 82326 295548
rect 178678 295536 178684 295548
rect 178736 295536 178742 295588
rect 84194 295468 84200 295520
rect 84252 295508 84258 295520
rect 196618 295508 196624 295520
rect 84252 295480 196624 295508
rect 84252 295468 84258 295480
rect 196618 295468 196624 295480
rect 196676 295468 196682 295520
rect 68554 295400 68560 295452
rect 68612 295440 68618 295452
rect 278038 295440 278044 295452
rect 68612 295412 278044 295440
rect 68612 295400 68618 295412
rect 278038 295400 278044 295412
rect 278096 295400 278102 295452
rect 109954 295332 109960 295384
rect 110012 295372 110018 295384
rect 347038 295372 347044 295384
rect 110012 295344 347044 295372
rect 110012 295332 110018 295344
rect 347038 295332 347044 295344
rect 347096 295332 347102 295384
rect 87414 294652 87420 294704
rect 87472 294692 87478 294704
rect 112438 294692 112444 294704
rect 87472 294664 112444 294692
rect 87472 294652 87478 294664
rect 112438 294652 112444 294664
rect 112496 294652 112502 294704
rect 73246 294584 73252 294636
rect 73304 294624 73310 294636
rect 111794 294624 111800 294636
rect 73304 294596 111800 294624
rect 73304 294584 73310 294596
rect 111794 294584 111800 294596
rect 111852 294584 111858 294636
rect 113818 294380 113824 294432
rect 113876 294420 113882 294432
rect 118418 294420 118424 294432
rect 113876 294392 118424 294420
rect 113876 294380 113882 294392
rect 118418 294380 118424 294392
rect 118476 294380 118482 294432
rect 106734 294312 106740 294364
rect 106792 294352 106798 294364
rect 170398 294352 170404 294364
rect 106792 294324 170404 294352
rect 106792 294312 106798 294324
rect 170398 294312 170404 294324
rect 170456 294312 170462 294364
rect 91922 294244 91928 294296
rect 91980 294284 91986 294296
rect 215938 294284 215944 294296
rect 91980 294256 215944 294284
rect 91980 294244 91986 294256
rect 215938 294244 215944 294256
rect 215996 294244 216002 294296
rect 82906 294176 82912 294228
rect 82964 294216 82970 294228
rect 255314 294216 255320 294228
rect 82964 294188 255320 294216
rect 82964 294176 82970 294188
rect 255314 294176 255320 294188
rect 255372 294176 255378 294228
rect 32398 294108 32404 294160
rect 32456 294148 32462 294160
rect 32456 294120 103514 294148
rect 32456 294108 32462 294120
rect 69474 294040 69480 294092
rect 69532 294080 69538 294092
rect 92566 294080 92572 294092
rect 69532 294052 92572 294080
rect 69532 294040 69538 294052
rect 92566 294040 92572 294052
rect 92624 294040 92630 294092
rect 103486 294080 103514 294120
rect 117682 294108 117688 294160
rect 117740 294148 117746 294160
rect 308490 294148 308496 294160
rect 117740 294120 308496 294148
rect 117740 294108 117746 294120
rect 308490 294108 308496 294120
rect 308548 294108 308554 294160
rect 118326 294080 118332 294092
rect 103486 294052 118332 294080
rect 118326 294040 118332 294052
rect 118384 294040 118390 294092
rect 118418 294040 118424 294092
rect 118476 294080 118482 294092
rect 345014 294080 345020 294092
rect 118476 294052 345020 294080
rect 118476 294040 118482 294052
rect 345014 294040 345020 294052
rect 345072 294040 345078 294092
rect 39298 293972 39304 294024
rect 39356 294012 39362 294024
rect 39356 293984 77708 294012
rect 39356 293972 39362 293984
rect 77680 293944 77708 293984
rect 77754 293972 77760 294024
rect 77812 294012 77818 294024
rect 80698 294012 80704 294024
rect 77812 293984 80704 294012
rect 77812 293972 77818 293984
rect 80698 293972 80704 293984
rect 80756 293972 80762 294024
rect 84286 293972 84292 294024
rect 84344 294012 84350 294024
rect 85206 294012 85212 294024
rect 84344 293984 85212 294012
rect 84344 293972 84350 293984
rect 85206 293972 85212 293984
rect 85264 293972 85270 294024
rect 93946 293972 93952 294024
rect 94004 294012 94010 294024
rect 94774 294012 94780 294024
rect 94004 293984 94780 294012
rect 94004 293972 94010 293984
rect 94774 293972 94780 293984
rect 94832 293972 94838 294024
rect 111886 293972 111892 294024
rect 111944 294012 111950 294024
rect 350534 294012 350540 294024
rect 111944 293984 350540 294012
rect 111944 293972 111950 293984
rect 350534 293972 350540 293984
rect 350592 293972 350598 294024
rect 78766 293944 78772 293956
rect 77680 293916 78772 293944
rect 78766 293904 78772 293916
rect 78824 293904 78830 293956
rect 93854 292884 93860 292936
rect 93912 292924 93918 292936
rect 120258 292924 120264 292936
rect 93912 292896 120264 292924
rect 93912 292884 93918 292896
rect 120258 292884 120264 292896
rect 120316 292884 120322 292936
rect 2774 292816 2780 292868
rect 2832 292856 2838 292868
rect 4798 292856 4804 292868
rect 2832 292828 4804 292856
rect 2832 292816 2838 292828
rect 4798 292816 4804 292828
rect 4856 292816 4862 292868
rect 83550 292816 83556 292868
rect 83608 292856 83614 292868
rect 220078 292856 220084 292868
rect 83608 292828 220084 292856
rect 83608 292816 83614 292828
rect 220078 292816 220084 292828
rect 220136 292816 220142 292868
rect 100938 292748 100944 292800
rect 100996 292788 101002 292800
rect 263594 292788 263600 292800
rect 100996 292760 263600 292788
rect 100996 292748 101002 292760
rect 263594 292748 263600 292760
rect 263652 292748 263658 292800
rect 103514 292680 103520 292732
rect 103572 292720 103578 292732
rect 318058 292720 318064 292732
rect 103572 292692 318064 292720
rect 103572 292680 103578 292692
rect 318058 292680 318064 292692
rect 318116 292680 318122 292732
rect 48958 292612 48964 292664
rect 49016 292652 49022 292664
rect 97074 292652 97080 292664
rect 49016 292624 97080 292652
rect 49016 292612 49022 292624
rect 97074 292612 97080 292624
rect 97132 292612 97138 292664
rect 97718 292612 97724 292664
rect 97776 292652 97782 292664
rect 320174 292652 320180 292664
rect 97776 292624 320180 292652
rect 97776 292612 97782 292624
rect 320174 292612 320180 292624
rect 320232 292612 320238 292664
rect 8202 292544 8208 292596
rect 8260 292584 8266 292596
rect 96430 292584 96436 292596
rect 8260 292556 96436 292584
rect 8260 292544 8266 292556
rect 96430 292544 96436 292556
rect 96488 292544 96494 292596
rect 109310 292544 109316 292596
rect 109368 292584 109374 292596
rect 336734 292584 336740 292596
rect 109368 292556 336740 292584
rect 109368 292544 109374 292556
rect 336734 292544 336740 292556
rect 336792 292544 336798 292596
rect 115842 291864 115848 291916
rect 115900 291864 115906 291916
rect 117222 291864 117228 291916
rect 117280 291864 117286 291916
rect 119062 291864 119068 291916
rect 119120 291904 119126 291916
rect 119890 291904 119896 291916
rect 119120 291876 119896 291904
rect 119120 291864 119126 291876
rect 119890 291864 119896 291876
rect 119948 291864 119954 291916
rect 3418 291796 3424 291848
rect 3476 291836 3482 291848
rect 69474 291836 69480 291848
rect 3476 291808 69480 291836
rect 3476 291796 3482 291808
rect 69474 291796 69480 291808
rect 69532 291796 69538 291848
rect 115860 291292 115888 291864
rect 117240 291360 117268 291864
rect 148318 291360 148324 291372
rect 117240 291332 148324 291360
rect 148318 291320 148324 291332
rect 148376 291320 148382 291372
rect 345106 291292 345112 291304
rect 115860 291264 345112 291292
rect 345106 291252 345112 291264
rect 345164 291252 345170 291304
rect 69750 291184 69756 291236
rect 69808 291224 69814 291236
rect 582650 291224 582656 291236
rect 69808 291196 582656 291224
rect 69808 291184 69814 291196
rect 582650 291184 582656 291196
rect 582708 291184 582714 291236
rect 121638 289892 121644 289944
rect 121696 289932 121702 289944
rect 246298 289932 246304 289944
rect 121696 289904 246304 289932
rect 121696 289892 121702 289904
rect 246298 289892 246304 289904
rect 246356 289892 246362 289944
rect 25498 289824 25504 289876
rect 25556 289864 25562 289876
rect 67634 289864 67640 289876
rect 25556 289836 67640 289864
rect 25556 289824 25562 289836
rect 67634 289824 67640 289836
rect 67692 289824 67698 289876
rect 121730 289824 121736 289876
rect 121788 289864 121794 289876
rect 269114 289864 269120 289876
rect 121788 289836 269120 289864
rect 121788 289824 121794 289836
rect 269114 289824 269120 289836
rect 269172 289824 269178 289876
rect 121638 289756 121644 289808
rect 121696 289796 121702 289808
rect 124950 289796 124956 289808
rect 121696 289768 124956 289796
rect 121696 289756 121702 289768
rect 124950 289756 124956 289768
rect 125008 289756 125014 289808
rect 68554 289484 68560 289536
rect 68612 289524 68618 289536
rect 68922 289524 68928 289536
rect 68612 289496 68928 289524
rect 68612 289484 68618 289496
rect 68922 289484 68928 289496
rect 68980 289484 68986 289536
rect 120258 289076 120264 289128
rect 120316 289116 120322 289128
rect 202138 289116 202144 289128
rect 120316 289088 202144 289116
rect 120316 289076 120322 289088
rect 202138 289076 202144 289088
rect 202196 289076 202202 289128
rect 66070 288396 66076 288448
rect 66128 288436 66134 288448
rect 68186 288436 68192 288448
rect 66128 288408 68192 288436
rect 66128 288396 66134 288408
rect 68186 288396 68192 288408
rect 68244 288396 68250 288448
rect 121638 288396 121644 288448
rect 121696 288436 121702 288448
rect 313918 288436 313924 288448
rect 121696 288408 313924 288436
rect 121696 288396 121702 288408
rect 313918 288396 313924 288408
rect 313976 288396 313982 288448
rect 55030 287036 55036 287088
rect 55088 287076 55094 287088
rect 67634 287076 67640 287088
rect 55088 287048 67640 287076
rect 55088 287036 55094 287048
rect 67634 287036 67640 287048
rect 67692 287036 67698 287088
rect 121638 286968 121644 287020
rect 121696 287008 121702 287020
rect 123662 287008 123668 287020
rect 121696 286980 123668 287008
rect 121696 286968 121702 286980
rect 123662 286968 123668 286980
rect 123720 286968 123726 287020
rect 26878 286900 26884 286952
rect 26936 286940 26942 286952
rect 67634 286940 67640 286952
rect 26936 286912 67640 286940
rect 26936 286900 26942 286912
rect 67634 286900 67640 286912
rect 67692 286900 67698 286952
rect 121822 286288 121828 286340
rect 121880 286328 121886 286340
rect 327074 286328 327080 286340
rect 121880 286300 327080 286328
rect 121880 286288 121886 286300
rect 327074 286288 327080 286300
rect 327132 286288 327138 286340
rect 60642 285676 60648 285728
rect 60700 285716 60706 285728
rect 67726 285716 67732 285728
rect 60700 285688 67732 285716
rect 60700 285676 60706 285688
rect 67726 285676 67732 285688
rect 67784 285676 67790 285728
rect 121546 285676 121552 285728
rect 121604 285716 121610 285728
rect 193122 285716 193128 285728
rect 121604 285688 193128 285716
rect 121604 285676 121610 285688
rect 193122 285676 193128 285688
rect 193180 285676 193186 285728
rect 121638 285608 121644 285660
rect 121696 285648 121702 285660
rect 138658 285648 138664 285660
rect 121696 285620 138664 285648
rect 121696 285608 121702 285620
rect 138658 285608 138664 285620
rect 138716 285608 138722 285660
rect 52362 284316 52368 284368
rect 52420 284356 52426 284368
rect 67634 284356 67640 284368
rect 52420 284328 67640 284356
rect 52420 284316 52426 284328
rect 67634 284316 67640 284328
rect 67692 284316 67698 284368
rect 121546 284316 121552 284368
rect 121604 284356 121610 284368
rect 335354 284356 335360 284368
rect 121604 284328 335360 284356
rect 121604 284316 121610 284328
rect 335354 284316 335360 284328
rect 335412 284316 335418 284368
rect 121546 284112 121552 284164
rect 121604 284152 121610 284164
rect 124858 284152 124864 284164
rect 121604 284124 124864 284152
rect 121604 284112 121610 284124
rect 124858 284112 124864 284124
rect 124916 284112 124922 284164
rect 121546 282888 121552 282940
rect 121604 282928 121610 282940
rect 307018 282928 307024 282940
rect 121604 282900 307024 282928
rect 121604 282888 121610 282900
rect 307018 282888 307024 282900
rect 307076 282888 307082 282940
rect 193122 282140 193128 282192
rect 193180 282180 193186 282192
rect 580258 282180 580264 282192
rect 193180 282152 580264 282180
rect 193180 282140 193186 282152
rect 580258 282140 580264 282152
rect 580316 282140 580322 282192
rect 121546 281528 121552 281580
rect 121604 281568 121610 281580
rect 242158 281568 242164 281580
rect 121604 281540 242164 281568
rect 121604 281528 121610 281540
rect 242158 281528 242164 281540
rect 242216 281528 242222 281580
rect 121546 280236 121552 280288
rect 121604 280276 121610 280288
rect 238018 280276 238024 280288
rect 121604 280248 238024 280276
rect 121604 280236 121610 280248
rect 238018 280236 238024 280248
rect 238076 280236 238082 280288
rect 46842 280168 46848 280220
rect 46900 280208 46906 280220
rect 67634 280208 67640 280220
rect 46900 280180 67640 280208
rect 46900 280168 46906 280180
rect 67634 280168 67640 280180
rect 67692 280168 67698 280220
rect 121638 280168 121644 280220
rect 121696 280208 121702 280220
rect 342346 280208 342352 280220
rect 121696 280180 342352 280208
rect 121696 280168 121702 280180
rect 342346 280168 342352 280180
rect 342404 280168 342410 280220
rect 121546 278808 121552 278860
rect 121604 278848 121610 278860
rect 206278 278848 206284 278860
rect 121604 278820 206284 278848
rect 121604 278808 121610 278820
rect 206278 278808 206284 278820
rect 206336 278808 206342 278860
rect 57238 278740 57244 278792
rect 57296 278780 57302 278792
rect 67634 278780 67640 278792
rect 57296 278752 67640 278780
rect 57296 278740 57302 278752
rect 67634 278740 67640 278752
rect 67692 278740 67698 278792
rect 121638 278740 121644 278792
rect 121696 278780 121702 278792
rect 318150 278780 318156 278792
rect 121696 278752 318156 278780
rect 121696 278740 121702 278752
rect 318150 278740 318156 278752
rect 318208 278740 318214 278792
rect 56502 277448 56508 277500
rect 56560 277488 56566 277500
rect 67634 277488 67640 277500
rect 56560 277460 67640 277488
rect 56560 277448 56566 277460
rect 67634 277448 67640 277460
rect 67692 277448 67698 277500
rect 121638 277448 121644 277500
rect 121696 277488 121702 277500
rect 328454 277488 328460 277500
rect 121696 277460 328460 277488
rect 121696 277448 121702 277460
rect 328454 277448 328460 277460
rect 328512 277448 328518 277500
rect 50890 277380 50896 277432
rect 50948 277420 50954 277432
rect 67726 277420 67732 277432
rect 50948 277392 67732 277420
rect 50948 277380 50954 277392
rect 67726 277380 67732 277392
rect 67784 277380 67790 277432
rect 121546 277380 121552 277432
rect 121604 277420 121610 277432
rect 347774 277420 347780 277432
rect 121604 277392 347780 277420
rect 121604 277380 121610 277392
rect 347774 277380 347780 277392
rect 347832 277380 347838 277432
rect 53650 276088 53656 276140
rect 53708 276128 53714 276140
rect 67726 276128 67732 276140
rect 53708 276100 67732 276128
rect 53708 276088 53714 276100
rect 67726 276088 67732 276100
rect 67784 276088 67790 276140
rect 121638 276088 121644 276140
rect 121696 276128 121702 276140
rect 247678 276128 247684 276140
rect 121696 276100 247684 276128
rect 121696 276088 121702 276100
rect 247678 276088 247684 276100
rect 247736 276088 247742 276140
rect 45462 276020 45468 276072
rect 45520 276060 45526 276072
rect 67634 276060 67640 276072
rect 45520 276032 67640 276060
rect 45520 276020 45526 276032
rect 67634 276020 67640 276032
rect 67692 276020 67698 276072
rect 121546 276020 121552 276072
rect 121604 276060 121610 276072
rect 331214 276060 331220 276072
rect 121604 276032 331220 276060
rect 121604 276020 121610 276032
rect 331214 276020 331220 276032
rect 331272 276020 331278 276072
rect 122190 275272 122196 275324
rect 122248 275312 122254 275324
rect 392578 275312 392584 275324
rect 122248 275284 392584 275312
rect 122248 275272 122254 275284
rect 392578 275272 392584 275284
rect 392636 275272 392642 275324
rect 61930 274728 61936 274780
rect 61988 274768 61994 274780
rect 67634 274768 67640 274780
rect 61988 274740 67640 274768
rect 61988 274728 61994 274740
rect 67634 274728 67640 274740
rect 67692 274728 67698 274780
rect 48222 274660 48228 274712
rect 48280 274700 48286 274712
rect 67726 274700 67732 274712
rect 48280 274672 67732 274700
rect 48280 274660 48286 274672
rect 67726 274660 67732 274672
rect 67784 274660 67790 274712
rect 121546 274660 121552 274712
rect 121604 274700 121610 274712
rect 253934 274700 253940 274712
rect 121604 274672 253940 274700
rect 121604 274660 121610 274672
rect 253934 274660 253940 274672
rect 253992 274660 253998 274712
rect 46198 274592 46204 274644
rect 46256 274632 46262 274644
rect 67634 274632 67640 274644
rect 46256 274604 67640 274632
rect 46256 274592 46262 274604
rect 67634 274592 67640 274604
rect 67692 274592 67698 274644
rect 121638 274592 121644 274644
rect 121696 274632 121702 274644
rect 126330 274632 126336 274644
rect 121696 274604 126336 274632
rect 121696 274592 121702 274604
rect 126330 274592 126336 274604
rect 126388 274592 126394 274644
rect 66162 273232 66168 273284
rect 66220 273272 66226 273284
rect 68002 273272 68008 273284
rect 66220 273244 68008 273272
rect 66220 273232 66226 273244
rect 68002 273232 68008 273244
rect 68060 273232 68066 273284
rect 121546 273232 121552 273284
rect 121604 273272 121610 273284
rect 211798 273272 211804 273284
rect 121604 273244 211804 273272
rect 121604 273232 121610 273244
rect 211798 273232 211804 273244
rect 211856 273232 211862 273284
rect 121638 273164 121644 273216
rect 121696 273204 121702 273216
rect 126974 273204 126980 273216
rect 121696 273176 126980 273204
rect 121696 273164 121702 273176
rect 126974 273164 126980 273176
rect 127032 273164 127038 273216
rect 121730 272484 121736 272536
rect 121788 272524 121794 272536
rect 395338 272524 395344 272536
rect 121788 272496 395344 272524
rect 121788 272484 121794 272496
rect 395338 272484 395344 272496
rect 395396 272484 395402 272536
rect 64506 271940 64512 271992
rect 64564 271980 64570 271992
rect 67634 271980 67640 271992
rect 64564 271952 67640 271980
rect 64564 271940 64570 271952
rect 67634 271940 67640 271952
rect 67692 271940 67698 271992
rect 57698 271872 57704 271924
rect 57756 271912 57762 271924
rect 67818 271912 67824 271924
rect 57756 271884 67824 271912
rect 57756 271872 57762 271884
rect 67818 271872 67824 271884
rect 67876 271872 67882 271924
rect 57882 271804 57888 271856
rect 57940 271844 57946 271856
rect 67726 271844 67732 271856
rect 57940 271816 67732 271844
rect 57940 271804 57946 271816
rect 67726 271804 67732 271816
rect 67784 271804 67790 271856
rect 54938 270512 54944 270564
rect 54996 270552 55002 270564
rect 67634 270552 67640 270564
rect 54996 270524 67640 270552
rect 54996 270512 55002 270524
rect 67634 270512 67640 270524
rect 67692 270512 67698 270564
rect 121546 270512 121552 270564
rect 121604 270552 121610 270564
rect 249794 270552 249800 270564
rect 121604 270524 249800 270552
rect 121604 270512 121610 270524
rect 249794 270512 249800 270524
rect 249852 270512 249858 270564
rect 121638 269152 121644 269204
rect 121696 269192 121702 269204
rect 207658 269192 207664 269204
rect 121696 269164 207664 269192
rect 121696 269152 121702 269164
rect 207658 269152 207664 269164
rect 207716 269152 207722 269204
rect 60550 269084 60556 269136
rect 60608 269124 60614 269136
rect 67634 269124 67640 269136
rect 60608 269096 67640 269124
rect 60608 269084 60614 269096
rect 67634 269084 67640 269096
rect 67692 269084 67698 269136
rect 121546 269084 121552 269136
rect 121604 269124 121610 269136
rect 239398 269124 239404 269136
rect 121604 269096 239404 269124
rect 121604 269084 121610 269096
rect 239398 269084 239404 269096
rect 239456 269084 239462 269136
rect 46198 267724 46204 267776
rect 46256 267764 46262 267776
rect 67634 267764 67640 267776
rect 46256 267736 67640 267764
rect 46256 267724 46262 267736
rect 67634 267724 67640 267736
rect 67692 267724 67698 267776
rect 121546 267724 121552 267776
rect 121604 267764 121610 267776
rect 311158 267764 311164 267776
rect 121604 267736 311164 267764
rect 121604 267724 121610 267736
rect 311158 267724 311164 267736
rect 311216 267724 311222 267776
rect 8938 267656 8944 267708
rect 8996 267696 9002 267708
rect 67726 267696 67732 267708
rect 8996 267668 67732 267696
rect 8996 267656 9002 267668
rect 67726 267656 67732 267668
rect 67784 267656 67790 267708
rect 64138 267588 64144 267640
rect 64196 267628 64202 267640
rect 67634 267628 67640 267640
rect 64196 267600 67640 267628
rect 64196 267588 64202 267600
rect 67634 267588 67640 267600
rect 67692 267588 67698 267640
rect 122098 266976 122104 267028
rect 122156 267016 122162 267028
rect 255406 267016 255412 267028
rect 122156 266988 255412 267016
rect 122156 266976 122162 266988
rect 255406 266976 255412 266988
rect 255464 266976 255470 267028
rect 121454 266364 121460 266416
rect 121512 266404 121518 266416
rect 345106 266404 345112 266416
rect 121512 266376 345112 266404
rect 121512 266364 121518 266376
rect 345106 266364 345112 266376
rect 345164 266364 345170 266416
rect 21358 266296 21364 266348
rect 21416 266336 21422 266348
rect 67634 266336 67640 266348
rect 21416 266308 67640 266336
rect 21416 266296 21422 266308
rect 67634 266296 67640 266308
rect 67692 266296 67698 266348
rect 57790 265616 57796 265668
rect 57848 265656 57854 265668
rect 68370 265656 68376 265668
rect 57848 265628 68376 265656
rect 57848 265616 57854 265628
rect 68370 265616 68376 265628
rect 68428 265616 68434 265668
rect 121454 265004 121460 265056
rect 121512 265044 121518 265056
rect 308582 265044 308588 265056
rect 121512 265016 308588 265044
rect 121512 265004 121518 265016
rect 308582 265004 308588 265016
rect 308640 265004 308646 265056
rect 121546 264936 121552 264988
rect 121604 264976 121610 264988
rect 349154 264976 349160 264988
rect 121604 264948 349160 264976
rect 121604 264936 121610 264948
rect 349154 264936 349160 264948
rect 349212 264936 349218 264988
rect 121454 264868 121460 264920
rect 121512 264908 121518 264920
rect 129090 264908 129096 264920
rect 121512 264880 129096 264908
rect 121512 264868 121518 264880
rect 129090 264868 129096 264880
rect 129148 264868 129154 264920
rect 56410 263644 56416 263696
rect 56468 263684 56474 263696
rect 67634 263684 67640 263696
rect 56468 263656 67640 263684
rect 56468 263644 56474 263656
rect 67634 263644 67640 263656
rect 67692 263644 67698 263696
rect 8938 263576 8944 263628
rect 8996 263616 9002 263628
rect 67726 263616 67732 263628
rect 8996 263588 67732 263616
rect 8996 263576 9002 263588
rect 67726 263576 67732 263588
rect 67784 263576 67790 263628
rect 18598 263508 18604 263560
rect 18656 263548 18662 263560
rect 67634 263548 67640 263560
rect 18656 263520 67640 263548
rect 18656 263508 18662 263520
rect 67634 263508 67640 263520
rect 67692 263508 67698 263560
rect 121454 262828 121460 262880
rect 121512 262868 121518 262880
rect 254026 262868 254032 262880
rect 121512 262840 254032 262868
rect 121512 262828 121518 262840
rect 254026 262828 254032 262840
rect 254084 262828 254090 262880
rect 64598 262216 64604 262268
rect 64656 262256 64662 262268
rect 67634 262256 67640 262268
rect 64656 262228 67640 262256
rect 64656 262216 64662 262228
rect 67634 262216 67640 262228
rect 67692 262216 67698 262268
rect 121454 262216 121460 262268
rect 121512 262256 121518 262268
rect 327166 262256 327172 262268
rect 121512 262228 327172 262256
rect 121512 262216 121518 262228
rect 327166 262216 327172 262228
rect 327224 262216 327230 262268
rect 53466 260856 53472 260908
rect 53524 260896 53530 260908
rect 67726 260896 67732 260908
rect 53524 260868 67732 260896
rect 53524 260856 53530 260868
rect 67726 260856 67732 260868
rect 67784 260856 67790 260908
rect 121454 260856 121460 260908
rect 121512 260896 121518 260908
rect 342438 260896 342444 260908
rect 121512 260868 342444 260896
rect 121512 260856 121518 260868
rect 342438 260856 342444 260868
rect 342496 260856 342502 260908
rect 36538 260788 36544 260840
rect 36596 260828 36602 260840
rect 67634 260828 67640 260840
rect 36596 260800 67640 260828
rect 36596 260788 36602 260800
rect 67634 260788 67640 260800
rect 67692 260788 67698 260840
rect 62022 259428 62028 259480
rect 62080 259468 62086 259480
rect 67634 259468 67640 259480
rect 62080 259440 67640 259468
rect 62080 259428 62086 259440
rect 67634 259428 67640 259440
rect 67692 259428 67698 259480
rect 121454 259428 121460 259480
rect 121512 259468 121518 259480
rect 267734 259468 267740 259480
rect 121512 259440 267740 259468
rect 121512 259428 121518 259440
rect 267734 259428 267740 259440
rect 267792 259428 267798 259480
rect 126422 259360 126428 259412
rect 126480 259400 126486 259412
rect 579614 259400 579620 259412
rect 126480 259372 579620 259400
rect 126480 259360 126486 259372
rect 579614 259360 579620 259372
rect 579672 259360 579678 259412
rect 121454 259292 121460 259344
rect 121512 259332 121518 259344
rect 149698 259332 149704 259344
rect 121512 259304 149704 259332
rect 121512 259292 121518 259304
rect 149698 259292 149704 259304
rect 149756 259292 149762 259344
rect 60458 258680 60464 258732
rect 60516 258720 60522 258732
rect 67818 258720 67824 258732
rect 60516 258692 67824 258720
rect 60516 258680 60522 258692
rect 67818 258680 67824 258692
rect 67876 258680 67882 258732
rect 63310 258136 63316 258188
rect 63368 258176 63374 258188
rect 67634 258176 67640 258188
rect 63368 258148 67640 258176
rect 63368 258136 63374 258148
rect 67634 258136 67640 258148
rect 67692 258136 67698 258188
rect 59078 258068 59084 258120
rect 59136 258108 59142 258120
rect 67726 258108 67732 258120
rect 59136 258080 67732 258108
rect 59136 258068 59142 258080
rect 67726 258068 67732 258080
rect 67784 258068 67790 258120
rect 122190 257320 122196 257372
rect 122248 257360 122254 257372
rect 332870 257360 332876 257372
rect 122248 257332 332876 257360
rect 122248 257320 122254 257332
rect 332870 257320 332876 257332
rect 332928 257320 332934 257372
rect 121454 257116 121460 257168
rect 121512 257156 121518 257168
rect 123570 257156 123576 257168
rect 121512 257128 123576 257156
rect 121512 257116 121518 257128
rect 123570 257116 123576 257128
rect 123628 257116 123634 257168
rect 53558 256776 53564 256828
rect 53616 256816 53622 256828
rect 67634 256816 67640 256828
rect 53616 256788 67640 256816
rect 53616 256776 53622 256788
rect 67634 256776 67640 256788
rect 67692 256776 67698 256828
rect 14458 256708 14464 256760
rect 14516 256748 14522 256760
rect 67726 256748 67732 256760
rect 14516 256720 67732 256748
rect 14516 256708 14522 256720
rect 67726 256708 67732 256720
rect 67784 256708 67790 256760
rect 121638 256708 121644 256760
rect 121696 256748 121702 256760
rect 232498 256748 232504 256760
rect 121696 256720 232504 256748
rect 121696 256708 121702 256720
rect 232498 256708 232504 256720
rect 232556 256708 232562 256760
rect 121546 256640 121552 256692
rect 121604 256680 121610 256692
rect 130378 256680 130384 256692
rect 121604 256652 130384 256680
rect 121604 256640 121610 256652
rect 130378 256640 130384 256652
rect 130436 256640 130442 256692
rect 121454 256436 121460 256488
rect 121512 256476 121518 256488
rect 123478 256476 123484 256488
rect 121512 256448 123484 256476
rect 121512 256436 121518 256448
rect 123478 256436 123484 256448
rect 123536 256436 123542 256488
rect 61746 255348 61752 255400
rect 61804 255388 61810 255400
rect 67634 255388 67640 255400
rect 61804 255360 67640 255388
rect 61804 255348 61810 255360
rect 67634 255348 67640 255360
rect 67692 255348 67698 255400
rect 50982 255280 50988 255332
rect 51040 255320 51046 255332
rect 67726 255320 67732 255332
rect 51040 255292 67732 255320
rect 51040 255280 51046 255292
rect 67726 255280 67732 255292
rect 67784 255280 67790 255332
rect 63402 255212 63408 255264
rect 63460 255252 63466 255264
rect 67634 255252 67640 255264
rect 63460 255224 67640 255252
rect 63460 255212 63466 255224
rect 67634 255212 67640 255224
rect 67692 255212 67698 255264
rect 121454 253988 121460 254040
rect 121512 254028 121518 254040
rect 197998 254028 198004 254040
rect 121512 254000 198004 254028
rect 121512 253988 121518 254000
rect 197998 253988 198004 254000
rect 198056 253988 198062 254040
rect 3142 253920 3148 253972
rect 3200 253960 3206 253972
rect 13078 253960 13084 253972
rect 3200 253932 13084 253960
rect 3200 253920 3206 253932
rect 13078 253920 13084 253932
rect 13136 253920 13142 253972
rect 121546 253920 121552 253972
rect 121604 253960 121610 253972
rect 323670 253960 323676 253972
rect 121604 253932 323676 253960
rect 121604 253920 121610 253932
rect 323670 253920 323676 253932
rect 323728 253920 323734 253972
rect 121638 253172 121644 253224
rect 121696 253212 121702 253224
rect 144178 253212 144184 253224
rect 121696 253184 144184 253212
rect 121696 253172 121702 253184
rect 144178 253172 144184 253184
rect 144236 253172 144242 253224
rect 65886 252628 65892 252680
rect 65944 252668 65950 252680
rect 68094 252668 68100 252680
rect 65944 252640 68100 252668
rect 65944 252628 65950 252640
rect 68094 252628 68100 252640
rect 68152 252628 68158 252680
rect 121546 252628 121552 252680
rect 121604 252668 121610 252680
rect 233878 252668 233884 252680
rect 121604 252640 233884 252668
rect 121604 252628 121610 252640
rect 233878 252628 233884 252640
rect 233936 252628 233942 252680
rect 44818 252560 44824 252612
rect 44876 252600 44882 252612
rect 67634 252600 67640 252612
rect 44876 252572 67640 252600
rect 44876 252560 44882 252572
rect 67634 252560 67640 252572
rect 67692 252560 67698 252612
rect 121454 252560 121460 252612
rect 121512 252600 121518 252612
rect 347866 252600 347872 252612
rect 121512 252572 347872 252600
rect 121512 252560 121518 252572
rect 347866 252560 347872 252572
rect 347924 252560 347930 252612
rect 119798 251812 119804 251864
rect 119856 251852 119862 251864
rect 142798 251852 142804 251864
rect 119856 251824 142804 251852
rect 119856 251812 119862 251824
rect 142798 251812 142804 251824
rect 142856 251812 142862 251864
rect 121454 251200 121460 251252
rect 121512 251240 121518 251252
rect 346486 251240 346492 251252
rect 121512 251212 346492 251240
rect 121512 251200 121518 251212
rect 346486 251200 346492 251212
rect 346544 251200 346550 251252
rect 122098 250452 122104 250504
rect 122156 250492 122162 250504
rect 331306 250492 331312 250504
rect 122156 250464 331312 250492
rect 122156 250452 122162 250464
rect 331306 250452 331312 250464
rect 331364 250452 331370 250504
rect 64690 249840 64696 249892
rect 64748 249880 64754 249892
rect 67634 249880 67640 249892
rect 64748 249852 67640 249880
rect 64748 249840 64754 249852
rect 67634 249840 67640 249852
rect 67692 249840 67698 249892
rect 63126 249772 63132 249824
rect 63184 249812 63190 249824
rect 67726 249812 67732 249824
rect 63184 249784 67732 249812
rect 63184 249772 63190 249784
rect 67726 249772 67732 249784
rect 67784 249772 67790 249824
rect 121546 249772 121552 249824
rect 121604 249812 121610 249824
rect 203518 249812 203524 249824
rect 121604 249784 203524 249812
rect 121604 249772 121610 249784
rect 203518 249772 203524 249784
rect 203576 249772 203582 249824
rect 59262 249704 59268 249756
rect 59320 249744 59326 249756
rect 67634 249744 67640 249756
rect 59320 249716 67640 249744
rect 59320 249704 59326 249716
rect 67634 249704 67640 249716
rect 67692 249704 67698 249756
rect 121454 249704 121460 249756
rect 121512 249744 121518 249756
rect 140038 249744 140044 249756
rect 121512 249716 140044 249744
rect 121512 249704 121518 249716
rect 140038 249704 140044 249716
rect 140096 249704 140102 249756
rect 166258 249024 166264 249076
rect 166316 249064 166322 249076
rect 305638 249064 305644 249076
rect 166316 249036 305644 249064
rect 166316 249024 166322 249036
rect 305638 249024 305644 249036
rect 305696 249024 305702 249076
rect 58986 248412 58992 248464
rect 59044 248452 59050 248464
rect 67634 248452 67640 248464
rect 59044 248424 67640 248452
rect 59044 248412 59050 248424
rect 67634 248412 67640 248424
rect 67692 248412 67698 248464
rect 121454 248412 121460 248464
rect 121512 248452 121518 248464
rect 309778 248452 309784 248464
rect 121512 248424 309784 248452
rect 121512 248412 121518 248424
rect 309778 248412 309784 248424
rect 309836 248412 309842 248464
rect 247678 247664 247684 247716
rect 247736 247704 247742 247716
rect 580442 247704 580448 247716
rect 247736 247676 580448 247704
rect 247736 247664 247742 247676
rect 580442 247664 580448 247676
rect 580500 247664 580506 247716
rect 61838 247120 61844 247172
rect 61896 247160 61902 247172
rect 67634 247160 67640 247172
rect 61896 247132 67640 247160
rect 61896 247120 61902 247132
rect 67634 247120 67640 247132
rect 67692 247120 67698 247172
rect 59262 247052 59268 247104
rect 59320 247092 59326 247104
rect 67726 247092 67732 247104
rect 59320 247064 67732 247092
rect 59320 247052 59326 247064
rect 67726 247052 67732 247064
rect 67784 247052 67790 247104
rect 121454 247052 121460 247104
rect 121512 247092 121518 247104
rect 229738 247092 229744 247104
rect 121512 247064 229744 247092
rect 121512 247052 121518 247064
rect 229738 247052 229744 247064
rect 229796 247052 229802 247104
rect 49602 246984 49608 247036
rect 49660 247024 49666 247036
rect 67634 247024 67640 247036
rect 49660 246996 67640 247024
rect 49660 246984 49666 246996
rect 67634 246984 67640 246996
rect 67692 246984 67698 247036
rect 121546 245624 121552 245676
rect 121604 245664 121610 245676
rect 270494 245664 270500 245676
rect 121604 245636 270500 245664
rect 121604 245624 121610 245636
rect 270494 245624 270500 245636
rect 270552 245624 270558 245676
rect 17218 245556 17224 245608
rect 17276 245596 17282 245608
rect 67634 245596 67640 245608
rect 17276 245568 67640 245596
rect 17276 245556 17282 245568
rect 67634 245556 67640 245568
rect 67692 245556 67698 245608
rect 121454 245556 121460 245608
rect 121512 245596 121518 245608
rect 128998 245596 129004 245608
rect 121512 245568 129004 245596
rect 121512 245556 121518 245568
rect 128998 245556 129004 245568
rect 129056 245556 129062 245608
rect 63402 244264 63408 244316
rect 63460 244304 63466 244316
rect 67634 244304 67640 244316
rect 63460 244276 67640 244304
rect 63460 244264 63466 244276
rect 67634 244264 67640 244276
rect 67692 244264 67698 244316
rect 121546 244264 121552 244316
rect 121604 244304 121610 244316
rect 323578 244304 323584 244316
rect 121604 244276 323584 244304
rect 121604 244264 121610 244276
rect 323578 244264 323584 244276
rect 323636 244264 323642 244316
rect 4798 244196 4804 244248
rect 4856 244236 4862 244248
rect 67726 244236 67732 244248
rect 4856 244208 67732 244236
rect 4856 244196 4862 244208
rect 67726 244196 67732 244208
rect 67784 244196 67790 244248
rect 121454 243720 121460 243772
rect 121512 243760 121518 243772
rect 125134 243760 125140 243772
rect 121512 243732 125140 243760
rect 121512 243720 121518 243732
rect 125134 243720 125140 243732
rect 125192 243720 125198 243772
rect 340966 243516 340972 243568
rect 341024 243556 341030 243568
rect 579890 243556 579896 243568
rect 341024 243528 579896 243556
rect 341024 243516 341030 243528
rect 579890 243516 579896 243528
rect 579948 243516 579954 243568
rect 65978 242904 65984 242956
rect 66036 242944 66042 242956
rect 67818 242944 67824 242956
rect 66036 242916 67824 242944
rect 66036 242904 66042 242916
rect 67818 242904 67824 242916
rect 67876 242904 67882 242956
rect 121546 242904 121552 242956
rect 121604 242944 121610 242956
rect 311250 242944 311256 242956
rect 121604 242916 311256 242944
rect 121604 242904 121610 242916
rect 311250 242904 311256 242916
rect 311308 242904 311314 242956
rect 53742 242836 53748 242888
rect 53800 242876 53806 242888
rect 67634 242876 67640 242888
rect 53800 242848 67640 242876
rect 53800 242836 53806 242848
rect 67634 242836 67640 242848
rect 67692 242836 67698 242888
rect 121454 242836 121460 242888
rect 121512 242876 121518 242888
rect 340966 242876 340972 242888
rect 121512 242848 340972 242876
rect 121512 242836 121518 242848
rect 340966 242836 340972 242848
rect 341024 242836 341030 242888
rect 121546 242768 121552 242820
rect 121604 242808 121610 242820
rect 134518 242808 134524 242820
rect 121604 242780 134524 242808
rect 121604 242768 121610 242780
rect 134518 242768 134524 242780
rect 134576 242768 134582 242820
rect 63218 241476 63224 241528
rect 63276 241516 63282 241528
rect 67726 241516 67732 241528
rect 63276 241488 67732 241516
rect 63276 241476 63282 241488
rect 67726 241476 67732 241488
rect 67784 241476 67790 241528
rect 59170 241408 59176 241460
rect 59228 241448 59234 241460
rect 67634 241448 67640 241460
rect 59228 241420 67640 241448
rect 59228 241408 59234 241420
rect 67634 241408 67640 241420
rect 67692 241408 67698 241460
rect 119798 240184 119804 240236
rect 119856 240184 119862 240236
rect 121546 240184 121552 240236
rect 121604 240224 121610 240236
rect 328546 240224 328552 240236
rect 121604 240196 328552 240224
rect 121604 240184 121610 240196
rect 328546 240184 328552 240196
rect 328604 240184 328610 240236
rect 3050 240116 3056 240168
rect 3108 240156 3114 240168
rect 16574 240156 16580 240168
rect 3108 240128 16580 240156
rect 3108 240116 3114 240128
rect 16574 240116 16580 240128
rect 16632 240116 16638 240168
rect 65886 239912 65892 239964
rect 65944 239952 65950 239964
rect 71038 239952 71044 239964
rect 65944 239924 71044 239952
rect 65944 239912 65950 239924
rect 71038 239912 71044 239924
rect 71096 239912 71102 239964
rect 118970 239912 118976 239964
rect 119028 239952 119034 239964
rect 119816 239952 119844 240184
rect 119890 240116 119896 240168
rect 119948 240156 119954 240168
rect 330110 240156 330116 240168
rect 119948 240128 330116 240156
rect 119948 240116 119954 240128
rect 330110 240116 330116 240128
rect 330168 240116 330174 240168
rect 119028 239924 119844 239952
rect 119028 239912 119034 239924
rect 70578 239368 70584 239420
rect 70636 239408 70642 239420
rect 86218 239408 86224 239420
rect 70636 239380 86224 239408
rect 70636 239368 70642 239380
rect 86218 239368 86224 239380
rect 86276 239368 86282 239420
rect 117038 238824 117044 238876
rect 117096 238864 117102 238876
rect 126238 238864 126244 238876
rect 117096 238836 126244 238864
rect 117096 238824 117102 238836
rect 126238 238824 126244 238836
rect 126296 238824 126302 238876
rect 40034 238756 40040 238808
rect 40092 238796 40098 238808
rect 95786 238796 95792 238808
rect 40092 238768 95792 238796
rect 40092 238756 40098 238768
rect 95786 238756 95792 238768
rect 95844 238756 95850 238808
rect 115106 238756 115112 238808
rect 115164 238796 115170 238808
rect 582466 238796 582472 238808
rect 115164 238768 582472 238796
rect 115164 238756 115170 238768
rect 582466 238756 582472 238768
rect 582524 238756 582530 238808
rect 3510 238688 3516 238740
rect 3568 238728 3574 238740
rect 86770 238728 86776 238740
rect 3568 238700 86776 238728
rect 3568 238688 3574 238700
rect 86770 238688 86776 238700
rect 86828 238688 86834 238740
rect 113818 238688 113824 238740
rect 113876 238728 113882 238740
rect 494054 238728 494060 238740
rect 113876 238700 494060 238728
rect 113876 238688 113882 238700
rect 494054 238688 494060 238700
rect 494112 238688 494118 238740
rect 72602 238620 72608 238672
rect 72660 238660 72666 238672
rect 130470 238660 130476 238672
rect 72660 238632 130476 238660
rect 72660 238620 72666 238632
rect 130470 238620 130476 238632
rect 130528 238620 130534 238672
rect 50338 238552 50344 238604
rect 50396 238592 50402 238604
rect 99006 238592 99012 238604
rect 50396 238564 99012 238592
rect 50396 238552 50402 238564
rect 99006 238552 99012 238564
rect 99064 238552 99070 238604
rect 135898 238592 135904 238604
rect 103486 238564 135904 238592
rect 55122 238484 55128 238536
rect 55180 238524 55186 238536
rect 89346 238524 89352 238536
rect 55180 238496 89352 238524
rect 55180 238484 55186 238496
rect 89346 238484 89352 238496
rect 89404 238484 89410 238536
rect 98362 238484 98368 238536
rect 98420 238524 98426 238536
rect 103486 238524 103514 238564
rect 135898 238552 135904 238564
rect 135956 238552 135962 238604
rect 98420 238496 103514 238524
rect 98420 238484 98426 238496
rect 95142 238144 95148 238196
rect 95200 238184 95206 238196
rect 106918 238184 106924 238196
rect 95200 238156 106924 238184
rect 95200 238144 95206 238156
rect 106918 238144 106924 238156
rect 106976 238144 106982 238196
rect 105446 238076 105452 238128
rect 105504 238116 105510 238128
rect 188338 238116 188344 238128
rect 105504 238088 188344 238116
rect 105504 238076 105510 238088
rect 188338 238076 188344 238088
rect 188396 238076 188402 238128
rect 74534 238008 74540 238060
rect 74592 238048 74598 238060
rect 338114 238048 338120 238060
rect 74592 238020 338120 238048
rect 74592 238008 74598 238020
rect 338114 238008 338120 238020
rect 338172 238008 338178 238060
rect 79042 237600 79048 237652
rect 79100 237640 79106 237652
rect 80698 237640 80704 237652
rect 79100 237612 80704 237640
rect 79100 237600 79106 237612
rect 80698 237600 80704 237612
rect 80756 237600 80762 237652
rect 71314 237396 71320 237448
rect 71372 237436 71378 237448
rect 75178 237436 75184 237448
rect 71372 237408 75184 237436
rect 71372 237396 71378 237408
rect 75178 237396 75184 237408
rect 75236 237396 75242 237448
rect 43438 237328 43444 237380
rect 43496 237368 43502 237380
rect 82262 237368 82268 237380
rect 43496 237340 82268 237368
rect 43496 237328 43502 237340
rect 82262 237328 82268 237340
rect 82320 237328 82326 237380
rect 91922 237328 91928 237380
rect 91980 237368 91986 237380
rect 582742 237368 582748 237380
rect 91980 237340 582748 237368
rect 91980 237328 91986 237340
rect 582742 237328 582748 237340
rect 582800 237328 582806 237380
rect 16574 237260 16580 237312
rect 16632 237300 16638 237312
rect 103514 237300 103520 237312
rect 16632 237272 103520 237300
rect 16632 237260 16638 237272
rect 103514 237260 103520 237272
rect 103572 237260 103578 237312
rect 31018 237192 31024 237244
rect 31076 237232 31082 237244
rect 114462 237232 114468 237244
rect 31076 237204 114468 237232
rect 31076 237192 31082 237204
rect 114462 237192 114468 237204
rect 114520 237192 114526 237244
rect 97718 236648 97724 236700
rect 97776 236688 97782 236700
rect 340966 236688 340972 236700
rect 97776 236660 340972 236688
rect 97776 236648 97782 236660
rect 340966 236648 340972 236660
rect 341024 236648 341030 236700
rect 106734 235900 106740 235952
rect 106792 235940 106798 235952
rect 264238 235940 264244 235952
rect 106792 235912 264244 235940
rect 106792 235900 106798 235912
rect 264238 235900 264244 235912
rect 264296 235900 264302 235952
rect 13078 235832 13084 235884
rect 13136 235872 13142 235884
rect 112530 235872 112536 235884
rect 13136 235844 112536 235872
rect 13136 235832 13142 235844
rect 112530 235832 112536 235844
rect 112588 235832 112594 235884
rect 63402 235356 63408 235408
rect 63460 235396 63466 235408
rect 280154 235396 280160 235408
rect 63460 235368 280160 235396
rect 63460 235356 63466 235368
rect 280154 235356 280160 235368
rect 280212 235356 280218 235408
rect 108022 235288 108028 235340
rect 108080 235328 108086 235340
rect 327350 235328 327356 235340
rect 108080 235300 327356 235328
rect 108080 235288 108086 235300
rect 327350 235288 327356 235300
rect 327408 235288 327414 235340
rect 64782 235220 64788 235272
rect 64840 235260 64846 235272
rect 121454 235260 121460 235272
rect 64840 235232 121460 235260
rect 64840 235220 64846 235232
rect 121454 235220 121460 235232
rect 121512 235220 121518 235272
rect 60458 233928 60464 233980
rect 60516 233968 60522 233980
rect 192570 233968 192576 233980
rect 60516 233940 192576 233968
rect 60516 233928 60522 233940
rect 192570 233928 192576 233940
rect 192628 233928 192634 233980
rect 84286 233860 84292 233912
rect 84344 233900 84350 233912
rect 85482 233900 85488 233912
rect 84344 233872 85488 233900
rect 84344 233860 84350 233872
rect 85482 233860 85488 233872
rect 85540 233860 85546 233912
rect 95234 233860 95240 233912
rect 95292 233900 95298 233912
rect 96430 233900 96436 233912
rect 95292 233872 96436 233900
rect 95292 233860 95298 233872
rect 96430 233860 96436 233872
rect 96488 233860 96494 233912
rect 99374 233860 99380 233912
rect 99432 233900 99438 233912
rect 100294 233900 100300 233912
rect 99432 233872 100300 233900
rect 99432 233860 99438 233872
rect 100294 233860 100300 233872
rect 100352 233860 100358 233912
rect 103606 233860 103612 233912
rect 103664 233900 103670 233912
rect 104802 233900 104808 233912
rect 103664 233872 104808 233900
rect 103664 233860 103670 233872
rect 104802 233860 104808 233872
rect 104860 233860 104866 233912
rect 104894 233860 104900 233912
rect 104952 233900 104958 233912
rect 106090 233900 106096 233912
rect 104952 233872 106096 233900
rect 104952 233860 104958 233872
rect 106090 233860 106096 233872
rect 106148 233860 106154 233912
rect 110414 233860 110420 233912
rect 110472 233900 110478 233912
rect 111242 233900 111248 233912
rect 110472 233872 111248 233900
rect 110472 233860 110478 233872
rect 111242 233860 111248 233872
rect 111300 233860 111306 233912
rect 117682 233860 117688 233912
rect 117740 233900 117746 233912
rect 582466 233900 582472 233912
rect 117740 233872 582472 233900
rect 117740 233860 117746 233872
rect 582466 233860 582472 233872
rect 582524 233860 582530 233912
rect 75822 233180 75828 233232
rect 75880 233220 75886 233232
rect 582374 233220 582380 233232
rect 75880 233192 582380 233220
rect 75880 233180 75886 233192
rect 582374 233180 582380 233192
rect 582432 233180 582438 233232
rect 73154 232976 73160 233028
rect 73212 233016 73218 233028
rect 73890 233016 73896 233028
rect 73212 232988 73896 233016
rect 73212 232976 73218 232988
rect 73890 232976 73896 232988
rect 73948 232976 73954 233028
rect 67358 232500 67364 232552
rect 67416 232540 67422 232552
rect 324406 232540 324412 232552
rect 67416 232512 324412 232540
rect 67416 232500 67422 232512
rect 324406 232500 324412 232512
rect 324464 232500 324470 232552
rect 114554 232160 114560 232212
rect 114612 232200 114618 232212
rect 115750 232200 115756 232212
rect 114612 232172 115756 232200
rect 114612 232160 114618 232172
rect 115750 232160 115756 232172
rect 115808 232160 115814 232212
rect 84102 231820 84108 231872
rect 84160 231860 84166 231872
rect 84838 231860 84844 231872
rect 84160 231832 84844 231860
rect 84160 231820 84166 231832
rect 84838 231820 84844 231832
rect 84896 231820 84902 231872
rect 81618 231752 81624 231804
rect 81676 231792 81682 231804
rect 214558 231792 214564 231804
rect 81676 231764 214564 231792
rect 81676 231752 81682 231764
rect 214558 231752 214564 231764
rect 214616 231752 214622 231804
rect 93210 231072 93216 231124
rect 93268 231112 93274 231124
rect 331398 231112 331404 231124
rect 93268 231084 331404 231112
rect 93268 231072 93274 231084
rect 331398 231072 331404 231084
rect 331456 231072 331462 231124
rect 100754 231004 100760 231056
rect 100812 231044 100818 231056
rect 101582 231044 101588 231056
rect 100812 231016 101588 231044
rect 100812 231004 100818 231016
rect 101582 231004 101588 231016
rect 101640 231004 101646 231056
rect 82906 229848 82912 229900
rect 82964 229888 82970 229900
rect 175918 229888 175924 229900
rect 82964 229860 175924 229888
rect 82964 229848 82970 229860
rect 175918 229848 175924 229860
rect 175976 229848 175982 229900
rect 88058 229780 88064 229832
rect 88116 229820 88122 229832
rect 252554 229820 252560 229832
rect 88116 229792 252560 229820
rect 88116 229780 88122 229792
rect 252554 229780 252560 229792
rect 252612 229780 252618 229832
rect 80054 229712 80060 229764
rect 80112 229752 80118 229764
rect 80974 229752 80980 229764
rect 80112 229724 80980 229752
rect 80112 229712 80118 229724
rect 80974 229712 80980 229724
rect 81032 229712 81038 229764
rect 86126 229712 86132 229764
rect 86184 229752 86190 229764
rect 582374 229752 582380 229764
rect 86184 229724 582380 229752
rect 86184 229712 86190 229724
rect 582374 229712 582380 229724
rect 582432 229712 582438 229764
rect 106826 229032 106832 229084
rect 106884 229072 106890 229084
rect 542354 229072 542360 229084
rect 106884 229044 542360 229072
rect 106884 229032 106890 229044
rect 542354 229032 542360 229044
rect 542412 229032 542418 229084
rect 69106 228352 69112 228404
rect 69164 228392 69170 228404
rect 321646 228392 321652 228404
rect 69164 228364 321652 228392
rect 69164 228352 69170 228364
rect 321646 228352 321652 228364
rect 321704 228352 321710 228404
rect 61746 227060 61752 227112
rect 61804 227100 61810 227112
rect 276014 227100 276020 227112
rect 61804 227072 276020 227100
rect 61804 227060 61810 227072
rect 276014 227060 276020 227072
rect 276072 227060 276078 227112
rect 99650 226992 99656 227044
rect 99708 227032 99714 227044
rect 343726 227032 343732 227044
rect 99708 227004 343732 227032
rect 99708 226992 99714 227004
rect 343726 226992 343732 227004
rect 343784 226992 343790 227044
rect 80330 225632 80336 225684
rect 80388 225672 80394 225684
rect 315298 225672 315304 225684
rect 80388 225644 315304 225672
rect 80388 225632 80394 225644
rect 315298 225632 315304 225644
rect 315356 225632 315362 225684
rect 50890 225564 50896 225616
rect 50948 225604 50954 225616
rect 309870 225604 309876 225616
rect 50948 225576 309876 225604
rect 50948 225564 50954 225576
rect 309870 225564 309876 225576
rect 309928 225564 309934 225616
rect 64506 224204 64512 224256
rect 64564 224244 64570 224256
rect 214558 224244 214564 224256
rect 64564 224216 214564 224244
rect 64564 224204 64570 224216
rect 214558 224204 214564 224216
rect 214616 224204 214622 224256
rect 13078 223048 13084 223100
rect 13136 223088 13142 223100
rect 110598 223088 110604 223100
rect 13136 223060 110604 223088
rect 13136 223048 13142 223060
rect 110598 223048 110604 223060
rect 110656 223048 110662 223100
rect 94498 222980 94504 223032
rect 94556 223020 94562 223032
rect 287698 223020 287704 223032
rect 94556 222992 287704 223020
rect 94556 222980 94562 222992
rect 287698 222980 287704 222992
rect 287756 222980 287762 223032
rect 108666 222912 108672 222964
rect 108724 222952 108730 222964
rect 329926 222952 329932 222964
rect 108724 222924 329932 222952
rect 108724 222912 108730 222924
rect 329926 222912 329932 222924
rect 329984 222912 329990 222964
rect 45462 222844 45468 222896
rect 45520 222884 45526 222896
rect 312538 222884 312544 222896
rect 45520 222856 312544 222884
rect 45520 222844 45526 222856
rect 312538 222844 312544 222856
rect 312596 222844 312602 222896
rect 4798 221416 4804 221468
rect 4856 221456 4862 221468
rect 83550 221456 83556 221468
rect 4856 221428 83556 221456
rect 4856 221416 4862 221428
rect 83550 221416 83556 221428
rect 83608 221416 83614 221468
rect 102870 221416 102876 221468
rect 102928 221456 102934 221468
rect 252646 221456 252652 221468
rect 102928 221428 252652 221456
rect 102928 221416 102934 221428
rect 252646 221416 252652 221428
rect 252704 221416 252710 221468
rect 74902 220192 74908 220244
rect 74960 220232 74966 220244
rect 254118 220232 254124 220244
rect 74960 220204 254124 220232
rect 74960 220192 74966 220204
rect 254118 220192 254124 220204
rect 254176 220192 254182 220244
rect 80698 220124 80704 220176
rect 80756 220164 80762 220176
rect 263686 220164 263692 220176
rect 80756 220136 263692 220164
rect 80756 220124 80762 220136
rect 263686 220124 263692 220136
rect 263744 220124 263750 220176
rect 71038 220056 71044 220108
rect 71096 220096 71102 220108
rect 334250 220096 334256 220108
rect 71096 220068 334256 220096
rect 71096 220056 71102 220068
rect 334250 220056 334256 220068
rect 334308 220056 334314 220108
rect 63218 218764 63224 218816
rect 63276 218804 63282 218816
rect 228358 218804 228364 218816
rect 63276 218776 228364 218804
rect 63276 218764 63282 218776
rect 228358 218764 228364 218776
rect 228416 218764 228422 218816
rect 48222 218696 48228 218748
rect 48280 218736 48286 218748
rect 346578 218736 346584 218748
rect 48280 218708 346584 218736
rect 48280 218696 48286 218708
rect 346578 218696 346584 218708
rect 346636 218696 346642 218748
rect 61930 217404 61936 217456
rect 61988 217444 61994 217456
rect 262214 217444 262220 217456
rect 61988 217416 262220 217444
rect 61988 217404 61994 217416
rect 262214 217404 262220 217416
rect 262272 217404 262278 217456
rect 58986 217336 58992 217388
rect 59044 217376 59050 217388
rect 277394 217376 277400 217388
rect 59044 217348 277400 217376
rect 59044 217336 59050 217348
rect 277394 217336 277400 217348
rect 277452 217336 277458 217388
rect 53466 217268 53472 217320
rect 53524 217308 53530 217320
rect 318242 217308 318248 217320
rect 53524 217280 318248 217308
rect 53524 217268 53530 217280
rect 318242 217268 318248 217280
rect 318300 217268 318306 217320
rect 86218 215976 86224 216028
rect 86276 216016 86282 216028
rect 314010 216016 314016 216028
rect 86276 215988 314016 216016
rect 86276 215976 86282 215988
rect 314010 215976 314016 215988
rect 314068 215976 314074 216028
rect 56410 215908 56416 215960
rect 56468 215948 56474 215960
rect 291838 215948 291844 215960
rect 56468 215920 291844 215948
rect 56468 215908 56474 215920
rect 291838 215908 291844 215920
rect 291896 215908 291902 215960
rect 3510 214956 3516 215008
rect 3568 214996 3574 215008
rect 8938 214996 8944 215008
rect 3568 214968 8944 214996
rect 3568 214956 3574 214968
rect 8938 214956 8944 214968
rect 8996 214956 9002 215008
rect 66070 214616 66076 214668
rect 66128 214656 66134 214668
rect 251174 214656 251180 214668
rect 66128 214628 251180 214656
rect 66128 214616 66134 214628
rect 251174 214616 251180 214628
rect 251232 214616 251238 214668
rect 78674 214548 78680 214600
rect 78732 214588 78738 214600
rect 330018 214588 330024 214600
rect 78732 214560 330024 214588
rect 78732 214548 78738 214560
rect 330018 214548 330024 214560
rect 330076 214548 330082 214600
rect 63310 213324 63316 213376
rect 63368 213364 63374 213376
rect 224310 213364 224316 213376
rect 63368 213336 224316 213364
rect 63368 213324 63374 213336
rect 224310 213324 224316 213336
rect 224368 213324 224374 213376
rect 93854 213256 93860 213308
rect 93912 213296 93918 213308
rect 278866 213296 278872 213308
rect 93912 213268 278872 213296
rect 93912 213256 93918 213268
rect 278866 213256 278872 213268
rect 278924 213256 278930 213308
rect 106918 213188 106924 213240
rect 106976 213228 106982 213240
rect 341058 213228 341064 213240
rect 106976 213200 341064 213228
rect 106976 213188 106982 213200
rect 341058 213188 341064 213200
rect 341116 213188 341122 213240
rect 67542 211828 67548 211880
rect 67600 211868 67606 211880
rect 251266 211868 251272 211880
rect 67600 211840 251272 211868
rect 67600 211828 67606 211840
rect 251266 211828 251272 211840
rect 251324 211828 251330 211880
rect 57698 211760 57704 211812
rect 57756 211800 57762 211812
rect 271874 211800 271880 211812
rect 57756 211772 271880 211800
rect 57756 211760 57762 211772
rect 271874 211760 271880 211772
rect 271932 211760 271938 211812
rect 192570 210468 192576 210520
rect 192628 210508 192634 210520
rect 307110 210508 307116 210520
rect 192628 210480 307116 210508
rect 192628 210468 192634 210480
rect 307110 210468 307116 210480
rect 307168 210468 307174 210520
rect 84286 210400 84292 210452
rect 84344 210440 84350 210452
rect 249886 210440 249892 210452
rect 84344 210412 249892 210440
rect 84344 210400 84350 210412
rect 249886 210400 249892 210412
rect 249944 210400 249950 210452
rect 160738 209108 160744 209160
rect 160796 209148 160802 209160
rect 300118 209148 300124 209160
rect 160796 209120 300124 209148
rect 160796 209108 160802 209120
rect 300118 209108 300124 209120
rect 300176 209108 300182 209160
rect 67450 209040 67456 209092
rect 67508 209080 67514 209092
rect 324590 209080 324596 209092
rect 67508 209052 324596 209080
rect 67508 209040 67514 209052
rect 324590 209040 324596 209052
rect 324648 209040 324654 209092
rect 125042 206932 125048 206984
rect 125100 206972 125106 206984
rect 580166 206972 580172 206984
rect 125100 206944 580172 206972
rect 125100 206932 125106 206944
rect 580166 206932 580172 206944
rect 580224 206932 580230 206984
rect 56502 206252 56508 206304
rect 56560 206292 56566 206304
rect 266446 206292 266452 206304
rect 56560 206264 266452 206292
rect 56560 206252 56566 206264
rect 266446 206252 266452 206264
rect 266504 206252 266510 206304
rect 92474 204960 92480 205012
rect 92532 205000 92538 205012
rect 252738 205000 252744 205012
rect 92532 204972 252744 205000
rect 92532 204960 92538 204972
rect 252738 204960 252744 204972
rect 252796 204960 252802 205012
rect 63126 204892 63132 204944
rect 63184 204932 63190 204944
rect 242250 204932 242256 204944
rect 63184 204904 242256 204932
rect 63184 204892 63190 204904
rect 242250 204892 242256 204904
rect 242308 204892 242314 204944
rect 100846 203668 100852 203720
rect 100904 203708 100910 203720
rect 270586 203708 270592 203720
rect 100904 203680 270592 203708
rect 100904 203668 100910 203680
rect 270586 203668 270592 203680
rect 270644 203668 270650 203720
rect 100754 203600 100760 203652
rect 100812 203640 100818 203652
rect 274726 203640 274732 203652
rect 100812 203612 274732 203640
rect 100812 203600 100818 203612
rect 274726 203600 274732 203612
rect 274784 203600 274790 203652
rect 114554 203532 114560 203584
rect 114612 203572 114618 203584
rect 327258 203572 327264 203584
rect 114612 203544 327264 203572
rect 114612 203532 114618 203544
rect 327258 203532 327264 203544
rect 327316 203532 327322 203584
rect 3050 202784 3056 202836
rect 3108 202824 3114 202836
rect 120166 202824 120172 202836
rect 3108 202796 120172 202824
rect 3108 202784 3114 202796
rect 120166 202784 120172 202796
rect 120224 202784 120230 202836
rect 115934 202240 115940 202292
rect 115992 202280 115998 202292
rect 266354 202280 266360 202292
rect 115992 202252 266360 202280
rect 115992 202240 115998 202252
rect 266354 202240 266360 202252
rect 266412 202240 266418 202292
rect 60550 202172 60556 202224
rect 60608 202212 60614 202224
rect 271966 202212 271972 202224
rect 60608 202184 271972 202212
rect 60608 202172 60614 202184
rect 271966 202172 271972 202184
rect 272024 202172 272030 202224
rect 104894 202104 104900 202156
rect 104952 202144 104958 202156
rect 339586 202144 339592 202156
rect 104952 202116 339592 202144
rect 104952 202104 104958 202116
rect 339586 202104 339592 202116
rect 339644 202104 339650 202156
rect 89806 200880 89812 200932
rect 89864 200920 89870 200932
rect 254210 200920 254216 200932
rect 89864 200892 254216 200920
rect 89864 200880 89870 200892
rect 254210 200880 254216 200892
rect 254268 200880 254274 200932
rect 64598 200812 64604 200864
rect 64656 200852 64662 200864
rect 260834 200852 260840 200864
rect 64656 200824 260840 200852
rect 64656 200812 64662 200824
rect 260834 200812 260840 200824
rect 260892 200812 260898 200864
rect 103698 200744 103704 200796
rect 103756 200784 103762 200796
rect 321554 200784 321560 200796
rect 103756 200756 321560 200784
rect 103756 200744 103762 200756
rect 321554 200744 321560 200756
rect 321612 200744 321618 200796
rect 86954 199588 86960 199640
rect 87012 199628 87018 199640
rect 196710 199628 196716 199640
rect 87012 199600 196716 199628
rect 87012 199588 87018 199600
rect 196710 199588 196716 199600
rect 196768 199588 196774 199640
rect 99374 199520 99380 199572
rect 99432 199560 99438 199572
rect 249978 199560 249984 199572
rect 99432 199532 249984 199560
rect 99432 199520 99438 199532
rect 249978 199520 249984 199532
rect 250036 199520 250042 199572
rect 148318 199452 148324 199504
rect 148376 199492 148382 199504
rect 334158 199492 334164 199504
rect 148376 199464 334164 199492
rect 148376 199452 148382 199464
rect 334158 199452 334164 199464
rect 334216 199452 334222 199504
rect 59262 199384 59268 199436
rect 59320 199424 59326 199436
rect 258166 199424 258172 199436
rect 59320 199396 258172 199424
rect 59320 199384 59326 199396
rect 258166 199384 258172 199396
rect 258224 199384 258230 199436
rect 96614 198024 96620 198076
rect 96672 198064 96678 198076
rect 259546 198064 259552 198076
rect 96672 198036 259552 198064
rect 96672 198024 96678 198036
rect 259546 198024 259552 198036
rect 259604 198024 259610 198076
rect 59078 197956 59084 198008
rect 59136 197996 59142 198008
rect 273346 197996 273352 198008
rect 59136 197968 273352 197996
rect 59136 197956 59142 197968
rect 273346 197956 273352 197968
rect 273404 197956 273410 198008
rect 111794 196664 111800 196716
rect 111852 196704 111858 196716
rect 262306 196704 262312 196716
rect 111852 196676 262312 196704
rect 111852 196664 111858 196676
rect 262306 196664 262312 196676
rect 262364 196664 262370 196716
rect 77386 196596 77392 196648
rect 77444 196636 77450 196648
rect 264974 196636 264980 196648
rect 77444 196608 264980 196636
rect 77444 196596 77450 196608
rect 264974 196596 264980 196608
rect 265032 196596 265038 196648
rect 53650 195372 53656 195424
rect 53708 195412 53714 195424
rect 240778 195412 240784 195424
rect 53708 195384 240784 195412
rect 53708 195372 53714 195384
rect 240778 195372 240784 195384
rect 240836 195372 240842 195424
rect 69014 195304 69020 195356
rect 69072 195344 69078 195356
rect 324498 195344 324504 195356
rect 69072 195316 324504 195344
rect 69072 195304 69078 195316
rect 324498 195304 324504 195316
rect 324556 195304 324562 195356
rect 53558 195236 53564 195288
rect 53616 195276 53622 195288
rect 336826 195276 336832 195288
rect 53616 195248 336832 195276
rect 53616 195236 53622 195248
rect 336826 195236 336832 195248
rect 336884 195236 336890 195288
rect 75178 193808 75184 193860
rect 75236 193848 75242 193860
rect 269206 193848 269212 193860
rect 75236 193820 269212 193848
rect 75236 193808 75242 193820
rect 269206 193808 269212 193820
rect 269264 193808 269270 193860
rect 89714 192516 89720 192568
rect 89772 192556 89778 192568
rect 252830 192556 252836 192568
rect 89772 192528 252836 192556
rect 89772 192516 89778 192528
rect 252830 192516 252836 192528
rect 252888 192516 252894 192568
rect 84194 192448 84200 192500
rect 84252 192488 84258 192500
rect 337010 192488 337016 192500
rect 84252 192460 337016 192488
rect 84252 192448 84258 192460
rect 337010 192448 337016 192460
rect 337068 192448 337074 192500
rect 224218 191224 224224 191276
rect 224276 191264 224282 191276
rect 256694 191264 256700 191276
rect 224276 191236 256700 191264
rect 224276 191224 224282 191236
rect 256694 191224 256700 191236
rect 256752 191224 256758 191276
rect 122098 191156 122104 191208
rect 122156 191196 122162 191208
rect 250070 191196 250076 191208
rect 122156 191168 250076 191196
rect 122156 191156 122162 191168
rect 250070 191156 250076 191168
rect 250128 191156 250134 191208
rect 75914 191088 75920 191140
rect 75972 191128 75978 191140
rect 582742 191128 582748 191140
rect 75972 191100 582748 191128
rect 75972 191088 75978 191100
rect 582742 191088 582748 191100
rect 582800 191088 582806 191140
rect 43438 189728 43444 189780
rect 43496 189768 43502 189780
rect 109034 189768 109040 189780
rect 43496 189740 109040 189768
rect 43496 189728 43502 189740
rect 109034 189728 109040 189740
rect 109092 189728 109098 189780
rect 157978 189728 157984 189780
rect 158036 189768 158042 189780
rect 339770 189768 339776 189780
rect 158036 189740 339776 189768
rect 158036 189728 158042 189740
rect 339770 189728 339776 189740
rect 339828 189728 339834 189780
rect 106182 189048 106188 189100
rect 106240 189088 106246 189100
rect 211890 189088 211896 189100
rect 106240 189060 211896 189088
rect 106240 189048 106246 189060
rect 211890 189048 211896 189060
rect 211948 189048 211954 189100
rect 207658 188436 207664 188488
rect 207716 188476 207722 188488
rect 269298 188476 269304 188488
rect 207716 188448 269304 188476
rect 207716 188436 207722 188448
rect 269298 188436 269304 188448
rect 269356 188436 269362 188488
rect 192478 188368 192484 188420
rect 192536 188408 192542 188420
rect 267918 188408 267924 188420
rect 192536 188380 267924 188408
rect 192536 188368 192542 188380
rect 267918 188368 267924 188380
rect 267976 188368 267982 188420
rect 88426 188300 88432 188352
rect 88484 188340 88490 188352
rect 328638 188340 328644 188352
rect 88484 188312 328644 188340
rect 88484 188300 88490 188312
rect 328638 188300 328644 188312
rect 328696 188300 328702 188352
rect 100662 187756 100668 187808
rect 100720 187796 100726 187808
rect 171778 187796 171784 187808
rect 100720 187768 171784 187796
rect 100720 187756 100726 187768
rect 171778 187756 171784 187768
rect 171836 187756 171842 187808
rect 107562 187688 107568 187740
rect 107620 187728 107626 187740
rect 207750 187728 207756 187740
rect 107620 187700 207756 187728
rect 107620 187688 107626 187700
rect 207750 187688 207756 187700
rect 207808 187688 207814 187740
rect 197998 187008 198004 187060
rect 198056 187048 198062 187060
rect 256786 187048 256792 187060
rect 198056 187020 256792 187048
rect 198056 187008 198062 187020
rect 256786 187008 256792 187020
rect 256844 187008 256850 187060
rect 50982 186940 50988 186992
rect 51040 186980 51046 186992
rect 338206 186980 338212 186992
rect 51040 186952 338212 186980
rect 51040 186940 51046 186952
rect 338206 186940 338212 186952
rect 338264 186940 338270 186992
rect 126790 186396 126796 186448
rect 126848 186436 126854 186448
rect 171962 186436 171968 186448
rect 126848 186408 171968 186436
rect 126848 186396 126854 186408
rect 171962 186396 171968 186408
rect 172020 186396 172026 186448
rect 117222 186328 117228 186380
rect 117280 186368 117286 186380
rect 214650 186368 214656 186380
rect 117280 186340 214656 186368
rect 117280 186328 117286 186340
rect 214650 186328 214656 186340
rect 214708 186328 214714 186380
rect 185578 185716 185584 185768
rect 185636 185756 185642 185768
rect 255498 185756 255504 185768
rect 185636 185728 255504 185756
rect 185636 185716 185642 185728
rect 255498 185716 255504 185728
rect 255556 185716 255562 185768
rect 95234 185648 95240 185700
rect 95292 185688 95298 185700
rect 321830 185688 321836 185700
rect 95292 185660 321836 185688
rect 95292 185648 95298 185660
rect 321830 185648 321836 185660
rect 321888 185648 321894 185700
rect 80054 185580 80060 185632
rect 80112 185620 80118 185632
rect 322934 185620 322940 185632
rect 80112 185592 322940 185620
rect 80112 185580 80118 185592
rect 322934 185580 322940 185592
rect 322992 185580 322998 185632
rect 118602 184900 118608 184952
rect 118660 184940 118666 184952
rect 170582 184940 170588 184952
rect 118660 184912 170588 184940
rect 118660 184900 118666 184912
rect 170582 184900 170588 184912
rect 170640 184900 170646 184952
rect 102134 184152 102140 184204
rect 102192 184192 102198 184204
rect 321278 184192 321284 184204
rect 102192 184164 321284 184192
rect 102192 184152 102198 184164
rect 321278 184152 321284 184164
rect 321336 184152 321342 184204
rect 124122 183540 124128 183592
rect 124180 183580 124186 183592
rect 167822 183580 167828 183592
rect 124180 183552 167828 183580
rect 124180 183540 124186 183552
rect 167822 183540 167828 183552
rect 167880 183540 167886 183592
rect 233878 183132 233884 183184
rect 233936 183172 233942 183184
rect 260926 183172 260932 183184
rect 233936 183144 260932 183172
rect 233936 183132 233942 183144
rect 260926 183132 260932 183144
rect 260984 183132 260990 183184
rect 211798 183064 211804 183116
rect 211856 183104 211862 183116
rect 261110 183104 261116 183116
rect 211856 183076 261116 183104
rect 211856 183064 211862 183076
rect 261110 183064 261116 183076
rect 261168 183064 261174 183116
rect 166258 182996 166264 183048
rect 166316 183036 166322 183048
rect 332778 183036 332784 183048
rect 166316 183008 332784 183036
rect 166316 182996 166322 183008
rect 332778 182996 332784 183008
rect 332836 182996 332842 183048
rect 73154 182928 73160 182980
rect 73212 182968 73218 182980
rect 321922 182968 321928 182980
rect 73212 182940 321928 182968
rect 73212 182928 73218 182940
rect 321922 182928 321928 182940
rect 321980 182928 321986 182980
rect 65978 182860 65984 182912
rect 66036 182900 66042 182912
rect 338390 182900 338396 182912
rect 66036 182872 338396 182900
rect 66036 182860 66042 182872
rect 338390 182860 338396 182872
rect 338448 182860 338454 182912
rect 62022 182792 62028 182844
rect 62080 182832 62086 182844
rect 345198 182832 345204 182844
rect 62080 182804 345204 182832
rect 62080 182792 62086 182804
rect 345198 182792 345204 182804
rect 345256 182792 345262 182844
rect 128170 182248 128176 182300
rect 128228 182288 128234 182300
rect 166442 182288 166448 182300
rect 128228 182260 166448 182288
rect 128228 182248 128234 182260
rect 166442 182248 166448 182260
rect 166500 182248 166506 182300
rect 114370 182180 114376 182232
rect 114428 182220 114434 182232
rect 169202 182220 169208 182232
rect 114428 182192 169208 182220
rect 114428 182180 114434 182192
rect 169202 182180 169208 182192
rect 169260 182180 169266 182232
rect 215938 181636 215944 181688
rect 215996 181676 216002 181688
rect 259638 181676 259644 181688
rect 215996 181648 259644 181676
rect 215996 181636 216002 181648
rect 259638 181636 259644 181648
rect 259696 181636 259702 181688
rect 202138 181568 202144 181620
rect 202196 181608 202202 181620
rect 259454 181608 259460 181620
rect 202196 181580 259460 181608
rect 202196 181568 202202 181580
rect 259454 181568 259460 181580
rect 259512 181568 259518 181620
rect 174538 181500 174544 181552
rect 174596 181540 174602 181552
rect 265066 181540 265072 181552
rect 174596 181512 265072 181540
rect 174596 181500 174602 181512
rect 265066 181500 265072 181512
rect 265124 181500 265130 181552
rect 291838 181500 291844 181552
rect 291896 181540 291902 181552
rect 332686 181540 332692 181552
rect 291896 181512 332692 181540
rect 291896 181500 291902 181512
rect 332686 181500 332692 181512
rect 332744 181500 332750 181552
rect 66162 181432 66168 181484
rect 66220 181472 66226 181484
rect 251450 181472 251456 181484
rect 66220 181444 251456 181472
rect 66220 181432 66226 181444
rect 251450 181432 251456 181444
rect 251508 181432 251514 181484
rect 283558 181432 283564 181484
rect 283616 181472 283622 181484
rect 343818 181472 343824 181484
rect 283616 181444 343824 181472
rect 283616 181432 283622 181444
rect 343818 181432 343824 181444
rect 343876 181432 343882 181484
rect 112162 180956 112168 181008
rect 112220 180996 112226 181008
rect 167730 180996 167736 181008
rect 112220 180968 167736 180996
rect 112220 180956 112226 180968
rect 167730 180956 167736 180968
rect 167788 180956 167794 181008
rect 110690 180888 110696 180940
rect 110748 180928 110754 180940
rect 169110 180928 169116 180940
rect 110748 180900 169116 180928
rect 110748 180888 110754 180900
rect 169110 180888 169116 180900
rect 169168 180888 169174 180940
rect 125042 180820 125048 180872
rect 125100 180860 125106 180872
rect 211798 180860 211804 180872
rect 125100 180832 211804 180860
rect 125100 180820 125106 180832
rect 211798 180820 211804 180832
rect 211856 180820 211862 180872
rect 220078 180276 220084 180328
rect 220136 180316 220142 180328
rect 258442 180316 258448 180328
rect 220136 180288 258448 180316
rect 220136 180276 220142 180288
rect 258442 180276 258448 180288
rect 258500 180276 258506 180328
rect 287698 180276 287704 180328
rect 287756 180316 287762 180328
rect 335538 180316 335544 180328
rect 287756 180288 335544 180316
rect 287756 180276 287762 180288
rect 335538 180276 335544 180288
rect 335596 180276 335602 180328
rect 113358 180208 113364 180260
rect 113416 180248 113422 180260
rect 336918 180248 336924 180260
rect 113416 180220 336924 180248
rect 113416 180208 113422 180220
rect 336918 180208 336924 180220
rect 336976 180208 336982 180260
rect 71774 180140 71780 180192
rect 71832 180180 71838 180192
rect 339678 180180 339684 180192
rect 71832 180152 339684 180180
rect 71832 180140 71838 180152
rect 339678 180140 339684 180152
rect 339736 180140 339742 180192
rect 64690 180072 64696 180124
rect 64748 180112 64754 180124
rect 342530 180112 342536 180124
rect 64748 180084 342536 180112
rect 64748 180072 64754 180084
rect 342530 180072 342536 180084
rect 342588 180072 342594 180124
rect 133138 179528 133144 179580
rect 133196 179568 133202 179580
rect 165062 179568 165068 179580
rect 133196 179540 165068 179568
rect 133196 179528 133202 179540
rect 165062 179528 165068 179540
rect 165120 179528 165126 179580
rect 121178 179460 121184 179512
rect 121236 179500 121242 179512
rect 166350 179500 166356 179512
rect 121236 179472 166356 179500
rect 121236 179460 121242 179472
rect 166350 179460 166356 179472
rect 166408 179460 166414 179512
rect 110046 179392 110052 179444
rect 110104 179432 110110 179444
rect 214742 179432 214748 179444
rect 110104 179404 214748 179432
rect 110104 179392 110110 179404
rect 214742 179392 214748 179404
rect 214800 179392 214806 179444
rect 347038 179324 347044 179376
rect 347096 179364 347102 179376
rect 579982 179364 579988 179376
rect 347096 179336 579988 179364
rect 347096 179324 347102 179336
rect 579982 179324 579988 179336
rect 580040 179324 580046 179376
rect 238018 179052 238024 179104
rect 238076 179092 238082 179104
rect 258350 179092 258356 179104
rect 238076 179064 258356 179092
rect 238076 179052 238082 179064
rect 258350 179052 258356 179064
rect 258408 179052 258414 179104
rect 225598 178916 225604 178968
rect 225656 178956 225662 178968
rect 258258 178956 258264 178968
rect 225656 178928 258264 178956
rect 225656 178916 225662 178928
rect 258258 178916 258264 178928
rect 258316 178916 258322 178968
rect 229738 178848 229744 178900
rect 229796 178888 229802 178900
rect 258074 178888 258080 178900
rect 229796 178860 258080 178888
rect 229796 178848 229802 178860
rect 258074 178848 258080 178860
rect 258132 178848 258138 178900
rect 206278 178780 206284 178832
rect 206336 178820 206342 178832
rect 249058 178820 249064 178832
rect 206336 178792 249064 178820
rect 206336 178780 206342 178792
rect 249058 178780 249064 178792
rect 249116 178780 249122 178832
rect 184198 178712 184204 178764
rect 184256 178752 184262 178764
rect 242802 178752 242808 178764
rect 184256 178724 242808 178752
rect 184256 178712 184262 178724
rect 242802 178712 242808 178724
rect 242860 178712 242866 178764
rect 311158 178712 311164 178764
rect 311216 178752 311222 178764
rect 335446 178752 335452 178764
rect 311216 178724 335452 178752
rect 311216 178712 311222 178724
rect 335446 178712 335452 178724
rect 335504 178712 335510 178764
rect 70394 178644 70400 178696
rect 70452 178684 70458 178696
rect 328730 178684 328736 178696
rect 70452 178656 328736 178684
rect 70452 178644 70458 178656
rect 328730 178644 328736 178656
rect 328788 178644 328794 178696
rect 148226 178304 148232 178356
rect 148284 178344 148290 178356
rect 169018 178344 169024 178356
rect 148284 178316 169024 178344
rect 148284 178304 148290 178316
rect 169018 178304 169024 178316
rect 169076 178304 169082 178356
rect 134702 178236 134708 178288
rect 134760 178276 134766 178288
rect 165430 178276 165436 178288
rect 134760 178248 165436 178276
rect 134760 178236 134766 178248
rect 165430 178236 165436 178248
rect 165488 178236 165494 178288
rect 115842 178168 115848 178220
rect 115900 178208 115906 178220
rect 166258 178208 166264 178220
rect 115900 178180 166264 178208
rect 115900 178168 115906 178180
rect 166258 178168 166264 178180
rect 166316 178168 166322 178220
rect 99098 178100 99104 178152
rect 99156 178140 99162 178152
rect 170490 178140 170496 178152
rect 99156 178112 170496 178140
rect 99156 178100 99162 178112
rect 170490 178100 170496 178112
rect 170548 178100 170554 178152
rect 129458 178032 129464 178084
rect 129516 178072 129522 178084
rect 208394 178072 208400 178084
rect 129516 178044 208400 178072
rect 129516 178032 129522 178044
rect 208394 178032 208400 178044
rect 208452 178032 208458 178084
rect 242802 177624 242808 177676
rect 242860 177664 242866 177676
rect 261018 177664 261024 177676
rect 242860 177636 261024 177664
rect 242860 177624 242866 177636
rect 261018 177624 261024 177636
rect 261076 177624 261082 177676
rect 232498 177556 232504 177608
rect 232556 177596 232562 177608
rect 259730 177596 259736 177608
rect 232556 177568 259736 177596
rect 232556 177556 232562 177568
rect 259730 177556 259736 177568
rect 259788 177556 259794 177608
rect 314010 177556 314016 177608
rect 314068 177596 314074 177608
rect 334066 177596 334072 177608
rect 314068 177568 334072 177596
rect 314068 177556 314074 177568
rect 334066 177556 334072 177568
rect 334124 177556 334130 177608
rect 239398 177488 239404 177540
rect 239456 177528 239462 177540
rect 267826 177528 267832 177540
rect 239456 177500 267832 177528
rect 239456 177488 239462 177500
rect 267826 177488 267832 177500
rect 267884 177488 267890 177540
rect 318058 177488 318064 177540
rect 318116 177528 318122 177540
rect 338298 177528 338304 177540
rect 318116 177500 338304 177528
rect 318116 177488 318122 177500
rect 338298 177488 338304 177500
rect 338356 177488 338362 177540
rect 228358 177420 228364 177472
rect 228416 177460 228422 177472
rect 266538 177460 266544 177472
rect 228416 177432 266544 177460
rect 228416 177420 228422 177432
rect 266538 177420 266544 177432
rect 266596 177420 266602 177472
rect 311250 177420 311256 177472
rect 311308 177460 311314 177472
rect 331490 177460 331496 177472
rect 311308 177432 331496 177460
rect 311308 177420 311314 177432
rect 331490 177420 331496 177432
rect 331548 177420 331554 177472
rect 203518 177352 203524 177404
rect 203576 177392 203582 177404
rect 249242 177392 249248 177404
rect 203576 177364 249248 177392
rect 203576 177352 203582 177364
rect 249242 177352 249248 177364
rect 249300 177352 249306 177404
rect 307018 177352 307024 177404
rect 307076 177392 307082 177404
rect 341150 177392 341156 177404
rect 307076 177364 341156 177392
rect 307076 177352 307082 177364
rect 341150 177352 341156 177364
rect 341208 177352 341214 177404
rect 170398 177284 170404 177336
rect 170456 177324 170462 177336
rect 321370 177324 321376 177336
rect 170456 177296 321376 177324
rect 170456 177284 170462 177296
rect 321370 177284 321376 177296
rect 321428 177284 321434 177336
rect 132034 176944 132040 176996
rect 132092 176984 132098 176996
rect 165522 176984 165528 176996
rect 132092 176956 165528 176984
rect 132092 176944 132098 176956
rect 165522 176944 165528 176956
rect 165580 176944 165586 176996
rect 108114 176876 108120 176928
rect 108172 176916 108178 176928
rect 170674 176916 170680 176928
rect 108172 176888 170680 176916
rect 108172 176876 108178 176888
rect 170674 176876 170680 176888
rect 170732 176876 170738 176928
rect 102042 176808 102048 176860
rect 102100 176848 102106 176860
rect 171870 176848 171876 176860
rect 102100 176820 171876 176848
rect 102100 176808 102106 176820
rect 171870 176808 171876 176820
rect 171928 176808 171934 176860
rect 135714 176740 135720 176792
rect 135772 176780 135778 176792
rect 213914 176780 213920 176792
rect 135772 176752 213920 176780
rect 135772 176740 135778 176752
rect 213914 176740 213920 176752
rect 213972 176740 213978 176792
rect 127066 176672 127072 176724
rect 127124 176712 127130 176724
rect 211982 176712 211988 176724
rect 127124 176684 211988 176712
rect 127124 176672 127130 176684
rect 211982 176672 211988 176684
rect 212040 176672 212046 176724
rect 196618 176604 196624 176656
rect 196676 176644 196682 176656
rect 248046 176644 248052 176656
rect 196676 176616 248052 176644
rect 196676 176604 196682 176616
rect 248046 176604 248052 176616
rect 248104 176604 248110 176656
rect 249150 176644 249156 176656
rect 248386 176616 249156 176644
rect 242158 176536 242164 176588
rect 242216 176576 242222 176588
rect 248386 176576 248414 176616
rect 249150 176604 249156 176616
rect 249208 176604 249214 176656
rect 309870 176604 309876 176656
rect 309928 176644 309934 176656
rect 321462 176644 321468 176656
rect 309928 176616 321468 176644
rect 309928 176604 309934 176616
rect 321462 176604 321468 176616
rect 321520 176604 321526 176656
rect 242216 176548 248414 176576
rect 242216 176536 242222 176548
rect 121914 176196 121920 176248
rect 121972 176236 121978 176248
rect 167914 176236 167920 176248
rect 121972 176208 167920 176236
rect 121972 176196 121978 176208
rect 167914 176196 167920 176208
rect 167972 176196 167978 176248
rect 119430 176128 119436 176180
rect 119488 176168 119494 176180
rect 166534 176168 166540 176180
rect 119488 176140 166540 176168
rect 119488 176128 119494 176140
rect 166534 176128 166540 176140
rect 166592 176128 166598 176180
rect 158898 176060 158904 176112
rect 158956 176100 158962 176112
rect 214558 176100 214564 176112
rect 158956 176072 214564 176100
rect 158956 176060 158962 176072
rect 214558 176060 214564 176072
rect 214616 176060 214622 176112
rect 130746 175992 130752 176044
rect 130804 176032 130810 176044
rect 214098 176032 214104 176044
rect 130804 176004 214104 176032
rect 130804 175992 130810 176004
rect 214098 175992 214104 176004
rect 214156 175992 214162 176044
rect 242250 175992 242256 176044
rect 242308 176032 242314 176044
rect 255590 176032 255596 176044
rect 242308 176004 255596 176032
rect 242308 175992 242314 176004
rect 255590 175992 255596 176004
rect 255648 175992 255654 176044
rect 315298 175992 315304 176044
rect 315356 176032 315362 176044
rect 332594 176032 332600 176044
rect 315356 176004 332600 176032
rect 315356 175992 315362 176004
rect 332594 175992 332600 176004
rect 332652 175992 332658 176044
rect 100754 175924 100760 175976
rect 100812 175964 100818 175976
rect 210510 175964 210516 175976
rect 100812 175936 210516 175964
rect 100812 175924 100818 175936
rect 210510 175924 210516 175936
rect 210568 175924 210574 175976
rect 246298 175924 246304 175976
rect 246356 175964 246362 175976
rect 262490 175964 262496 175976
rect 246356 175936 262496 175964
rect 246356 175924 246362 175936
rect 262490 175924 262496 175936
rect 262548 175924 262554 175976
rect 318242 175924 318248 175976
rect 318300 175964 318306 175976
rect 335630 175964 335636 175976
rect 318300 175936 335636 175964
rect 318300 175924 318306 175936
rect 335630 175924 335636 175936
rect 335688 175924 335694 175976
rect 318150 175584 318156 175636
rect 318208 175624 318214 175636
rect 321462 175624 321468 175636
rect 318208 175596 321468 175624
rect 318208 175584 318214 175596
rect 321462 175584 321468 175596
rect 321520 175584 321526 175636
rect 165430 175176 165436 175228
rect 165488 175216 165494 175228
rect 213914 175216 213920 175228
rect 165488 175188 213920 175216
rect 165488 175176 165494 175188
rect 213914 175176 213920 175188
rect 213972 175176 213978 175228
rect 165062 175108 165068 175160
rect 165120 175148 165126 175160
rect 214006 175148 214012 175160
rect 165120 175120 214012 175148
rect 165120 175108 165126 175120
rect 214006 175108 214012 175120
rect 214064 175108 214070 175160
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 39298 164200 39304 164212
rect 3292 164172 39304 164200
rect 3292 164160 3298 164172
rect 39298 164160 39304 164172
rect 39356 164160 39362 164212
rect 3418 150356 3424 150408
rect 3476 150396 3482 150408
rect 25498 150396 25504 150408
rect 3476 150368 25504 150396
rect 3476 150356 3482 150368
rect 25498 150356 25504 150368
rect 25556 150356 25562 150408
rect 3234 137912 3240 137964
rect 3292 137952 3298 137964
rect 14458 137952 14464 137964
rect 3292 137924 14464 137952
rect 3292 137912 3298 137924
rect 14458 137912 14464 137924
rect 14516 137912 14522 137964
rect 63402 122816 63408 122868
rect 63460 122856 63466 122868
rect 66070 122856 66076 122868
rect 63460 122828 66076 122856
rect 63460 122816 63466 122828
rect 66070 122816 66076 122828
rect 66128 122816 66134 122868
rect 3418 111732 3424 111784
rect 3476 111772 3482 111784
rect 13078 111772 13084 111784
rect 3476 111744 13084 111772
rect 3476 111732 3482 111744
rect 13078 111732 13084 111744
rect 13136 111732 13142 111784
rect 2774 97724 2780 97776
rect 2832 97764 2838 97776
rect 4798 97764 4804 97776
rect 2832 97736 4804 97764
rect 2832 97724 2838 97736
rect 4798 97724 4804 97736
rect 4856 97724 4862 97776
rect 291838 174020 291844 174072
rect 291896 174060 291902 174072
rect 307662 174060 307668 174072
rect 291896 174032 307668 174060
rect 291896 174020 291902 174032
rect 307662 174020 307668 174032
rect 307720 174020 307726 174072
rect 278222 173952 278228 174004
rect 278280 173992 278286 174004
rect 306742 173992 306748 174004
rect 278280 173964 306748 173992
rect 278280 173952 278286 173964
rect 306742 173952 306748 173964
rect 306800 173952 306806 174004
rect 266998 173884 267004 173936
rect 267056 173924 267062 173936
rect 307570 173924 307576 173936
rect 267056 173896 307576 173924
rect 267056 173884 267062 173896
rect 307570 173884 307576 173896
rect 307628 173884 307634 173936
rect 165522 173816 165528 173868
rect 165580 173856 165586 173868
rect 213914 173856 213920 173868
rect 165580 173828 213920 173856
rect 165580 173816 165586 173828
rect 213914 173816 213920 173828
rect 213972 173816 213978 173868
rect 251818 172660 251824 172712
rect 251876 172700 251882 172712
rect 259454 172700 259460 172712
rect 251876 172672 259460 172700
rect 251876 172660 251882 172672
rect 259454 172660 259460 172672
rect 259512 172660 259518 172712
rect 282178 172660 282184 172712
rect 282236 172700 282242 172712
rect 307294 172700 307300 172712
rect 282236 172672 307300 172700
rect 282236 172660 282242 172672
rect 307294 172660 307300 172672
rect 307352 172660 307358 172712
rect 273990 172592 273996 172644
rect 274048 172632 274054 172644
rect 307662 172632 307668 172644
rect 274048 172604 307668 172632
rect 274048 172592 274054 172604
rect 307662 172592 307668 172604
rect 307720 172592 307726 172644
rect 260282 172524 260288 172576
rect 260340 172564 260346 172576
rect 306926 172564 306932 172576
rect 260340 172536 306932 172564
rect 260340 172524 260346 172536
rect 306926 172524 306932 172536
rect 306984 172524 306990 172576
rect 166442 172456 166448 172508
rect 166500 172496 166506 172508
rect 214006 172496 214012 172508
rect 166500 172468 214012 172496
rect 166500 172456 166506 172468
rect 214006 172456 214012 172468
rect 214064 172456 214070 172508
rect 252002 172456 252008 172508
rect 252060 172496 252066 172508
rect 258074 172496 258080 172508
rect 252060 172468 258080 172496
rect 252060 172456 252066 172468
rect 258074 172456 258080 172468
rect 258132 172456 258138 172508
rect 208394 172388 208400 172440
rect 208452 172428 208458 172440
rect 213914 172428 213920 172440
rect 208452 172400 213920 172428
rect 208452 172388 208458 172400
rect 213914 172388 213920 172400
rect 213972 172388 213978 172440
rect 252462 172388 252468 172440
rect 252520 172428 252526 172440
rect 261110 172428 261116 172440
rect 252520 172400 261116 172428
rect 252520 172388 252526 172400
rect 261110 172388 261116 172400
rect 261168 172388 261174 172440
rect 258074 172320 258080 172372
rect 258132 172360 258138 172372
rect 258258 172360 258264 172372
rect 258132 172332 258264 172360
rect 258132 172320 258138 172332
rect 258258 172320 258264 172332
rect 258316 172320 258322 172372
rect 258258 172184 258264 172236
rect 258316 172224 258322 172236
rect 258442 172224 258448 172236
rect 258316 172196 258448 172224
rect 258316 172184 258322 172196
rect 258442 172184 258448 172196
rect 258500 172184 258506 172236
rect 289262 171232 289268 171284
rect 289320 171272 289326 171284
rect 307478 171272 307484 171284
rect 289320 171244 307484 171272
rect 289320 171232 289326 171244
rect 307478 171232 307484 171244
rect 307536 171232 307542 171284
rect 264330 171164 264336 171216
rect 264388 171204 264394 171216
rect 307570 171204 307576 171216
rect 264388 171176 307576 171204
rect 264388 171164 264394 171176
rect 307570 171164 307576 171176
rect 307628 171164 307634 171216
rect 261754 171096 261760 171148
rect 261812 171136 261818 171148
rect 307662 171136 307668 171148
rect 261812 171108 307668 171136
rect 261812 171096 261818 171108
rect 307662 171096 307668 171108
rect 307720 171096 307726 171148
rect 171962 171028 171968 171080
rect 172020 171068 172026 171080
rect 213914 171068 213920 171080
rect 172020 171040 213920 171068
rect 172020 171028 172026 171040
rect 213914 171028 213920 171040
rect 213972 171028 213978 171080
rect 252094 171028 252100 171080
rect 252152 171068 252158 171080
rect 262214 171068 262220 171080
rect 252152 171040 262220 171068
rect 252152 171028 252158 171040
rect 262214 171028 262220 171040
rect 262272 171028 262278 171080
rect 211982 170960 211988 171012
rect 212040 171000 212046 171012
rect 214006 171000 214012 171012
rect 212040 170972 214012 171000
rect 212040 170960 212046 170972
rect 214006 170960 214012 170972
rect 214064 170960 214070 171012
rect 252462 170892 252468 170944
rect 252520 170932 252526 170944
rect 256970 170932 256976 170944
rect 252520 170904 256976 170932
rect 252520 170892 252526 170904
rect 256970 170892 256976 170904
rect 257028 170892 257034 170944
rect 251818 169940 251824 169992
rect 251876 169980 251882 169992
rect 258166 169980 258172 169992
rect 251876 169952 258172 169980
rect 251876 169940 251882 169952
rect 258166 169940 258172 169952
rect 258224 169940 258230 169992
rect 287882 169872 287888 169924
rect 287940 169912 287946 169924
rect 306926 169912 306932 169924
rect 287940 169884 306932 169912
rect 287940 169872 287946 169884
rect 306926 169872 306932 169884
rect 306984 169872 306990 169924
rect 271322 169804 271328 169856
rect 271380 169844 271386 169856
rect 307478 169844 307484 169856
rect 271380 169816 307484 169844
rect 271380 169804 271386 169816
rect 307478 169804 307484 169816
rect 307536 169804 307542 169856
rect 258810 169736 258816 169788
rect 258868 169776 258874 169788
rect 307662 169776 307668 169788
rect 258868 169748 307668 169776
rect 258868 169736 258874 169748
rect 307662 169736 307668 169748
rect 307720 169736 307726 169788
rect 167822 169668 167828 169720
rect 167880 169708 167886 169720
rect 213914 169708 213920 169720
rect 167880 169680 213920 169708
rect 167880 169668 167886 169680
rect 213914 169668 213920 169680
rect 213972 169668 213978 169720
rect 324314 169668 324320 169720
rect 324372 169708 324378 169720
rect 332594 169708 332600 169720
rect 324372 169680 332600 169708
rect 324372 169668 324378 169680
rect 332594 169668 332600 169680
rect 332652 169668 332658 169720
rect 211798 169600 211804 169652
rect 211856 169640 211862 169652
rect 214006 169640 214012 169652
rect 211856 169612 214012 169640
rect 211856 169600 211862 169612
rect 214006 169600 214012 169612
rect 214064 169600 214070 169652
rect 252002 169192 252008 169244
rect 252060 169232 252066 169244
rect 258074 169232 258080 169244
rect 252060 169204 258080 169232
rect 252060 169192 252066 169204
rect 258074 169192 258080 169204
rect 258132 169192 258138 169244
rect 283558 168512 283564 168564
rect 283616 168552 283622 168564
rect 307294 168552 307300 168564
rect 283616 168524 307300 168552
rect 283616 168512 283622 168524
rect 307294 168512 307300 168524
rect 307352 168512 307358 168564
rect 252462 168444 252468 168496
rect 252520 168484 252526 168496
rect 259546 168484 259552 168496
rect 252520 168456 259552 168484
rect 252520 168444 252526 168456
rect 259546 168444 259552 168456
rect 259604 168444 259610 168496
rect 279602 168444 279608 168496
rect 279660 168484 279666 168496
rect 307478 168484 307484 168496
rect 279660 168456 307484 168484
rect 279660 168444 279666 168456
rect 307478 168444 307484 168456
rect 307536 168444 307542 168496
rect 264238 168376 264244 168428
rect 264296 168416 264302 168428
rect 307662 168416 307668 168428
rect 264296 168388 307668 168416
rect 264296 168376 264302 168388
rect 307662 168376 307668 168388
rect 307720 168376 307726 168428
rect 166350 168308 166356 168360
rect 166408 168348 166414 168360
rect 214006 168348 214012 168360
rect 166408 168320 214012 168348
rect 166408 168308 166414 168320
rect 214006 168308 214012 168320
rect 214064 168308 214070 168360
rect 252094 168308 252100 168360
rect 252152 168348 252158 168360
rect 260926 168348 260932 168360
rect 252152 168320 260932 168348
rect 252152 168308 252158 168320
rect 260926 168308 260932 168320
rect 260984 168308 260990 168360
rect 324406 168308 324412 168360
rect 324464 168348 324470 168360
rect 338390 168348 338396 168360
rect 324464 168320 338396 168348
rect 324464 168308 324470 168320
rect 338390 168308 338396 168320
rect 338448 168308 338454 168360
rect 167914 168240 167920 168292
rect 167972 168280 167978 168292
rect 213914 168280 213920 168292
rect 167972 168252 213920 168280
rect 167972 168240 167978 168252
rect 213914 168240 213920 168252
rect 213972 168240 213978 168292
rect 324314 168240 324320 168292
rect 324372 168280 324378 168292
rect 334250 168280 334256 168292
rect 324372 168252 334256 168280
rect 324372 168240 324378 168252
rect 334250 168240 334256 168252
rect 334308 168240 334314 168292
rect 251910 168172 251916 168224
rect 251968 168212 251974 168224
rect 255314 168212 255320 168224
rect 251968 168184 255320 168212
rect 251968 168172 251974 168184
rect 255314 168172 255320 168184
rect 255372 168172 255378 168224
rect 252462 168036 252468 168088
rect 252520 168076 252526 168088
rect 259638 168076 259644 168088
rect 252520 168048 259644 168076
rect 252520 168036 252526 168048
rect 259638 168036 259644 168048
rect 259696 168036 259702 168088
rect 283650 167152 283656 167204
rect 283708 167192 283714 167204
rect 307662 167192 307668 167204
rect 283708 167164 307668 167192
rect 283708 167152 283714 167164
rect 307662 167152 307668 167164
rect 307720 167152 307726 167204
rect 272518 167084 272524 167136
rect 272576 167124 272582 167136
rect 307478 167124 307484 167136
rect 272576 167096 307484 167124
rect 272576 167084 272582 167096
rect 307478 167084 307484 167096
rect 307536 167084 307542 167136
rect 265894 167016 265900 167068
rect 265952 167056 265958 167068
rect 307570 167056 307576 167068
rect 265952 167028 307576 167056
rect 265952 167016 265958 167028
rect 307570 167016 307576 167028
rect 307628 167016 307634 167068
rect 166534 166948 166540 167000
rect 166592 166988 166598 167000
rect 213914 166988 213920 167000
rect 166592 166960 213920 166988
rect 166592 166948 166598 166960
rect 213914 166948 213920 166960
rect 213972 166948 213978 167000
rect 324314 166948 324320 167000
rect 324372 166988 324378 167000
rect 345290 166988 345296 167000
rect 324372 166960 345296 166988
rect 324372 166948 324378 166960
rect 345290 166948 345296 166960
rect 345348 166948 345354 167000
rect 170582 166880 170588 166932
rect 170640 166920 170646 166932
rect 214006 166920 214012 166932
rect 170640 166892 214012 166920
rect 170640 166880 170646 166892
rect 214006 166880 214012 166892
rect 214064 166880 214070 166932
rect 251818 166880 251824 166932
rect 251876 166920 251882 166932
rect 260834 166920 260840 166932
rect 251876 166892 260840 166920
rect 251876 166880 251882 166892
rect 260834 166880 260840 166892
rect 260892 166880 260898 166932
rect 293218 165724 293224 165776
rect 293276 165764 293282 165776
rect 307294 165764 307300 165776
rect 293276 165736 307300 165764
rect 293276 165724 293282 165736
rect 307294 165724 307300 165736
rect 307352 165724 307358 165776
rect 271138 165656 271144 165708
rect 271196 165696 271202 165708
rect 307662 165696 307668 165708
rect 271196 165668 307668 165696
rect 271196 165656 271202 165668
rect 307662 165656 307668 165668
rect 307720 165656 307726 165708
rect 261662 165588 261668 165640
rect 261720 165628 261726 165640
rect 307478 165628 307484 165640
rect 261720 165600 307484 165628
rect 261720 165588 261726 165600
rect 307478 165588 307484 165600
rect 307536 165588 307542 165640
rect 166258 165520 166264 165572
rect 166316 165560 166322 165572
rect 213914 165560 213920 165572
rect 166316 165532 213920 165560
rect 166316 165520 166322 165532
rect 213914 165520 213920 165532
rect 213972 165520 213978 165572
rect 169202 165452 169208 165504
rect 169260 165492 169266 165504
rect 214006 165492 214012 165504
rect 169260 165464 214012 165492
rect 169260 165452 169266 165464
rect 214006 165452 214012 165464
rect 214064 165452 214070 165504
rect 252462 165452 252468 165504
rect 252520 165492 252526 165504
rect 261018 165492 261024 165504
rect 252520 165464 261024 165492
rect 252520 165452 252526 165464
rect 261018 165452 261024 165464
rect 261076 165452 261082 165504
rect 252370 165384 252376 165436
rect 252428 165424 252434 165436
rect 266446 165424 266452 165436
rect 252428 165396 266452 165424
rect 252428 165384 252434 165396
rect 266446 165384 266452 165396
rect 266504 165384 266510 165436
rect 251358 164976 251364 165028
rect 251416 165016 251422 165028
rect 252830 165016 252836 165028
rect 251416 164988 252836 165016
rect 251416 164976 251422 164988
rect 252830 164976 252836 164988
rect 252888 164976 252894 165028
rect 265802 164432 265808 164484
rect 265860 164472 265866 164484
rect 307662 164472 307668 164484
rect 265860 164444 307668 164472
rect 265860 164432 265866 164444
rect 307662 164432 307668 164444
rect 307720 164432 307726 164484
rect 294782 164364 294788 164416
rect 294840 164404 294846 164416
rect 307570 164404 307576 164416
rect 294840 164376 307576 164404
rect 294840 164364 294846 164376
rect 307570 164364 307576 164376
rect 307628 164364 307634 164416
rect 269850 164296 269856 164348
rect 269908 164336 269914 164348
rect 307478 164336 307484 164348
rect 269908 164308 307484 164336
rect 269908 164296 269914 164308
rect 307478 164296 307484 164308
rect 307536 164296 307542 164348
rect 304350 164228 304356 164280
rect 304408 164268 304414 164280
rect 306558 164268 306564 164280
rect 304408 164240 306564 164268
rect 304408 164228 304414 164240
rect 306558 164228 306564 164240
rect 306616 164228 306622 164280
rect 167730 164160 167736 164212
rect 167788 164200 167794 164212
rect 213914 164200 213920 164212
rect 167788 164172 213920 164200
rect 167788 164160 167794 164172
rect 213914 164160 213920 164172
rect 213972 164160 213978 164212
rect 252462 164160 252468 164212
rect 252520 164200 252526 164212
rect 267918 164200 267924 164212
rect 252520 164172 267924 164200
rect 252520 164160 252526 164172
rect 267918 164160 267924 164172
rect 267976 164160 267982 164212
rect 324406 164160 324412 164212
rect 324464 164200 324470 164212
rect 345198 164200 345204 164212
rect 324464 164172 345204 164200
rect 324464 164160 324470 164172
rect 345198 164160 345204 164172
rect 345256 164160 345262 164212
rect 324314 164092 324320 164144
rect 324372 164132 324378 164144
rect 335630 164132 335636 164144
rect 324372 164104 335636 164132
rect 324372 164092 324378 164104
rect 335630 164092 335636 164104
rect 335688 164092 335694 164144
rect 251358 163072 251364 163124
rect 251416 163112 251422 163124
rect 254026 163112 254032 163124
rect 251416 163084 254032 163112
rect 251416 163072 251422 163084
rect 254026 163072 254032 163084
rect 254084 163072 254090 163124
rect 300118 163004 300124 163056
rect 300176 163044 300182 163056
rect 307478 163044 307484 163056
rect 300176 163016 307484 163044
rect 300176 163004 300182 163016
rect 307478 163004 307484 163016
rect 307536 163004 307542 163056
rect 268378 162936 268384 162988
rect 268436 162976 268442 162988
rect 307662 162976 307668 162988
rect 268436 162948 307668 162976
rect 268436 162936 268442 162948
rect 307662 162936 307668 162948
rect 307720 162936 307726 162988
rect 261570 162868 261576 162920
rect 261628 162908 261634 162920
rect 307294 162908 307300 162920
rect 261628 162880 307300 162908
rect 261628 162868 261634 162880
rect 307294 162868 307300 162880
rect 307352 162868 307358 162920
rect 169110 162800 169116 162852
rect 169168 162840 169174 162852
rect 213914 162840 213920 162852
rect 169168 162812 213920 162840
rect 169168 162800 169174 162812
rect 213914 162800 213920 162812
rect 213972 162800 213978 162852
rect 252462 162800 252468 162852
rect 252520 162840 252526 162852
rect 269298 162840 269304 162852
rect 252520 162812 269304 162840
rect 252520 162800 252526 162812
rect 269298 162800 269304 162812
rect 269356 162800 269362 162852
rect 324314 162800 324320 162852
rect 324372 162840 324378 162852
rect 336734 162840 336740 162852
rect 324372 162812 336740 162840
rect 324372 162800 324378 162812
rect 336734 162800 336740 162812
rect 336792 162800 336798 162852
rect 252094 162732 252100 162784
rect 252152 162772 252158 162784
rect 264974 162772 264980 162784
rect 252152 162744 264980 162772
rect 252152 162732 252158 162744
rect 264974 162732 264980 162744
rect 265032 162732 265038 162784
rect 324406 162732 324412 162784
rect 324464 162772 324470 162784
rect 331490 162772 331496 162784
rect 324464 162744 331496 162772
rect 324464 162732 324470 162744
rect 331490 162732 331496 162744
rect 331548 162732 331554 162784
rect 296070 161576 296076 161628
rect 296128 161616 296134 161628
rect 307478 161616 307484 161628
rect 296128 161588 307484 161616
rect 296128 161576 296134 161588
rect 307478 161576 307484 161588
rect 307536 161576 307542 161628
rect 269758 161508 269764 161560
rect 269816 161548 269822 161560
rect 307294 161548 307300 161560
rect 269816 161520 307300 161548
rect 269816 161508 269822 161520
rect 307294 161508 307300 161520
rect 307352 161508 307358 161560
rect 260190 161440 260196 161492
rect 260248 161480 260254 161492
rect 307662 161480 307668 161492
rect 260248 161452 307668 161480
rect 260248 161440 260254 161452
rect 307662 161440 307668 161452
rect 307720 161440 307726 161492
rect 170674 161372 170680 161424
rect 170732 161412 170738 161424
rect 213914 161412 213920 161424
rect 170732 161384 213920 161412
rect 170732 161372 170738 161384
rect 213914 161372 213920 161384
rect 213972 161372 213978 161424
rect 252462 161372 252468 161424
rect 252520 161412 252526 161424
rect 266354 161412 266360 161424
rect 252520 161384 266360 161412
rect 252520 161372 252526 161384
rect 266354 161372 266360 161384
rect 266412 161372 266418 161424
rect 324682 161372 324688 161424
rect 324740 161412 324746 161424
rect 339770 161412 339776 161424
rect 324740 161384 339776 161412
rect 324740 161372 324746 161384
rect 339770 161372 339776 161384
rect 339828 161372 339834 161424
rect 207750 161304 207756 161356
rect 207808 161344 207814 161356
rect 214006 161344 214012 161356
rect 207808 161316 214012 161344
rect 207808 161304 207814 161316
rect 214006 161304 214012 161316
rect 214064 161304 214070 161356
rect 324314 161304 324320 161356
rect 324372 161344 324378 161356
rect 335354 161344 335360 161356
rect 324372 161316 335360 161344
rect 324372 161304 324378 161316
rect 335354 161304 335360 161316
rect 335412 161304 335418 161356
rect 252002 160828 252008 160880
rect 252060 160868 252066 160880
rect 255406 160868 255412 160880
rect 252060 160840 255412 160868
rect 252060 160828 252066 160840
rect 255406 160828 255412 160840
rect 255464 160828 255470 160880
rect 171870 160692 171876 160744
rect 171928 160732 171934 160744
rect 213914 160732 213920 160744
rect 171928 160704 213920 160732
rect 171928 160692 171934 160704
rect 213914 160692 213920 160704
rect 213972 160692 213978 160744
rect 285030 160692 285036 160744
rect 285088 160732 285094 160744
rect 307202 160732 307208 160744
rect 285088 160704 307208 160732
rect 285088 160692 285094 160704
rect 307202 160692 307208 160704
rect 307260 160692 307266 160744
rect 252094 160284 252100 160336
rect 252152 160324 252158 160336
rect 258258 160324 258264 160336
rect 252152 160296 258264 160324
rect 252152 160284 252158 160296
rect 258258 160284 258264 160296
rect 258316 160284 258322 160336
rect 265710 160148 265716 160200
rect 265768 160188 265774 160200
rect 307662 160188 307668 160200
rect 265768 160160 307668 160188
rect 265768 160148 265774 160160
rect 307662 160148 307668 160160
rect 307720 160148 307726 160200
rect 258718 160080 258724 160132
rect 258776 160120 258782 160132
rect 306558 160120 306564 160132
rect 258776 160092 306564 160120
rect 258776 160080 258782 160092
rect 306558 160080 306564 160092
rect 306616 160080 306622 160132
rect 211890 160012 211896 160064
rect 211948 160052 211954 160064
rect 214466 160052 214472 160064
rect 211948 160024 214472 160052
rect 211948 160012 211954 160024
rect 214466 160012 214472 160024
rect 214524 160012 214530 160064
rect 252462 160012 252468 160064
rect 252520 160052 252526 160064
rect 262490 160052 262496 160064
rect 252520 160024 262496 160052
rect 252520 160012 252526 160024
rect 262490 160012 262496 160024
rect 262548 160012 262554 160064
rect 324314 160012 324320 160064
rect 324372 160052 324378 160064
rect 328730 160052 328736 160064
rect 324372 160024 328736 160052
rect 324372 160012 324378 160024
rect 328730 160012 328736 160024
rect 328788 160012 328794 160064
rect 296254 158856 296260 158908
rect 296312 158896 296318 158908
rect 307662 158896 307668 158908
rect 296312 158868 307668 158896
rect 296312 158856 296318 158868
rect 307662 158856 307668 158868
rect 307720 158856 307726 158908
rect 275278 158788 275284 158840
rect 275336 158828 275342 158840
rect 307478 158828 307484 158840
rect 275336 158800 307484 158828
rect 275336 158788 275342 158800
rect 307478 158788 307484 158800
rect 307536 158788 307542 158840
rect 262950 158720 262956 158772
rect 263008 158760 263014 158772
rect 306926 158760 306932 158772
rect 263008 158732 306932 158760
rect 263008 158720 263014 158732
rect 306926 158720 306932 158732
rect 306984 158720 306990 158772
rect 252370 158652 252376 158704
rect 252428 158692 252434 158704
rect 276014 158692 276020 158704
rect 252428 158664 276020 158692
rect 252428 158652 252434 158664
rect 276014 158652 276020 158664
rect 276072 158652 276078 158704
rect 324406 158652 324412 158704
rect 324464 158692 324470 158704
rect 338298 158692 338304 158704
rect 324464 158664 338304 158692
rect 324464 158652 324470 158664
rect 338298 158652 338304 158664
rect 338356 158652 338362 158704
rect 252462 158584 252468 158636
rect 252520 158624 252526 158636
rect 265066 158624 265072 158636
rect 252520 158596 265072 158624
rect 252520 158584 252526 158596
rect 265066 158584 265072 158596
rect 265124 158584 265130 158636
rect 324314 158584 324320 158636
rect 324372 158624 324378 158636
rect 332870 158624 332876 158636
rect 324372 158596 332876 158624
rect 324372 158584 324378 158596
rect 332870 158584 332876 158596
rect 332928 158584 332934 158636
rect 293586 157496 293592 157548
rect 293644 157536 293650 157548
rect 307478 157536 307484 157548
rect 293644 157508 307484 157536
rect 293644 157496 293650 157508
rect 307478 157496 307484 157508
rect 307536 157496 307542 157548
rect 260098 157428 260104 157480
rect 260156 157468 260162 157480
rect 306926 157468 306932 157480
rect 260156 157440 306932 157468
rect 260156 157428 260162 157440
rect 306926 157428 306932 157440
rect 306984 157428 306990 157480
rect 253198 157360 253204 157412
rect 253256 157400 253262 157412
rect 307294 157400 307300 157412
rect 253256 157372 307300 157400
rect 253256 157360 253262 157372
rect 307294 157360 307300 157372
rect 307352 157360 307358 157412
rect 171778 157292 171784 157344
rect 171836 157332 171842 157344
rect 213914 157332 213920 157344
rect 171836 157304 213920 157332
rect 171836 157292 171842 157304
rect 213914 157292 213920 157304
rect 213972 157292 213978 157344
rect 252370 157292 252376 157344
rect 252428 157332 252434 157344
rect 267734 157332 267740 157344
rect 252428 157304 267740 157332
rect 252428 157292 252434 157304
rect 267734 157292 267740 157304
rect 267792 157292 267798 157344
rect 324314 157292 324320 157344
rect 324372 157332 324378 157344
rect 346394 157332 346400 157344
rect 324372 157304 346400 157332
rect 324372 157292 324378 157304
rect 346394 157292 346400 157304
rect 346452 157292 346458 157344
rect 210510 157224 210516 157276
rect 210568 157264 210574 157276
rect 214006 157264 214012 157276
rect 210568 157236 214012 157264
rect 210568 157224 210574 157236
rect 214006 157224 214012 157236
rect 214064 157224 214070 157276
rect 252462 157224 252468 157276
rect 252520 157264 252526 157276
rect 263594 157264 263600 157276
rect 252520 157236 263600 157264
rect 252520 157224 252526 157236
rect 263594 157224 263600 157236
rect 263652 157224 263658 157276
rect 324406 157224 324412 157276
rect 324464 157264 324470 157276
rect 343726 157264 343732 157276
rect 324464 157236 343732 157264
rect 324464 157224 324470 157236
rect 343726 157224 343732 157236
rect 343784 157224 343790 157276
rect 291930 156068 291936 156120
rect 291988 156108 291994 156120
rect 306742 156108 306748 156120
rect 291988 156080 306748 156108
rect 291988 156068 291994 156080
rect 306742 156068 306748 156080
rect 306800 156068 306806 156120
rect 275370 156000 275376 156052
rect 275428 156040 275434 156052
rect 307662 156040 307668 156052
rect 275428 156012 307668 156040
rect 275428 156000 275434 156012
rect 307662 156000 307668 156012
rect 307720 156000 307726 156052
rect 261478 155932 261484 155984
rect 261536 155972 261542 155984
rect 307570 155972 307576 155984
rect 261536 155944 307576 155972
rect 261536 155932 261542 155944
rect 307570 155932 307576 155944
rect 307628 155932 307634 155984
rect 170490 155864 170496 155916
rect 170548 155904 170554 155916
rect 213914 155904 213920 155916
rect 170548 155876 213920 155904
rect 170548 155864 170554 155876
rect 213914 155864 213920 155876
rect 213972 155864 213978 155916
rect 252370 155864 252376 155916
rect 252428 155904 252434 155916
rect 278774 155904 278780 155916
rect 252428 155876 278780 155904
rect 252428 155864 252434 155876
rect 278774 155864 278780 155876
rect 278832 155864 278838 155916
rect 324314 155864 324320 155916
rect 324372 155904 324378 155916
rect 347774 155904 347780 155916
rect 324372 155876 347780 155904
rect 324372 155864 324378 155876
rect 347774 155864 347780 155876
rect 347832 155864 347838 155916
rect 252462 155796 252468 155848
rect 252520 155836 252526 155848
rect 270586 155836 270592 155848
rect 252520 155808 270592 155836
rect 252520 155796 252526 155808
rect 270586 155796 270592 155808
rect 270644 155796 270650 155848
rect 298830 154708 298836 154760
rect 298888 154748 298894 154760
rect 307570 154748 307576 154760
rect 298888 154720 307576 154748
rect 298888 154708 298894 154720
rect 307570 154708 307576 154720
rect 307628 154708 307634 154760
rect 282362 154640 282368 154692
rect 282420 154680 282426 154692
rect 307662 154680 307668 154692
rect 282420 154652 307668 154680
rect 282420 154640 282426 154652
rect 307662 154640 307668 154652
rect 307720 154640 307726 154692
rect 262858 154572 262864 154624
rect 262916 154612 262922 154624
rect 307478 154612 307484 154624
rect 262916 154584 307484 154612
rect 262916 154572 262922 154584
rect 307478 154572 307484 154584
rect 307536 154572 307542 154624
rect 324314 154504 324320 154556
rect 324372 154544 324378 154556
rect 328638 154544 328644 154556
rect 324372 154516 328644 154544
rect 324372 154504 324378 154516
rect 328638 154504 328644 154516
rect 328696 154504 328702 154556
rect 252370 154436 252376 154488
rect 252428 154476 252434 154488
rect 269206 154476 269212 154488
rect 252428 154448 269212 154476
rect 252428 154436 252434 154448
rect 269206 154436 269212 154448
rect 269264 154436 269270 154488
rect 252462 154368 252468 154420
rect 252520 154408 252526 154420
rect 271966 154408 271972 154420
rect 252520 154380 271972 154408
rect 252520 154368 252526 154380
rect 271966 154368 271972 154380
rect 272024 154368 272030 154420
rect 251174 154096 251180 154148
rect 251232 154136 251238 154148
rect 253934 154136 253940 154148
rect 251232 154108 253940 154136
rect 251232 154096 251238 154108
rect 253934 154096 253940 154108
rect 253992 154096 253998 154148
rect 258902 153824 258908 153876
rect 258960 153864 258966 153876
rect 307386 153864 307392 153876
rect 258960 153836 307392 153864
rect 258960 153824 258966 153836
rect 307386 153824 307392 153836
rect 307444 153824 307450 153876
rect 301590 153280 301596 153332
rect 301648 153320 301654 153332
rect 307662 153320 307668 153332
rect 301648 153292 307668 153320
rect 301648 153280 301654 153292
rect 307662 153280 307668 153292
rect 307720 153280 307726 153332
rect 178678 153212 178684 153264
rect 178736 153252 178742 153264
rect 213914 153252 213920 153264
rect 178736 153224 213920 153252
rect 178736 153212 178742 153224
rect 213914 153212 213920 153224
rect 213972 153212 213978 153264
rect 254670 153212 254676 153264
rect 254728 153252 254734 153264
rect 307478 153252 307484 153264
rect 254728 153224 307484 153252
rect 254728 153212 254734 153224
rect 307478 153212 307484 153224
rect 307536 153212 307542 153264
rect 252462 153144 252468 153196
rect 252520 153184 252526 153196
rect 273254 153184 273260 153196
rect 252520 153156 273260 153184
rect 252520 153144 252526 153156
rect 273254 153144 273260 153156
rect 273312 153144 273318 153196
rect 324314 153144 324320 153196
rect 324372 153184 324378 153196
rect 347866 153184 347872 153196
rect 324372 153156 347872 153184
rect 324372 153144 324378 153156
rect 347866 153144 347872 153156
rect 347924 153144 347930 153196
rect 202138 151920 202144 151972
rect 202196 151960 202202 151972
rect 213914 151960 213920 151972
rect 202196 151932 213920 151960
rect 202196 151920 202202 151932
rect 213914 151920 213920 151932
rect 213972 151920 213978 151972
rect 301498 151920 301504 151972
rect 301556 151960 301562 151972
rect 307662 151960 307668 151972
rect 301556 151932 307668 151960
rect 301556 151920 301562 151932
rect 307662 151920 307668 151932
rect 307720 151920 307726 151972
rect 206278 151852 206284 151904
rect 206336 151892 206342 151904
rect 214006 151892 214012 151904
rect 206336 151864 214012 151892
rect 206336 151852 206342 151864
rect 214006 151852 214012 151864
rect 214064 151852 214070 151904
rect 257338 151852 257344 151904
rect 257396 151892 257402 151904
rect 307478 151892 307484 151904
rect 257396 151864 307484 151892
rect 257396 151852 257402 151864
rect 307478 151852 307484 151864
rect 307536 151852 307542 151904
rect 254762 151784 254768 151836
rect 254820 151824 254826 151836
rect 307662 151824 307668 151836
rect 254820 151796 307668 151824
rect 254820 151784 254826 151796
rect 307662 151784 307668 151796
rect 307720 151784 307726 151836
rect 252462 151716 252468 151768
rect 252520 151756 252526 151768
rect 262306 151756 262312 151768
rect 252520 151728 262312 151756
rect 252520 151716 252526 151728
rect 262306 151716 262312 151728
rect 262364 151716 262370 151768
rect 324314 151716 324320 151768
rect 324372 151756 324378 151768
rect 327350 151756 327356 151768
rect 324372 151728 327356 151756
rect 324372 151716 324378 151728
rect 327350 151716 327356 151728
rect 327408 151716 327414 151768
rect 251266 151444 251272 151496
rect 251324 151484 251330 151496
rect 254210 151484 254216 151496
rect 251324 151456 254216 151484
rect 251324 151444 251330 151456
rect 254210 151444 254216 151456
rect 254268 151444 254274 151496
rect 167638 151036 167644 151088
rect 167696 151076 167702 151088
rect 184842 151076 184848 151088
rect 167696 151048 184848 151076
rect 167696 151036 167702 151048
rect 184842 151036 184848 151048
rect 184900 151036 184906 151088
rect 289170 150560 289176 150612
rect 289228 150600 289234 150612
rect 307478 150600 307484 150612
rect 289228 150572 307484 150600
rect 289228 150560 289234 150572
rect 307478 150560 307484 150572
rect 307536 150560 307542 150612
rect 264422 150492 264428 150544
rect 264480 150532 264486 150544
rect 307662 150532 307668 150544
rect 264480 150504 307668 150532
rect 264480 150492 264486 150504
rect 307662 150492 307668 150504
rect 307720 150492 307726 150544
rect 178862 150424 178868 150476
rect 178920 150464 178926 150476
rect 214006 150464 214012 150476
rect 178920 150436 214012 150464
rect 178920 150424 178926 150436
rect 214006 150424 214012 150436
rect 214064 150424 214070 150476
rect 256142 150424 256148 150476
rect 256200 150464 256206 150476
rect 306926 150464 306932 150476
rect 256200 150436 306932 150464
rect 256200 150424 256206 150436
rect 306926 150424 306932 150436
rect 306984 150424 306990 150476
rect 169018 150356 169024 150408
rect 169076 150396 169082 150408
rect 213914 150396 213920 150408
rect 169076 150368 213920 150396
rect 169076 150356 169082 150368
rect 213914 150356 213920 150368
rect 213972 150356 213978 150408
rect 252278 150356 252284 150408
rect 252336 150396 252342 150408
rect 278866 150396 278872 150408
rect 252336 150368 278872 150396
rect 252336 150356 252342 150368
rect 278866 150356 278872 150368
rect 278924 150356 278930 150408
rect 324314 150356 324320 150408
rect 324372 150396 324378 150408
rect 346578 150396 346584 150408
rect 324372 150368 346584 150396
rect 324372 150356 324378 150368
rect 346578 150356 346584 150368
rect 346636 150356 346642 150408
rect 184842 150288 184848 150340
rect 184900 150328 184906 150340
rect 214006 150328 214012 150340
rect 184900 150300 214012 150328
rect 184900 150288 184906 150300
rect 214006 150288 214012 150300
rect 214064 150288 214070 150340
rect 324406 150288 324412 150340
rect 324464 150328 324470 150340
rect 346486 150328 346492 150340
rect 324464 150300 346492 150328
rect 324464 150288 324470 150300
rect 346486 150288 346492 150300
rect 346544 150288 346550 150340
rect 256050 149676 256056 149728
rect 256108 149716 256114 149728
rect 307018 149716 307024 149728
rect 256108 149688 307024 149716
rect 256108 149676 256114 149688
rect 307018 149676 307024 149688
rect 307076 149676 307082 149728
rect 251726 149268 251732 149320
rect 251784 149308 251790 149320
rect 256786 149308 256792 149320
rect 251784 149280 256792 149308
rect 251784 149268 251790 149280
rect 256786 149268 256792 149280
rect 256844 149268 256850 149320
rect 297634 149132 297640 149184
rect 297692 149172 297698 149184
rect 307662 149172 307668 149184
rect 297692 149144 307668 149172
rect 297692 149132 297698 149144
rect 307662 149132 307668 149144
rect 307720 149132 307726 149184
rect 282454 149064 282460 149116
rect 282512 149104 282518 149116
rect 306926 149104 306932 149116
rect 282512 149076 306932 149104
rect 282512 149064 282518 149076
rect 306926 149064 306932 149076
rect 306984 149064 306990 149116
rect 252462 148996 252468 149048
rect 252520 149036 252526 149048
rect 271874 149036 271880 149048
rect 252520 149008 271880 149036
rect 252520 148996 252526 149008
rect 271874 148996 271880 149008
rect 271932 148996 271938 149048
rect 324314 148996 324320 149048
rect 324372 149036 324378 149048
rect 345106 149036 345112 149048
rect 324372 149008 345112 149036
rect 324372 148996 324378 149008
rect 345106 148996 345112 149008
rect 345164 148996 345170 149048
rect 324406 148928 324412 148980
rect 324464 148968 324470 148980
rect 337010 148968 337016 148980
rect 324464 148940 337016 148968
rect 324464 148928 324470 148940
rect 337010 148928 337016 148940
rect 337068 148928 337074 148980
rect 251266 148860 251272 148912
rect 251324 148900 251330 148912
rect 254118 148900 254124 148912
rect 251324 148872 254124 148900
rect 251324 148860 251330 148872
rect 254118 148860 254124 148872
rect 254176 148860 254182 148912
rect 251910 148724 251916 148776
rect 251968 148764 251974 148776
rect 255498 148764 255504 148776
rect 251968 148736 255504 148764
rect 251968 148724 251974 148736
rect 255498 148724 255504 148736
rect 255556 148724 255562 148776
rect 303062 147772 303068 147824
rect 303120 147812 303126 147824
rect 307570 147812 307576 147824
rect 303120 147784 307576 147812
rect 303120 147772 303126 147784
rect 307570 147772 307576 147784
rect 307628 147772 307634 147824
rect 280890 147704 280896 147756
rect 280948 147744 280954 147756
rect 307662 147744 307668 147756
rect 280948 147716 307668 147744
rect 280948 147704 280954 147716
rect 307662 147704 307668 147716
rect 307720 147704 307726 147756
rect 170398 147636 170404 147688
rect 170456 147676 170462 147688
rect 213914 147676 213920 147688
rect 170456 147648 213920 147676
rect 170456 147636 170462 147648
rect 213914 147636 213920 147648
rect 213972 147636 213978 147688
rect 257522 147636 257528 147688
rect 257580 147676 257586 147688
rect 306926 147676 306932 147688
rect 257580 147648 306932 147676
rect 257580 147636 257586 147648
rect 306926 147636 306932 147648
rect 306984 147636 306990 147688
rect 252462 147568 252468 147620
rect 252520 147608 252526 147620
rect 281534 147608 281540 147620
rect 252520 147580 281540 147608
rect 252520 147568 252526 147580
rect 281534 147568 281540 147580
rect 281592 147568 281598 147620
rect 324314 147568 324320 147620
rect 324372 147608 324378 147620
rect 340874 147608 340880 147620
rect 324372 147580 340880 147608
rect 324372 147568 324378 147580
rect 340874 147568 340880 147580
rect 340932 147568 340938 147620
rect 251726 147500 251732 147552
rect 251784 147540 251790 147552
rect 274726 147540 274732 147552
rect 251784 147512 274732 147540
rect 251784 147500 251790 147512
rect 274726 147500 274732 147512
rect 274784 147500 274790 147552
rect 287974 146888 287980 146940
rect 288032 146928 288038 146940
rect 307110 146928 307116 146940
rect 288032 146900 307116 146928
rect 288032 146888 288038 146900
rect 307110 146888 307116 146900
rect 307168 146888 307174 146940
rect 251726 146820 251732 146872
rect 251784 146860 251790 146872
rect 255590 146860 255596 146872
rect 251784 146832 255596 146860
rect 251784 146820 251790 146832
rect 255590 146820 255596 146832
rect 255648 146820 255654 146872
rect 181438 146344 181444 146396
rect 181496 146384 181502 146396
rect 213914 146384 213920 146396
rect 181496 146356 213920 146384
rect 181496 146344 181502 146356
rect 213914 146344 213920 146356
rect 213972 146344 213978 146396
rect 274082 146344 274088 146396
rect 274140 146384 274146 146396
rect 307662 146384 307668 146396
rect 274140 146356 307668 146384
rect 274140 146344 274146 146356
rect 307662 146344 307668 146356
rect 307720 146344 307726 146396
rect 170490 146276 170496 146328
rect 170548 146316 170554 146328
rect 214006 146316 214012 146328
rect 170548 146288 214012 146316
rect 170548 146276 170554 146288
rect 214006 146276 214012 146288
rect 214064 146276 214070 146328
rect 256234 146276 256240 146328
rect 256292 146316 256298 146328
rect 306742 146316 306748 146328
rect 256292 146288 306748 146316
rect 256292 146276 256298 146288
rect 306742 146276 306748 146288
rect 306800 146276 306806 146328
rect 251910 146208 251916 146260
rect 251968 146248 251974 146260
rect 273346 146248 273352 146260
rect 251968 146220 273352 146248
rect 251968 146208 251974 146220
rect 273346 146208 273352 146220
rect 273404 146208 273410 146260
rect 324406 146208 324412 146260
rect 324464 146248 324470 146260
rect 338206 146248 338212 146260
rect 324464 146220 338212 146248
rect 324464 146208 324470 146220
rect 338206 146208 338212 146220
rect 338264 146208 338270 146260
rect 251726 146140 251732 146192
rect 251784 146180 251790 146192
rect 266538 146180 266544 146192
rect 251784 146152 266544 146180
rect 251784 146140 251790 146152
rect 266538 146140 266544 146152
rect 266596 146140 266602 146192
rect 324314 146140 324320 146192
rect 324372 146180 324378 146192
rect 334158 146180 334164 146192
rect 324372 146152 334164 146180
rect 324372 146140 324378 146152
rect 334158 146140 334164 146152
rect 334216 146140 334222 146192
rect 252094 146072 252100 146124
rect 252152 146112 252158 146124
rect 263686 146112 263692 146124
rect 252152 146084 263692 146112
rect 252152 146072 252158 146084
rect 263686 146072 263692 146084
rect 263744 146072 263750 146124
rect 300486 146072 300492 146124
rect 300544 146112 300550 146124
rect 306650 146112 306656 146124
rect 300544 146084 306656 146112
rect 300544 146072 300550 146084
rect 306650 146072 306656 146084
rect 306708 146072 306714 146124
rect 176010 144984 176016 145036
rect 176068 145024 176074 145036
rect 214006 145024 214012 145036
rect 176068 144996 214012 145024
rect 176068 144984 176074 144996
rect 214006 144984 214012 144996
rect 214064 144984 214070 145036
rect 267090 144984 267096 145036
rect 267148 145024 267154 145036
rect 307662 145024 307668 145036
rect 267148 144996 307668 145024
rect 267148 144984 267154 144996
rect 307662 144984 307668 144996
rect 307720 144984 307726 145036
rect 173158 144916 173164 144968
rect 173216 144956 173222 144968
rect 213914 144956 213920 144968
rect 173216 144928 213920 144956
rect 173216 144916 173222 144928
rect 213914 144916 213920 144928
rect 213972 144916 213978 144968
rect 253474 144916 253480 144968
rect 253532 144956 253538 144968
rect 307570 144956 307576 144968
rect 253532 144928 307576 144956
rect 253532 144916 253538 144928
rect 307570 144916 307576 144928
rect 307628 144916 307634 144968
rect 252370 144848 252376 144900
rect 252428 144888 252434 144900
rect 270494 144888 270500 144900
rect 252428 144860 270500 144888
rect 252428 144848 252434 144860
rect 270494 144848 270500 144860
rect 270552 144848 270558 144900
rect 324314 144848 324320 144900
rect 324372 144888 324378 144900
rect 342530 144888 342536 144900
rect 324372 144860 342536 144888
rect 324372 144848 324378 144860
rect 342530 144848 342536 144860
rect 342588 144848 342594 144900
rect 252462 144780 252468 144832
rect 252520 144820 252526 144832
rect 267826 144820 267832 144832
rect 252520 144792 267832 144820
rect 252520 144780 252526 144792
rect 267826 144780 267832 144792
rect 267884 144780 267890 144832
rect 324406 144780 324412 144832
rect 324464 144820 324470 144832
rect 331214 144820 331220 144832
rect 324464 144792 331220 144820
rect 324464 144780 324470 144792
rect 331214 144780 331220 144792
rect 331272 144780 331278 144832
rect 252094 144168 252100 144220
rect 252152 144208 252158 144220
rect 264238 144208 264244 144220
rect 252152 144180 264244 144208
rect 252152 144168 252158 144180
rect 264238 144168 264244 144180
rect 264296 144168 264302 144220
rect 279694 144168 279700 144220
rect 279752 144208 279758 144220
rect 307386 144208 307392 144220
rect 279752 144180 307392 144208
rect 279752 144168 279758 144180
rect 307386 144168 307392 144180
rect 307444 144168 307450 144220
rect 252462 144032 252468 144084
rect 252520 144072 252526 144084
rect 259730 144072 259736 144084
rect 252520 144044 259736 144072
rect 252520 144032 252526 144044
rect 259730 144032 259736 144044
rect 259788 144032 259794 144084
rect 210418 143624 210424 143676
rect 210476 143664 210482 143676
rect 214006 143664 214012 143676
rect 210476 143636 214012 143664
rect 210476 143624 210482 143636
rect 214006 143624 214012 143636
rect 214064 143624 214070 143676
rect 174538 143556 174544 143608
rect 174596 143596 174602 143608
rect 213914 143596 213920 143608
rect 174596 143568 213920 143596
rect 174596 143556 174602 143568
rect 213914 143556 213920 143568
rect 213972 143556 213978 143608
rect 286410 143556 286416 143608
rect 286468 143596 286474 143608
rect 307662 143596 307668 143608
rect 286468 143568 307668 143596
rect 286468 143556 286474 143568
rect 307662 143556 307668 143568
rect 307720 143556 307726 143608
rect 252462 143488 252468 143540
rect 252520 143528 252526 143540
rect 269114 143528 269120 143540
rect 252520 143500 269120 143528
rect 252520 143488 252526 143500
rect 269114 143488 269120 143500
rect 269172 143488 269178 143540
rect 251910 142808 251916 142860
rect 251968 142848 251974 142860
rect 293218 142848 293224 142860
rect 251968 142820 293224 142848
rect 251968 142808 251974 142820
rect 293218 142808 293224 142820
rect 293276 142808 293282 142860
rect 324314 142672 324320 142724
rect 324372 142712 324378 142724
rect 327074 142712 327080 142724
rect 324372 142684 327080 142712
rect 324372 142672 324378 142684
rect 327074 142672 327080 142684
rect 327132 142672 327138 142724
rect 171778 142196 171784 142248
rect 171836 142236 171842 142248
rect 213914 142236 213920 142248
rect 171836 142208 213920 142236
rect 171836 142196 171842 142208
rect 213914 142196 213920 142208
rect 213972 142196 213978 142248
rect 286318 142196 286324 142248
rect 286376 142236 286382 142248
rect 307662 142236 307668 142248
rect 286376 142208 307668 142236
rect 286376 142196 286382 142208
rect 307662 142196 307668 142208
rect 307720 142196 307726 142248
rect 169018 142128 169024 142180
rect 169076 142168 169082 142180
rect 214006 142168 214012 142180
rect 169076 142140 214012 142168
rect 169076 142128 169082 142140
rect 214006 142128 214012 142140
rect 214064 142128 214070 142180
rect 257430 142128 257436 142180
rect 257488 142168 257494 142180
rect 306742 142168 306748 142180
rect 257488 142140 306748 142168
rect 257488 142128 257494 142140
rect 306742 142128 306748 142140
rect 306800 142128 306806 142180
rect 252462 142060 252468 142112
rect 252520 142100 252526 142112
rect 258350 142100 258356 142112
rect 252520 142072 258356 142100
rect 252520 142060 252526 142072
rect 258350 142060 258356 142072
rect 258408 142060 258414 142112
rect 324314 142060 324320 142112
rect 324372 142100 324378 142112
rect 349154 142100 349160 142112
rect 324372 142072 349160 142100
rect 324372 142060 324378 142072
rect 349154 142060 349160 142072
rect 349212 142060 349218 142112
rect 324498 141992 324504 142044
rect 324556 142032 324562 142044
rect 333974 142032 333980 142044
rect 324556 142004 333980 142032
rect 324556 141992 324562 142004
rect 333974 141992 333980 142004
rect 334032 141992 334038 142044
rect 323670 141652 323676 141704
rect 323728 141692 323734 141704
rect 324406 141692 324412 141704
rect 323728 141664 324412 141692
rect 323728 141652 323734 141664
rect 324406 141652 324412 141664
rect 324464 141652 324470 141704
rect 251818 141380 251824 141432
rect 251876 141420 251882 141432
rect 275278 141420 275284 141432
rect 251876 141392 275284 141420
rect 251876 141380 251882 141392
rect 275278 141380 275284 141392
rect 275336 141380 275342 141432
rect 276750 141380 276756 141432
rect 276808 141420 276814 141432
rect 307202 141420 307208 141432
rect 276808 141392 307208 141420
rect 276808 141380 276814 141392
rect 307202 141380 307208 141392
rect 307260 141380 307266 141432
rect 305914 140836 305920 140888
rect 305972 140876 305978 140888
rect 307478 140876 307484 140888
rect 305972 140848 307484 140876
rect 305972 140836 305978 140848
rect 307478 140836 307484 140848
rect 307536 140836 307542 140888
rect 193858 140768 193864 140820
rect 193916 140808 193922 140820
rect 213914 140808 213920 140820
rect 193916 140780 213920 140808
rect 193916 140768 193922 140780
rect 213914 140768 213920 140780
rect 213972 140768 213978 140820
rect 254578 140768 254584 140820
rect 254636 140808 254642 140820
rect 307662 140808 307668 140820
rect 254636 140780 307668 140808
rect 254636 140768 254642 140780
rect 307662 140768 307668 140780
rect 307720 140768 307726 140820
rect 253382 140020 253388 140072
rect 253440 140060 253446 140072
rect 306558 140060 306564 140072
rect 253440 140032 306564 140060
rect 253440 140020 253446 140032
rect 306558 140020 306564 140032
rect 306616 140020 306622 140072
rect 251358 139884 251364 139936
rect 251416 139924 251422 139936
rect 256694 139924 256700 139936
rect 251416 139896 256700 139924
rect 251416 139884 251422 139896
rect 256694 139884 256700 139896
rect 256752 139884 256758 139936
rect 304442 139544 304448 139596
rect 304500 139584 304506 139596
rect 307386 139584 307392 139596
rect 304500 139556 307392 139584
rect 304500 139544 304506 139556
rect 307386 139544 307392 139556
rect 307444 139544 307450 139596
rect 289078 139476 289084 139528
rect 289136 139516 289142 139528
rect 307570 139516 307576 139528
rect 289136 139488 307576 139516
rect 289136 139476 289142 139488
rect 307570 139476 307576 139488
rect 307628 139476 307634 139528
rect 166258 139408 166264 139460
rect 166316 139448 166322 139460
rect 213914 139448 213920 139460
rect 166316 139420 213920 139448
rect 166316 139408 166322 139420
rect 213914 139408 213920 139420
rect 213972 139408 213978 139460
rect 280798 139408 280804 139460
rect 280856 139448 280862 139460
rect 307662 139448 307668 139460
rect 280856 139420 307668 139448
rect 280856 139408 280862 139420
rect 307662 139408 307668 139420
rect 307720 139408 307726 139460
rect 252462 139340 252468 139392
rect 252520 139380 252526 139392
rect 280154 139380 280160 139392
rect 252520 139352 280160 139380
rect 252520 139340 252526 139352
rect 280154 139340 280160 139352
rect 280212 139340 280218 139392
rect 324314 139340 324320 139392
rect 324372 139380 324378 139392
rect 350534 139380 350540 139392
rect 324372 139352 350540 139380
rect 324372 139340 324378 139352
rect 350534 139340 350540 139352
rect 350592 139340 350598 139392
rect 324498 139272 324504 139324
rect 324556 139312 324562 139324
rect 332778 139312 332784 139324
rect 324556 139284 332784 139312
rect 324556 139272 324562 139284
rect 332778 139272 332784 139284
rect 332836 139272 332842 139324
rect 324958 139204 324964 139256
rect 325016 139244 325022 139256
rect 327166 139244 327172 139256
rect 325016 139216 327172 139244
rect 325016 139204 325022 139216
rect 327166 139204 327172 139216
rect 327224 139204 327230 139256
rect 251542 138660 251548 138712
rect 251600 138700 251606 138712
rect 278222 138700 278228 138712
rect 251600 138672 278228 138700
rect 251600 138660 251606 138672
rect 278222 138660 278228 138672
rect 278280 138660 278286 138712
rect 298738 138116 298744 138168
rect 298796 138156 298802 138168
rect 307662 138156 307668 138168
rect 298796 138128 307668 138156
rect 298796 138116 298802 138128
rect 307662 138116 307668 138128
rect 307720 138116 307726 138168
rect 278130 138048 278136 138100
rect 278188 138088 278194 138100
rect 307570 138088 307576 138100
rect 278188 138060 307576 138088
rect 278188 138048 278194 138060
rect 307570 138048 307576 138060
rect 307628 138048 307634 138100
rect 171870 137980 171876 138032
rect 171928 138020 171934 138032
rect 213914 138020 213920 138032
rect 171928 137992 213920 138020
rect 171928 137980 171934 137992
rect 213914 137980 213920 137992
rect 213972 137980 213978 138032
rect 273898 137980 273904 138032
rect 273956 138020 273962 138032
rect 307478 138020 307484 138032
rect 273956 137992 307484 138020
rect 273956 137980 273962 137992
rect 307478 137980 307484 137992
rect 307536 137980 307542 138032
rect 252462 137912 252468 137964
rect 252520 137952 252526 137964
rect 277394 137952 277400 137964
rect 252520 137924 277400 137952
rect 252520 137912 252526 137924
rect 277394 137912 277400 137924
rect 277452 137912 277458 137964
rect 324314 137912 324320 137964
rect 324372 137952 324378 137964
rect 342438 137952 342444 137964
rect 324372 137924 342444 137952
rect 324372 137912 324378 137924
rect 342438 137912 342444 137924
rect 342496 137912 342502 137964
rect 251358 137844 251364 137896
rect 251416 137884 251422 137896
rect 274634 137884 274640 137896
rect 251416 137856 274640 137884
rect 251416 137844 251422 137856
rect 274634 137844 274640 137856
rect 274692 137844 274698 137896
rect 324498 137844 324504 137896
rect 324556 137884 324562 137896
rect 330018 137884 330024 137896
rect 324556 137856 330024 137884
rect 324556 137844 324562 137856
rect 330018 137844 330024 137856
rect 330076 137844 330082 137896
rect 174814 137232 174820 137284
rect 174872 137272 174878 137284
rect 214558 137272 214564 137284
rect 174872 137244 214564 137272
rect 174872 137232 174878 137244
rect 214558 137232 214564 137244
rect 214616 137232 214622 137284
rect 253290 137232 253296 137284
rect 253348 137272 253354 137284
rect 307294 137272 307300 137284
rect 253348 137244 307300 137272
rect 253348 137232 253354 137244
rect 307294 137232 307300 137244
rect 307352 137232 307358 137284
rect 282270 136688 282276 136740
rect 282328 136728 282334 136740
rect 307478 136728 307484 136740
rect 282328 136700 307484 136728
rect 282328 136688 282334 136700
rect 307478 136688 307484 136700
rect 307536 136688 307542 136740
rect 203518 136620 203524 136672
rect 203576 136660 203582 136672
rect 213914 136660 213920 136672
rect 203576 136632 213920 136660
rect 203576 136620 203582 136632
rect 213914 136620 213920 136632
rect 213972 136620 213978 136672
rect 264238 136620 264244 136672
rect 264296 136660 264302 136672
rect 306926 136660 306932 136672
rect 264296 136632 306932 136660
rect 264296 136620 264302 136632
rect 306926 136620 306932 136632
rect 306984 136620 306990 136672
rect 252462 136552 252468 136604
rect 252520 136592 252526 136604
rect 291838 136592 291844 136604
rect 252520 136564 291844 136592
rect 252520 136552 252526 136564
rect 291838 136552 291844 136564
rect 291896 136552 291902 136604
rect 324498 136552 324504 136604
rect 324556 136592 324562 136604
rect 343634 136592 343640 136604
rect 324556 136564 343640 136592
rect 324556 136552 324562 136564
rect 343634 136552 343640 136564
rect 343692 136552 343698 136604
rect 252370 136484 252376 136536
rect 252428 136524 252434 136536
rect 266998 136524 267004 136536
rect 252428 136496 267004 136524
rect 252428 136484 252434 136496
rect 266998 136484 267004 136496
rect 267056 136484 267062 136536
rect 324314 136484 324320 136536
rect 324372 136524 324378 136536
rect 339678 136524 339684 136536
rect 324372 136496 339684 136524
rect 324372 136484 324378 136496
rect 339678 136484 339684 136496
rect 339736 136484 339742 136536
rect 302878 135464 302884 135516
rect 302936 135504 302942 135516
rect 307570 135504 307576 135516
rect 302936 135476 307576 135504
rect 302936 135464 302942 135476
rect 307570 135464 307576 135476
rect 307628 135464 307634 135516
rect 297358 135396 297364 135448
rect 297416 135436 297422 135448
rect 307662 135436 307668 135448
rect 297416 135408 307668 135436
rect 297416 135396 297422 135408
rect 307662 135396 307668 135408
rect 307720 135396 307726 135448
rect 207750 135328 207756 135380
rect 207808 135368 207814 135380
rect 214006 135368 214012 135380
rect 207808 135340 214012 135368
rect 207808 135328 207814 135340
rect 214006 135328 214012 135340
rect 214064 135328 214070 135380
rect 284938 135328 284944 135380
rect 284996 135368 285002 135380
rect 307386 135368 307392 135380
rect 284996 135340 307392 135368
rect 284996 135328 285002 135340
rect 307386 135328 307392 135340
rect 307444 135328 307450 135380
rect 174630 135260 174636 135312
rect 174688 135300 174694 135312
rect 213914 135300 213920 135312
rect 174688 135272 213920 135300
rect 174688 135260 174694 135272
rect 213914 135260 213920 135272
rect 213972 135260 213978 135312
rect 271230 135260 271236 135312
rect 271288 135300 271294 135312
rect 307478 135300 307484 135312
rect 271288 135272 307484 135300
rect 271288 135260 271294 135272
rect 307478 135260 307484 135272
rect 307536 135260 307542 135312
rect 251634 135192 251640 135244
rect 251692 135232 251698 135244
rect 273990 135232 273996 135244
rect 251692 135204 273996 135232
rect 251692 135192 251698 135204
rect 273990 135192 273996 135204
rect 274048 135192 274054 135244
rect 252462 134580 252468 134632
rect 252520 134620 252526 134632
rect 260282 134620 260288 134632
rect 252520 134592 260288 134620
rect 252520 134580 252526 134592
rect 260282 134580 260288 134592
rect 260340 134580 260346 134632
rect 251542 134512 251548 134564
rect 251600 134552 251606 134564
rect 283650 134552 283656 134564
rect 251600 134524 283656 134552
rect 251600 134512 251606 134524
rect 283650 134512 283656 134524
rect 283708 134512 283714 134564
rect 290642 134036 290648 134088
rect 290700 134076 290706 134088
rect 307662 134076 307668 134088
rect 290700 134048 307668 134076
rect 290700 134036 290706 134048
rect 307662 134036 307668 134048
rect 307720 134036 307726 134088
rect 192478 133968 192484 134020
rect 192536 134008 192542 134020
rect 213914 134008 213920 134020
rect 192536 133980 213920 134008
rect 192536 133968 192542 133980
rect 213914 133968 213920 133980
rect 213972 133968 213978 134020
rect 283742 133968 283748 134020
rect 283800 134008 283806 134020
rect 307570 134008 307576 134020
rect 283800 133980 307576 134008
rect 283800 133968 283806 133980
rect 307570 133968 307576 133980
rect 307628 133968 307634 134020
rect 169110 133900 169116 133952
rect 169168 133940 169174 133952
rect 214006 133940 214012 133952
rect 169168 133912 214012 133940
rect 169168 133900 169174 133912
rect 214006 133900 214012 133912
rect 214064 133900 214070 133952
rect 275278 133900 275284 133952
rect 275336 133940 275342 133952
rect 306742 133940 306748 133952
rect 275336 133912 306748 133940
rect 275336 133900 275342 133912
rect 306742 133900 306748 133912
rect 306800 133900 306806 133952
rect 251450 133832 251456 133884
rect 251508 133872 251514 133884
rect 289262 133872 289268 133884
rect 251508 133844 289268 133872
rect 251508 133832 251514 133844
rect 289262 133832 289268 133844
rect 289320 133832 289326 133884
rect 324314 133832 324320 133884
rect 324372 133872 324378 133884
rect 328546 133872 328552 133884
rect 324372 133844 328552 133872
rect 324372 133832 324378 133844
rect 328546 133832 328552 133844
rect 328604 133832 328610 133884
rect 252462 133764 252468 133816
rect 252520 133804 252526 133816
rect 264330 133804 264336 133816
rect 252520 133776 264336 133804
rect 252520 133764 252526 133776
rect 264330 133764 264336 133776
rect 264388 133764 264394 133816
rect 176102 133152 176108 133204
rect 176160 133192 176166 133204
rect 214098 133192 214104 133204
rect 176160 133164 214104 133192
rect 176160 133152 176166 133164
rect 214098 133152 214104 133164
rect 214156 133152 214162 133204
rect 211890 132880 211896 132932
rect 211948 132920 211954 132932
rect 213914 132920 213920 132932
rect 211948 132892 213920 132920
rect 211948 132880 211954 132892
rect 213914 132880 213920 132892
rect 213972 132880 213978 132932
rect 293218 132540 293224 132592
rect 293276 132580 293282 132592
rect 307662 132580 307668 132592
rect 293276 132552 307668 132580
rect 293276 132540 293282 132552
rect 307662 132540 307668 132552
rect 307720 132540 307726 132592
rect 287698 132472 287704 132524
rect 287756 132512 287762 132524
rect 307478 132512 307484 132524
rect 287756 132484 307484 132512
rect 287756 132472 287762 132484
rect 307478 132472 307484 132484
rect 307536 132472 307542 132524
rect 252278 132404 252284 132456
rect 252336 132444 252342 132456
rect 287882 132444 287888 132456
rect 252336 132416 287888 132444
rect 252336 132404 252342 132416
rect 287882 132404 287888 132416
rect 287940 132404 287946 132456
rect 324498 132404 324504 132456
rect 324556 132444 324562 132456
rect 345014 132444 345020 132456
rect 324556 132416 345020 132444
rect 324556 132404 324562 132416
rect 345014 132404 345020 132416
rect 345072 132404 345078 132456
rect 252002 132336 252008 132388
rect 252060 132376 252066 132388
rect 271322 132376 271328 132388
rect 252060 132348 271328 132376
rect 252060 132336 252066 132348
rect 271322 132336 271328 132348
rect 271380 132336 271386 132388
rect 324314 132336 324320 132388
rect 324372 132376 324378 132388
rect 341150 132376 341156 132388
rect 324372 132348 341156 132376
rect 324372 132336 324378 132348
rect 341150 132336 341156 132348
rect 341208 132336 341214 132388
rect 251358 132268 251364 132320
rect 251416 132308 251422 132320
rect 261754 132308 261760 132320
rect 251416 132280 261760 132308
rect 251416 132268 251422 132280
rect 261754 132268 261760 132280
rect 261812 132268 261818 132320
rect 291838 131248 291844 131300
rect 291896 131288 291902 131300
rect 306742 131288 306748 131300
rect 291896 131260 306748 131288
rect 291896 131248 291902 131260
rect 306742 131248 306748 131260
rect 306800 131248 306806 131300
rect 287790 131180 287796 131232
rect 287848 131220 287854 131232
rect 307662 131220 307668 131232
rect 287848 131192 307668 131220
rect 287848 131180 287854 131192
rect 307662 131180 307668 131192
rect 307720 131180 307726 131232
rect 180150 131112 180156 131164
rect 180208 131152 180214 131164
rect 213914 131152 213920 131164
rect 180208 131124 213920 131152
rect 180208 131112 180214 131124
rect 213914 131112 213920 131124
rect 213972 131112 213978 131164
rect 279510 131112 279516 131164
rect 279568 131152 279574 131164
rect 307478 131152 307484 131164
rect 279568 131124 307484 131152
rect 279568 131112 279574 131124
rect 307478 131112 307484 131124
rect 307536 131112 307542 131164
rect 251726 131044 251732 131096
rect 251784 131084 251790 131096
rect 285030 131084 285036 131096
rect 251784 131056 285036 131084
rect 251784 131044 251790 131056
rect 285030 131044 285036 131056
rect 285088 131044 285094 131096
rect 324314 131044 324320 131096
rect 324372 131084 324378 131096
rect 331306 131084 331312 131096
rect 324372 131056 331312 131084
rect 324372 131044 324378 131056
rect 331306 131044 331312 131056
rect 331364 131044 331370 131096
rect 252002 130976 252008 131028
rect 252060 131016 252066 131028
rect 279602 131016 279608 131028
rect 252060 130988 279608 131016
rect 252060 130976 252066 130988
rect 279602 130976 279608 130988
rect 279660 130976 279666 131028
rect 324406 130976 324412 131028
rect 324464 131016 324470 131028
rect 331398 131016 331404 131028
rect 324464 130988 331404 131016
rect 324464 130976 324470 130988
rect 331398 130976 331404 130988
rect 331456 130976 331462 131028
rect 252462 129888 252468 129940
rect 252520 129928 252526 129940
rect 258810 129928 258816 129940
rect 252520 129900 258816 129928
rect 252520 129888 252526 129900
rect 258810 129888 258816 129900
rect 258868 129888 258874 129940
rect 290550 129888 290556 129940
rect 290608 129928 290614 129940
rect 306742 129928 306748 129940
rect 290608 129900 306748 129928
rect 290608 129888 290614 129900
rect 306742 129888 306748 129900
rect 306800 129888 306806 129940
rect 279418 129820 279424 129872
rect 279476 129860 279482 129872
rect 306926 129860 306932 129872
rect 279476 129832 306932 129860
rect 279476 129820 279482 129832
rect 306926 129820 306932 129832
rect 306984 129820 306990 129872
rect 189718 129752 189724 129804
rect 189776 129792 189782 129804
rect 213914 129792 213920 129804
rect 189776 129764 213920 129792
rect 189776 129752 189782 129764
rect 213914 129752 213920 129764
rect 213972 129752 213978 129804
rect 276658 129752 276664 129804
rect 276716 129792 276722 129804
rect 307662 129792 307668 129804
rect 276716 129764 307668 129792
rect 276716 129752 276722 129764
rect 307662 129752 307668 129764
rect 307720 129752 307726 129804
rect 251726 129684 251732 129736
rect 251784 129724 251790 129736
rect 283558 129724 283564 129736
rect 251784 129696 283564 129724
rect 251784 129684 251790 129696
rect 283558 129684 283564 129696
rect 283616 129684 283622 129736
rect 324314 129684 324320 129736
rect 324372 129724 324378 129736
rect 330110 129724 330116 129736
rect 324372 129696 330116 129724
rect 324372 129684 324378 129696
rect 330110 129684 330116 129696
rect 330168 129684 330174 129736
rect 252094 129616 252100 129668
rect 252152 129656 252158 129668
rect 272518 129656 272524 129668
rect 252152 129628 272524 129656
rect 252152 129616 252158 129628
rect 272518 129616 272524 129628
rect 272576 129616 272582 129668
rect 294598 128460 294604 128512
rect 294656 128500 294662 128512
rect 307662 128500 307668 128512
rect 294656 128472 307668 128500
rect 294656 128460 294662 128472
rect 307662 128460 307668 128472
rect 307720 128460 307726 128512
rect 197998 128392 198004 128444
rect 198056 128432 198062 128444
rect 214006 128432 214012 128444
rect 198056 128404 214012 128432
rect 198056 128392 198062 128404
rect 214006 128392 214012 128404
rect 214064 128392 214070 128444
rect 273990 128392 273996 128444
rect 274048 128432 274054 128444
rect 307570 128432 307576 128444
rect 274048 128404 307576 128432
rect 274048 128392 274054 128404
rect 307570 128392 307576 128404
rect 307628 128392 307634 128444
rect 173250 128324 173256 128376
rect 173308 128364 173314 128376
rect 213914 128364 213920 128376
rect 173308 128336 213920 128364
rect 173308 128324 173314 128336
rect 213914 128324 213920 128336
rect 213972 128324 213978 128376
rect 265618 128324 265624 128376
rect 265676 128364 265682 128376
rect 307478 128364 307484 128376
rect 265676 128336 307484 128364
rect 265676 128324 265682 128336
rect 307478 128324 307484 128336
rect 307536 128324 307542 128376
rect 252002 128256 252008 128308
rect 252060 128296 252066 128308
rect 271138 128296 271144 128308
rect 252060 128268 271144 128296
rect 252060 128256 252066 128268
rect 271138 128256 271144 128268
rect 271196 128256 271202 128308
rect 324314 128256 324320 128308
rect 324372 128296 324378 128308
rect 329926 128296 329932 128308
rect 324372 128268 329932 128296
rect 324372 128256 324378 128268
rect 329926 128256 329932 128268
rect 329984 128256 329990 128308
rect 252462 128188 252468 128240
rect 252520 128228 252526 128240
rect 265894 128228 265900 128240
rect 252520 128200 265900 128228
rect 252520 128188 252526 128200
rect 265894 128188 265900 128200
rect 265952 128188 265958 128240
rect 295978 127100 295984 127152
rect 296036 127140 296042 127152
rect 307662 127140 307668 127152
rect 296036 127112 307668 127140
rect 296036 127100 296042 127112
rect 307662 127100 307668 127112
rect 307720 127100 307726 127152
rect 178770 127032 178776 127084
rect 178828 127072 178834 127084
rect 213914 127072 213920 127084
rect 178828 127044 213920 127072
rect 178828 127032 178834 127044
rect 213914 127032 213920 127044
rect 213972 127032 213978 127084
rect 285030 127032 285036 127084
rect 285088 127072 285094 127084
rect 307570 127072 307576 127084
rect 285088 127044 307576 127072
rect 285088 127032 285094 127044
rect 307570 127032 307576 127044
rect 307628 127032 307634 127084
rect 177298 126964 177304 127016
rect 177356 127004 177362 127016
rect 214006 127004 214012 127016
rect 177356 126976 214012 127004
rect 177356 126964 177362 126976
rect 214006 126964 214012 126976
rect 214064 126964 214070 127016
rect 272518 126964 272524 127016
rect 272576 127004 272582 127016
rect 307478 127004 307484 127016
rect 272576 126976 307484 127004
rect 272576 126964 272582 126976
rect 307478 126964 307484 126976
rect 307536 126964 307542 127016
rect 252094 126896 252100 126948
rect 252152 126936 252158 126948
rect 269850 126936 269856 126948
rect 252152 126908 269856 126936
rect 252152 126896 252158 126908
rect 269850 126896 269856 126908
rect 269908 126896 269914 126948
rect 324314 126896 324320 126948
rect 324372 126936 324378 126948
rect 328454 126936 328460 126948
rect 324372 126908 328460 126936
rect 324372 126896 324378 126908
rect 328454 126896 328460 126908
rect 328512 126896 328518 126948
rect 392578 126896 392584 126948
rect 392636 126936 392642 126948
rect 580166 126936 580172 126948
rect 392636 126908 580172 126936
rect 392636 126896 392642 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 252462 126828 252468 126880
rect 252520 126868 252526 126880
rect 261662 126868 261668 126880
rect 252520 126840 261668 126868
rect 252520 126828 252526 126840
rect 261662 126828 261668 126840
rect 261720 126828 261726 126880
rect 251266 126216 251272 126268
rect 251324 126256 251330 126268
rect 294782 126256 294788 126268
rect 251324 126228 294788 126256
rect 251324 126216 251330 126228
rect 294782 126216 294788 126228
rect 294840 126216 294846 126268
rect 294690 125740 294696 125792
rect 294748 125780 294754 125792
rect 307662 125780 307668 125792
rect 294748 125752 307668 125780
rect 294748 125740 294754 125752
rect 307662 125740 307668 125752
rect 307720 125740 307726 125792
rect 169202 125672 169208 125724
rect 169260 125712 169266 125724
rect 214006 125712 214012 125724
rect 169260 125684 214012 125712
rect 169260 125672 169266 125684
rect 214006 125672 214012 125684
rect 214064 125672 214070 125724
rect 289354 125672 289360 125724
rect 289412 125712 289418 125724
rect 306742 125712 306748 125724
rect 289412 125684 306748 125712
rect 289412 125672 289418 125684
rect 306742 125672 306748 125684
rect 306800 125672 306806 125724
rect 166350 125604 166356 125656
rect 166408 125644 166414 125656
rect 213914 125644 213920 125656
rect 166408 125616 213920 125644
rect 166408 125604 166414 125616
rect 213914 125604 213920 125616
rect 213972 125604 213978 125656
rect 271138 125604 271144 125656
rect 271196 125644 271202 125656
rect 307478 125644 307484 125656
rect 271196 125616 307484 125644
rect 271196 125604 271202 125616
rect 307478 125604 307484 125616
rect 307536 125604 307542 125656
rect 252462 125536 252468 125588
rect 252520 125576 252526 125588
rect 304350 125576 304356 125588
rect 252520 125548 304356 125576
rect 252520 125536 252526 125548
rect 304350 125536 304356 125548
rect 304408 125536 304414 125588
rect 252370 125468 252376 125520
rect 252428 125508 252434 125520
rect 265802 125508 265808 125520
rect 252428 125480 265808 125508
rect 252428 125468 252434 125480
rect 265802 125468 265808 125480
rect 265860 125468 265866 125520
rect 252278 124856 252284 124908
rect 252336 124896 252342 124908
rect 300118 124896 300124 124908
rect 252336 124868 300124 124896
rect 252336 124856 252342 124868
rect 300118 124856 300124 124868
rect 300176 124856 300182 124908
rect 300302 124312 300308 124364
rect 300360 124352 300366 124364
rect 306742 124352 306748 124364
rect 300360 124324 306748 124352
rect 300360 124312 300366 124324
rect 306742 124312 306748 124324
rect 306800 124312 306806 124364
rect 173342 124244 173348 124296
rect 173400 124284 173406 124296
rect 213914 124284 213920 124296
rect 173400 124256 213920 124284
rect 173400 124244 173406 124256
rect 213914 124244 213920 124256
rect 213972 124244 213978 124296
rect 304258 124244 304264 124296
rect 304316 124284 304322 124296
rect 307478 124284 307484 124296
rect 304316 124256 307484 124284
rect 304316 124244 304322 124256
rect 307478 124244 307484 124256
rect 307536 124244 307542 124296
rect 170582 124176 170588 124228
rect 170640 124216 170646 124228
rect 214006 124216 214012 124228
rect 170640 124188 214012 124216
rect 170640 124176 170646 124188
rect 214006 124176 214012 124188
rect 214064 124176 214070 124228
rect 290458 124176 290464 124228
rect 290516 124216 290522 124228
rect 307662 124216 307668 124228
rect 290516 124188 307668 124216
rect 290516 124176 290522 124188
rect 307662 124176 307668 124188
rect 307720 124176 307726 124228
rect 252462 124108 252468 124160
rect 252520 124148 252526 124160
rect 268378 124148 268384 124160
rect 252520 124120 268384 124148
rect 252520 124108 252526 124120
rect 268378 124108 268384 124120
rect 268436 124108 268442 124160
rect 324314 124108 324320 124160
rect 324372 124148 324378 124160
rect 342346 124148 342352 124160
rect 324372 124120 342352 124148
rect 324372 124108 324378 124120
rect 342346 124108 342352 124120
rect 342404 124108 342410 124160
rect 252002 124040 252008 124092
rect 252060 124080 252066 124092
rect 261570 124080 261576 124092
rect 252060 124052 261576 124080
rect 252060 124040 252066 124052
rect 261570 124040 261576 124052
rect 261628 124040 261634 124092
rect 323578 124040 323584 124092
rect 323636 124080 323642 124092
rect 324498 124080 324504 124092
rect 323636 124052 324504 124080
rect 323636 124040 323642 124052
rect 324498 124040 324504 124052
rect 324556 124040 324562 124092
rect 252094 123428 252100 123480
rect 252152 123468 252158 123480
rect 301590 123468 301596 123480
rect 252152 123440 301596 123468
rect 252152 123428 252158 123440
rect 301590 123428 301596 123440
rect 301648 123428 301654 123480
rect 211798 123360 211804 123412
rect 211856 123400 211862 123412
rect 214006 123400 214012 123412
rect 211856 123372 214012 123400
rect 211856 123360 211862 123372
rect 214006 123360 214012 123372
rect 214064 123360 214070 123412
rect 300210 122952 300216 123004
rect 300268 122992 300274 123004
rect 307662 122992 307668 123004
rect 300268 122964 307668 122992
rect 300268 122952 300274 122964
rect 307662 122952 307668 122964
rect 307720 122952 307726 123004
rect 302970 122884 302976 122936
rect 303028 122924 303034 122936
rect 307570 122924 307576 122936
rect 303028 122896 307576 122924
rect 303028 122884 303034 122896
rect 307570 122884 307576 122896
rect 307628 122884 307634 122936
rect 174722 122816 174728 122868
rect 174780 122856 174786 122868
rect 213914 122856 213920 122868
rect 174780 122828 213920 122856
rect 174780 122816 174786 122828
rect 213914 122816 213920 122828
rect 213972 122816 213978 122868
rect 283558 122816 283564 122868
rect 283616 122856 283622 122868
rect 306558 122856 306564 122868
rect 283616 122828 306564 122856
rect 283616 122816 283622 122828
rect 306558 122816 306564 122828
rect 306616 122816 306622 122868
rect 252462 122748 252468 122800
rect 252520 122788 252526 122800
rect 296070 122788 296076 122800
rect 252520 122760 296076 122788
rect 252520 122748 252526 122760
rect 296070 122748 296076 122760
rect 296128 122748 296134 122800
rect 324682 122748 324688 122800
rect 324740 122788 324746 122800
rect 343818 122788 343824 122800
rect 324740 122760 343824 122788
rect 324740 122748 324746 122760
rect 343818 122748 343824 122760
rect 343876 122748 343882 122800
rect 252370 122680 252376 122732
rect 252428 122720 252434 122732
rect 269758 122720 269764 122732
rect 252428 122692 269764 122720
rect 252428 122680 252434 122692
rect 269758 122680 269764 122692
rect 269816 122680 269822 122732
rect 324314 122680 324320 122732
rect 324372 122720 324378 122732
rect 338114 122720 338120 122732
rect 324372 122692 338120 122720
rect 324372 122680 324378 122692
rect 338114 122680 338120 122692
rect 338172 122680 338178 122732
rect 252462 122000 252468 122052
rect 252520 122040 252526 122052
rect 260190 122040 260196 122052
rect 252520 122012 260196 122040
rect 252520 122000 252526 122012
rect 260190 122000 260196 122012
rect 260248 122000 260254 122052
rect 297542 121592 297548 121644
rect 297600 121632 297606 121644
rect 307662 121632 307668 121644
rect 297600 121604 307668 121632
rect 297600 121592 297606 121604
rect 307662 121592 307668 121604
rect 307720 121592 307726 121644
rect 207658 121524 207664 121576
rect 207716 121564 207722 121576
rect 214006 121564 214012 121576
rect 207716 121536 214012 121564
rect 207716 121524 207722 121536
rect 214006 121524 214012 121536
rect 214064 121524 214070 121576
rect 293310 121524 293316 121576
rect 293368 121564 293374 121576
rect 307570 121564 307576 121576
rect 293368 121536 307576 121564
rect 293368 121524 293374 121536
rect 307570 121524 307576 121536
rect 307628 121524 307634 121576
rect 180242 121456 180248 121508
rect 180300 121496 180306 121508
rect 213914 121496 213920 121508
rect 180300 121468 213920 121496
rect 180300 121456 180306 121468
rect 213914 121456 213920 121468
rect 213972 121456 213978 121508
rect 268378 121456 268384 121508
rect 268436 121496 268442 121508
rect 307478 121496 307484 121508
rect 268436 121468 307484 121496
rect 268436 121456 268442 121468
rect 307478 121456 307484 121468
rect 307536 121456 307542 121508
rect 251910 121388 251916 121440
rect 251968 121428 251974 121440
rect 287974 121428 287980 121440
rect 251968 121400 287980 121428
rect 251968 121388 251974 121400
rect 287974 121388 287980 121400
rect 288032 121388 288038 121440
rect 324406 121388 324412 121440
rect 324464 121428 324470 121440
rect 339494 121428 339500 121440
rect 324464 121400 339500 121428
rect 324464 121388 324470 121400
rect 339494 121388 339500 121400
rect 339552 121388 339558 121440
rect 252462 121320 252468 121372
rect 252520 121360 252526 121372
rect 265710 121360 265716 121372
rect 252520 121332 265716 121360
rect 252520 121320 252526 121332
rect 265710 121320 265716 121332
rect 265768 121320 265774 121372
rect 324314 121320 324320 121372
rect 324372 121360 324378 121372
rect 335538 121360 335544 121372
rect 324372 121332 335544 121360
rect 324372 121320 324378 121332
rect 335538 121320 335544 121332
rect 335596 121320 335602 121372
rect 252370 121252 252376 121304
rect 252428 121292 252434 121304
rect 258718 121292 258724 121304
rect 252428 121264 258724 121292
rect 252428 121252 252434 121264
rect 258718 121252 258724 121264
rect 258776 121252 258782 121304
rect 301682 120232 301688 120284
rect 301740 120272 301746 120284
rect 307662 120272 307668 120284
rect 301740 120244 307668 120272
rect 301740 120232 301746 120244
rect 307662 120232 307668 120244
rect 307720 120232 307726 120284
rect 185578 120164 185584 120216
rect 185636 120204 185642 120216
rect 214006 120204 214012 120216
rect 185636 120176 214012 120204
rect 185636 120164 185642 120176
rect 214006 120164 214012 120176
rect 214064 120164 214070 120216
rect 287882 120164 287888 120216
rect 287940 120204 287946 120216
rect 307478 120204 307484 120216
rect 287940 120176 307484 120204
rect 287940 120164 287946 120176
rect 307478 120164 307484 120176
rect 307536 120164 307542 120216
rect 167638 120096 167644 120148
rect 167696 120136 167702 120148
rect 213914 120136 213920 120148
rect 167696 120108 213920 120136
rect 167696 120096 167702 120108
rect 213914 120096 213920 120108
rect 213972 120096 213978 120148
rect 266998 120096 267004 120148
rect 267056 120136 267062 120148
rect 307570 120136 307576 120148
rect 267056 120108 307576 120136
rect 267056 120096 267062 120108
rect 307570 120096 307576 120108
rect 307628 120096 307634 120148
rect 252462 120028 252468 120080
rect 252520 120068 252526 120080
rect 296254 120068 296260 120080
rect 252520 120040 296260 120068
rect 252520 120028 252526 120040
rect 296254 120028 296260 120040
rect 296312 120028 296318 120080
rect 251358 119960 251364 120012
rect 251416 120000 251422 120012
rect 262950 120000 262956 120012
rect 251416 119972 262956 120000
rect 251416 119960 251422 119972
rect 262950 119960 262956 119972
rect 263008 119960 263014 120012
rect 263042 119348 263048 119400
rect 263100 119388 263106 119400
rect 307202 119388 307208 119400
rect 263100 119360 307208 119388
rect 263100 119348 263106 119360
rect 307202 119348 307208 119360
rect 307260 119348 307266 119400
rect 210510 118804 210516 118856
rect 210568 118844 210574 118856
rect 214098 118844 214104 118856
rect 210568 118816 214104 118844
rect 210568 118804 210574 118816
rect 214098 118804 214104 118816
rect 214156 118804 214162 118856
rect 296162 118804 296168 118856
rect 296220 118844 296226 118856
rect 306742 118844 306748 118856
rect 296220 118816 306748 118844
rect 296220 118804 296226 118816
rect 306742 118804 306748 118816
rect 306800 118804 306806 118856
rect 196618 118736 196624 118788
rect 196676 118776 196682 118788
rect 214006 118776 214012 118788
rect 196676 118748 214012 118776
rect 196676 118736 196682 118748
rect 214006 118736 214012 118748
rect 214064 118736 214070 118788
rect 251174 118736 251180 118788
rect 251232 118776 251238 118788
rect 253198 118776 253204 118788
rect 251232 118748 253204 118776
rect 251232 118736 251238 118748
rect 253198 118736 253204 118748
rect 253256 118736 253262 118788
rect 299014 118736 299020 118788
rect 299072 118776 299078 118788
rect 307662 118776 307668 118788
rect 299072 118748 307668 118776
rect 299072 118736 299078 118748
rect 307662 118736 307668 118748
rect 307720 118736 307726 118788
rect 166442 118668 166448 118720
rect 166500 118708 166506 118720
rect 213914 118708 213920 118720
rect 166500 118680 213920 118708
rect 166500 118668 166506 118680
rect 213914 118668 213920 118680
rect 213972 118668 213978 118720
rect 251818 118600 251824 118652
rect 251876 118640 251882 118652
rect 293586 118640 293592 118652
rect 251876 118612 293592 118640
rect 251876 118600 251882 118612
rect 293586 118600 293592 118612
rect 293644 118600 293650 118652
rect 324406 118600 324412 118652
rect 324464 118640 324470 118652
rect 341058 118640 341064 118652
rect 324464 118612 341064 118640
rect 324464 118600 324470 118612
rect 341058 118600 341064 118612
rect 341116 118600 341122 118652
rect 252462 118532 252468 118584
rect 252520 118572 252526 118584
rect 260098 118572 260104 118584
rect 252520 118544 260104 118572
rect 252520 118532 252526 118544
rect 260098 118532 260104 118544
rect 260156 118532 260162 118584
rect 324314 118532 324320 118584
rect 324372 118572 324378 118584
rect 339586 118572 339592 118584
rect 324372 118544 339592 118572
rect 324372 118532 324378 118544
rect 339586 118532 339592 118544
rect 339644 118532 339650 118584
rect 167730 117920 167736 117972
rect 167788 117960 167794 117972
rect 213270 117960 213276 117972
rect 167788 117932 213276 117960
rect 167788 117920 167794 117932
rect 213270 117920 213276 117932
rect 213328 117920 213334 117972
rect 251634 117920 251640 117972
rect 251692 117960 251698 117972
rect 298830 117960 298836 117972
rect 251692 117932 298836 117960
rect 251692 117920 251698 117932
rect 298830 117920 298836 117932
rect 298888 117920 298894 117972
rect 300394 117444 300400 117496
rect 300452 117484 300458 117496
rect 307570 117484 307576 117496
rect 300452 117456 307576 117484
rect 300452 117444 300458 117456
rect 307570 117444 307576 117456
rect 307628 117444 307634 117496
rect 296070 117376 296076 117428
rect 296128 117416 296134 117428
rect 307662 117416 307668 117428
rect 296128 117388 307668 117416
rect 296128 117376 296134 117388
rect 307662 117376 307668 117388
rect 307720 117376 307726 117428
rect 210602 117308 210608 117360
rect 210660 117348 210666 117360
rect 213914 117348 213920 117360
rect 210660 117320 213920 117348
rect 210660 117308 210666 117320
rect 213914 117308 213920 117320
rect 213972 117308 213978 117360
rect 293402 117308 293408 117360
rect 293460 117348 293466 117360
rect 307478 117348 307484 117360
rect 293460 117320 307484 117348
rect 293460 117308 293466 117320
rect 307478 117308 307484 117320
rect 307536 117308 307542 117360
rect 251910 117240 251916 117292
rect 251968 117280 251974 117292
rect 291930 117280 291936 117292
rect 251968 117252 291936 117280
rect 251968 117240 251974 117252
rect 291930 117240 291936 117252
rect 291988 117240 291994 117292
rect 324406 117240 324412 117292
rect 324464 117280 324470 117292
rect 336918 117280 336924 117292
rect 324464 117252 336924 117280
rect 324464 117240 324470 117252
rect 336918 117240 336924 117252
rect 336976 117240 336982 117292
rect 252370 117172 252376 117224
rect 252428 117212 252434 117224
rect 261478 117212 261484 117224
rect 252428 117184 261484 117212
rect 252428 117172 252434 117184
rect 261478 117172 261484 117184
rect 261536 117172 261542 117224
rect 324314 117172 324320 117224
rect 324372 117212 324378 117224
rect 332686 117212 332692 117224
rect 324372 117184 332692 117212
rect 324372 117172 324378 117184
rect 332686 117172 332692 117184
rect 332744 117172 332750 117224
rect 252462 117104 252468 117156
rect 252520 117144 252526 117156
rect 258902 117144 258908 117156
rect 252520 117116 258908 117144
rect 252520 117104 252526 117116
rect 258902 117104 258908 117116
rect 258960 117104 258966 117156
rect 189810 116016 189816 116068
rect 189868 116056 189874 116068
rect 213914 116056 213920 116068
rect 189868 116028 213920 116056
rect 189868 116016 189874 116028
rect 213914 116016 213920 116028
rect 213972 116016 213978 116068
rect 292022 116016 292028 116068
rect 292080 116056 292086 116068
rect 307662 116056 307668 116068
rect 292080 116028 307668 116056
rect 292080 116016 292086 116028
rect 307662 116016 307668 116028
rect 307720 116016 307726 116068
rect 169294 115948 169300 116000
rect 169352 115988 169358 116000
rect 214006 115988 214012 116000
rect 169352 115960 214012 115988
rect 169352 115948 169358 115960
rect 214006 115948 214012 115960
rect 214064 115948 214070 116000
rect 265710 115948 265716 116000
rect 265768 115988 265774 116000
rect 306742 115988 306748 116000
rect 265768 115960 306748 115988
rect 265768 115948 265774 115960
rect 306742 115948 306748 115960
rect 306800 115948 306806 116000
rect 252462 115880 252468 115932
rect 252520 115920 252526 115932
rect 275370 115920 275376 115932
rect 252520 115892 275376 115920
rect 252520 115880 252526 115892
rect 275370 115880 275376 115892
rect 275428 115880 275434 115932
rect 324314 115880 324320 115932
rect 324372 115920 324378 115932
rect 336826 115920 336832 115932
rect 324372 115892 336832 115920
rect 324372 115880 324378 115892
rect 336826 115880 336832 115892
rect 336884 115880 336890 115932
rect 252370 115812 252376 115864
rect 252428 115852 252434 115864
rect 262858 115852 262864 115864
rect 252428 115824 262864 115852
rect 252428 115812 252434 115824
rect 262858 115812 262864 115824
rect 262916 115812 262922 115864
rect 168190 115200 168196 115252
rect 168248 115240 168254 115252
rect 178862 115240 178868 115252
rect 168248 115212 178868 115240
rect 168248 115200 168254 115212
rect 178862 115200 178868 115212
rect 178920 115200 178926 115252
rect 211982 114588 211988 114640
rect 212040 114628 212046 114640
rect 214006 114628 214012 114640
rect 212040 114600 214012 114628
rect 212040 114588 212046 114600
rect 214006 114588 214012 114600
rect 214064 114588 214070 114640
rect 282178 114588 282184 114640
rect 282236 114628 282242 114640
rect 307662 114628 307668 114640
rect 282236 114600 307668 114628
rect 282236 114588 282242 114600
rect 307662 114588 307668 114600
rect 307720 114588 307726 114640
rect 178954 114520 178960 114572
rect 179012 114560 179018 114572
rect 213914 114560 213920 114572
rect 179012 114532 213920 114560
rect 179012 114520 179018 114532
rect 213914 114520 213920 114532
rect 213972 114520 213978 114572
rect 264330 114520 264336 114572
rect 264388 114560 264394 114572
rect 306742 114560 306748 114572
rect 264388 114532 306748 114560
rect 264388 114520 264394 114532
rect 306742 114520 306748 114532
rect 306800 114520 306806 114572
rect 252462 114452 252468 114504
rect 252520 114492 252526 114504
rect 282362 114492 282368 114504
rect 252520 114464 282368 114492
rect 252520 114452 252526 114464
rect 282362 114452 282368 114464
rect 282420 114452 282426 114504
rect 324314 114452 324320 114504
rect 324372 114492 324378 114504
rect 340966 114492 340972 114504
rect 324372 114464 340972 114492
rect 324372 114452 324378 114464
rect 340966 114452 340972 114464
rect 341024 114452 341030 114504
rect 252370 114384 252376 114436
rect 252428 114424 252434 114436
rect 276750 114424 276756 114436
rect 252428 114396 276756 114424
rect 252428 114384 252434 114396
rect 276750 114384 276756 114396
rect 276808 114384 276814 114436
rect 324406 114384 324412 114436
rect 324464 114424 324470 114436
rect 334066 114424 334072 114436
rect 324464 114396 334072 114424
rect 324464 114384 324470 114396
rect 334066 114384 334072 114396
rect 334124 114384 334130 114436
rect 252094 113704 252100 113756
rect 252152 113744 252158 113756
rect 254670 113744 254676 113756
rect 252152 113716 254676 113744
rect 252152 113704 252158 113716
rect 254670 113704 254676 113716
rect 254728 113704 254734 113756
rect 298830 113296 298836 113348
rect 298888 113336 298894 113348
rect 306742 113336 306748 113348
rect 298888 113308 306748 113336
rect 298888 113296 298894 113308
rect 306742 113296 306748 113308
rect 306800 113296 306806 113348
rect 184198 113228 184204 113280
rect 184256 113268 184262 113280
rect 214006 113268 214012 113280
rect 184256 113240 214012 113268
rect 184256 113228 184262 113240
rect 214006 113228 214012 113240
rect 214064 113228 214070 113280
rect 291930 113228 291936 113280
rect 291988 113268 291994 113280
rect 307570 113268 307576 113280
rect 291988 113240 307576 113268
rect 291988 113228 291994 113240
rect 307570 113228 307576 113240
rect 307628 113228 307634 113280
rect 171962 113160 171968 113212
rect 172020 113200 172026 113212
rect 213914 113200 213920 113212
rect 172020 113172 213920 113200
rect 172020 113160 172026 113172
rect 213914 113160 213920 113172
rect 213972 113160 213978 113212
rect 279602 113160 279608 113212
rect 279660 113200 279666 113212
rect 307662 113200 307668 113212
rect 279660 113172 307668 113200
rect 279660 113160 279666 113172
rect 307662 113160 307668 113172
rect 307720 113160 307726 113212
rect 252462 113092 252468 113144
rect 252520 113132 252526 113144
rect 300486 113132 300492 113144
rect 252520 113104 300492 113132
rect 252520 113092 252526 113104
rect 300486 113092 300492 113104
rect 300544 113092 300550 113144
rect 324314 113092 324320 113144
rect 324372 113132 324378 113144
rect 335446 113132 335452 113144
rect 324372 113104 335452 113132
rect 324372 113092 324378 113104
rect 335446 113092 335452 113104
rect 335504 113092 335510 113144
rect 252370 112412 252376 112464
rect 252428 112452 252434 112464
rect 264422 112452 264428 112464
rect 252428 112424 264428 112452
rect 252428 112412 252434 112424
rect 264422 112412 264428 112424
rect 264480 112412 264486 112464
rect 269390 112412 269396 112464
rect 269448 112452 269454 112464
rect 307018 112452 307024 112464
rect 269448 112424 307024 112452
rect 269448 112412 269454 112424
rect 307018 112412 307024 112424
rect 307076 112412 307082 112464
rect 177390 111868 177396 111920
rect 177448 111908 177454 111920
rect 214006 111908 214012 111920
rect 177448 111880 214012 111908
rect 177448 111868 177454 111880
rect 214006 111868 214012 111880
rect 214064 111868 214070 111920
rect 300118 111868 300124 111920
rect 300176 111908 300182 111920
rect 307570 111908 307576 111920
rect 300176 111880 307576 111908
rect 300176 111868 300182 111880
rect 307570 111868 307576 111880
rect 307628 111868 307634 111920
rect 170674 111800 170680 111852
rect 170732 111840 170738 111852
rect 213914 111840 213920 111852
rect 170732 111812 213920 111840
rect 170732 111800 170738 111812
rect 213914 111800 213920 111812
rect 213972 111800 213978 111852
rect 251542 111800 251548 111852
rect 251600 111840 251606 111852
rect 254762 111840 254768 111852
rect 251600 111812 254768 111840
rect 251600 111800 251606 111812
rect 254762 111800 254768 111812
rect 254820 111800 254826 111852
rect 297450 111800 297456 111852
rect 297508 111840 297514 111852
rect 307662 111840 307668 111852
rect 297508 111812 307668 111840
rect 297508 111800 297514 111812
rect 307662 111800 307668 111812
rect 307720 111800 307726 111852
rect 167914 111732 167920 111784
rect 167972 111772 167978 111784
rect 174814 111772 174820 111784
rect 167972 111744 174820 111772
rect 167972 111732 167978 111744
rect 174814 111732 174820 111744
rect 174872 111732 174878 111784
rect 252462 111732 252468 111784
rect 252520 111772 252526 111784
rect 301498 111772 301504 111784
rect 252520 111744 301504 111772
rect 252520 111732 252526 111744
rect 301498 111732 301504 111744
rect 301556 111732 301562 111784
rect 324314 111732 324320 111784
rect 324372 111772 324378 111784
rect 342254 111772 342260 111784
rect 324372 111744 342260 111772
rect 324372 111732 324378 111744
rect 342254 111732 342260 111744
rect 342312 111732 342318 111784
rect 252278 111664 252284 111716
rect 252336 111704 252342 111716
rect 257338 111704 257344 111716
rect 252336 111676 257344 111704
rect 252336 111664 252342 111676
rect 257338 111664 257344 111676
rect 257396 111664 257402 111716
rect 251726 111052 251732 111104
rect 251784 111092 251790 111104
rect 297634 111092 297640 111104
rect 251784 111064 297640 111092
rect 251784 111052 251790 111064
rect 297634 111052 297640 111064
rect 297692 111052 297698 111104
rect 301774 110576 301780 110628
rect 301832 110616 301838 110628
rect 307570 110616 307576 110628
rect 301832 110588 307576 110616
rect 301832 110576 301838 110588
rect 307570 110576 307576 110588
rect 307628 110576 307634 110628
rect 202230 110508 202236 110560
rect 202288 110548 202294 110560
rect 213914 110548 213920 110560
rect 202288 110520 213920 110548
rect 202288 110508 202294 110520
rect 213914 110508 213920 110520
rect 213972 110508 213978 110560
rect 303154 110508 303160 110560
rect 303212 110548 303218 110560
rect 307662 110548 307668 110560
rect 303212 110520 307668 110548
rect 303212 110508 303218 110520
rect 307662 110508 307668 110520
rect 307720 110508 307726 110560
rect 199378 110440 199384 110492
rect 199436 110480 199442 110492
rect 214006 110480 214012 110492
rect 199436 110452 214012 110480
rect 199436 110440 199442 110452
rect 214006 110440 214012 110452
rect 214064 110440 214070 110492
rect 296254 110440 296260 110492
rect 296312 110480 296318 110492
rect 307478 110480 307484 110492
rect 296312 110452 307484 110480
rect 296312 110440 296318 110452
rect 307478 110440 307484 110452
rect 307536 110440 307542 110492
rect 252462 110372 252468 110424
rect 252520 110412 252526 110424
rect 289170 110412 289176 110424
rect 252520 110384 289176 110412
rect 252520 110372 252526 110384
rect 289170 110372 289176 110384
rect 289228 110372 289234 110424
rect 251266 110304 251272 110356
rect 251324 110344 251330 110356
rect 257522 110344 257528 110356
rect 251324 110316 257528 110344
rect 251324 110304 251330 110316
rect 257522 110304 257528 110316
rect 257580 110304 257586 110356
rect 251910 109284 251916 109336
rect 251968 109324 251974 109336
rect 256142 109324 256148 109336
rect 251968 109296 256148 109324
rect 251968 109284 251974 109296
rect 256142 109284 256148 109296
rect 256200 109284 256206 109336
rect 304534 109148 304540 109200
rect 304592 109188 304598 109200
rect 307478 109188 307484 109200
rect 304592 109160 307484 109188
rect 304592 109148 304598 109160
rect 307478 109148 307484 109160
rect 307536 109148 307542 109200
rect 278222 109080 278228 109132
rect 278280 109120 278286 109132
rect 307570 109120 307576 109132
rect 278280 109092 307576 109120
rect 278280 109080 278286 109092
rect 307570 109080 307576 109092
rect 307628 109080 307634 109132
rect 206370 109012 206376 109064
rect 206428 109052 206434 109064
rect 213914 109052 213920 109064
rect 206428 109024 213920 109052
rect 206428 109012 206434 109024
rect 213914 109012 213920 109024
rect 213972 109012 213978 109064
rect 261478 109012 261484 109064
rect 261536 109052 261542 109064
rect 307662 109052 307668 109064
rect 261536 109024 307668 109052
rect 261536 109012 261542 109024
rect 307662 109012 307668 109024
rect 307720 109012 307726 109064
rect 251358 108944 251364 108996
rect 251416 108984 251422 108996
rect 303062 108984 303068 108996
rect 251416 108956 303068 108984
rect 251416 108944 251422 108956
rect 303062 108944 303068 108956
rect 303120 108944 303126 108996
rect 252462 108876 252468 108928
rect 252520 108916 252526 108928
rect 282454 108916 282460 108928
rect 252520 108888 282460 108916
rect 252520 108876 252526 108888
rect 282454 108876 282460 108888
rect 282512 108876 282518 108928
rect 324314 107992 324320 108044
rect 324372 108032 324378 108044
rect 327258 108032 327264 108044
rect 324372 108004 327264 108032
rect 324372 107992 324378 108004
rect 327258 107992 327264 108004
rect 327316 107992 327322 108044
rect 251174 107856 251180 107908
rect 251232 107896 251238 107908
rect 253474 107896 253480 107908
rect 251232 107868 253480 107896
rect 251232 107856 251238 107868
rect 253474 107856 253480 107868
rect 253532 107856 253538 107908
rect 282362 107856 282368 107908
rect 282420 107896 282426 107908
rect 307662 107896 307668 107908
rect 282420 107868 307668 107896
rect 282420 107856 282426 107868
rect 307662 107856 307668 107868
rect 307720 107856 307726 107908
rect 203610 107720 203616 107772
rect 203668 107760 203674 107772
rect 214006 107760 214012 107772
rect 203668 107732 214012 107760
rect 203668 107720 203674 107732
rect 214006 107720 214012 107732
rect 214064 107720 214070 107772
rect 301590 107720 301596 107772
rect 301648 107760 301654 107772
rect 306742 107760 306748 107772
rect 301648 107732 306748 107760
rect 301648 107720 301654 107732
rect 306742 107720 306748 107732
rect 306800 107720 306806 107772
rect 174814 107652 174820 107704
rect 174872 107692 174878 107704
rect 213914 107692 213920 107704
rect 174872 107664 213920 107692
rect 174872 107652 174878 107664
rect 213914 107652 213920 107664
rect 213972 107652 213978 107704
rect 304350 107652 304356 107704
rect 304408 107692 304414 107704
rect 307570 107692 307576 107704
rect 304408 107664 307576 107692
rect 304408 107652 304414 107664
rect 307570 107652 307576 107664
rect 307628 107652 307634 107704
rect 251358 107584 251364 107636
rect 251416 107624 251422 107636
rect 280890 107624 280896 107636
rect 251416 107596 280896 107624
rect 251416 107584 251422 107596
rect 280890 107584 280896 107596
rect 280948 107584 280954 107636
rect 252462 107516 252468 107568
rect 252520 107556 252526 107568
rect 269390 107556 269396 107568
rect 252520 107528 269396 107556
rect 252520 107516 252526 107528
rect 269390 107516 269396 107528
rect 269448 107516 269454 107568
rect 301498 106428 301504 106480
rect 301556 106468 301562 106480
rect 307478 106468 307484 106480
rect 301556 106440 307484 106468
rect 301556 106428 301562 106440
rect 307478 106428 307484 106440
rect 307536 106428 307542 106480
rect 283650 106360 283656 106412
rect 283708 106400 283714 106412
rect 307570 106400 307576 106412
rect 283708 106372 307576 106400
rect 283708 106360 283714 106372
rect 307570 106360 307576 106372
rect 307628 106360 307634 106412
rect 167730 106292 167736 106344
rect 167788 106332 167794 106344
rect 213914 106332 213920 106344
rect 167788 106304 213920 106332
rect 167788 106292 167794 106304
rect 213914 106292 213920 106304
rect 213972 106292 213978 106344
rect 269850 106292 269856 106344
rect 269908 106332 269914 106344
rect 307662 106332 307668 106344
rect 269908 106304 307668 106332
rect 269908 106292 269914 106304
rect 307662 106292 307668 106304
rect 307720 106292 307726 106344
rect 252002 106224 252008 106276
rect 252060 106264 252066 106276
rect 279694 106264 279700 106276
rect 252060 106236 279700 106264
rect 252060 106224 252066 106236
rect 279694 106224 279700 106236
rect 279752 106224 279758 106276
rect 252278 106156 252284 106208
rect 252336 106196 252342 106208
rect 256234 106196 256240 106208
rect 252336 106168 256240 106196
rect 252336 106156 252342 106168
rect 256234 106156 256240 106168
rect 256292 106156 256298 106208
rect 252002 105544 252008 105596
rect 252060 105584 252066 105596
rect 305822 105584 305828 105596
rect 252060 105556 305828 105584
rect 252060 105544 252066 105556
rect 305822 105544 305828 105556
rect 305880 105544 305886 105596
rect 280890 105000 280896 105052
rect 280948 105040 280954 105052
rect 307662 105040 307668 105052
rect 280948 105012 307668 105040
rect 280948 105000 280954 105012
rect 307662 105000 307668 105012
rect 307720 105000 307726 105052
rect 212074 104932 212080 104984
rect 212132 104972 212138 104984
rect 214006 104972 214012 104984
rect 212132 104944 214012 104972
rect 212132 104932 212138 104944
rect 214006 104932 214012 104944
rect 214064 104932 214070 104984
rect 289170 104932 289176 104984
rect 289228 104972 289234 104984
rect 306558 104972 306564 104984
rect 289228 104944 306564 104972
rect 289228 104932 289234 104944
rect 306558 104932 306564 104944
rect 306616 104932 306622 104984
rect 209038 104864 209044 104916
rect 209096 104904 209102 104916
rect 213914 104904 213920 104916
rect 209096 104876 213920 104904
rect 209096 104864 209102 104876
rect 213914 104864 213920 104876
rect 213972 104864 213978 104916
rect 252462 104796 252468 104848
rect 252520 104836 252526 104848
rect 305914 104836 305920 104848
rect 252520 104808 305920 104836
rect 252520 104796 252526 104808
rect 305914 104796 305920 104808
rect 305972 104796 305978 104848
rect 251542 104116 251548 104168
rect 251600 104156 251606 104168
rect 286410 104156 286416 104168
rect 251600 104128 286416 104156
rect 251600 104116 251606 104128
rect 286410 104116 286416 104128
rect 286468 104116 286474 104168
rect 253198 103640 253204 103692
rect 253256 103680 253262 103692
rect 307662 103680 307668 103692
rect 253256 103652 307668 103680
rect 253256 103640 253262 103652
rect 307662 103640 307668 103652
rect 307720 103640 307726 103692
rect 287974 103572 287980 103624
rect 288032 103612 288038 103624
rect 307570 103612 307576 103624
rect 288032 103584 307576 103612
rect 288032 103572 288038 103584
rect 307570 103572 307576 103584
rect 307628 103572 307634 103624
rect 209130 103504 209136 103556
rect 209188 103544 209194 103556
rect 213914 103544 213920 103556
rect 209188 103516 213920 103544
rect 209188 103504 209194 103516
rect 213914 103504 213920 103516
rect 213972 103504 213978 103556
rect 252462 103436 252468 103488
rect 252520 103476 252526 103488
rect 267090 103476 267096 103488
rect 252520 103448 267096 103476
rect 252520 103436 252526 103448
rect 267090 103436 267096 103448
rect 267148 103436 267154 103488
rect 251174 102756 251180 102808
rect 251232 102796 251238 102808
rect 253382 102796 253388 102808
rect 251232 102768 253388 102796
rect 251232 102756 251238 102768
rect 253382 102756 253388 102768
rect 253440 102756 253446 102808
rect 298922 102280 298928 102332
rect 298980 102320 298986 102332
rect 307478 102320 307484 102332
rect 298980 102292 307484 102320
rect 298980 102280 298986 102292
rect 307478 102280 307484 102292
rect 307536 102280 307542 102332
rect 252094 102212 252100 102264
rect 252152 102252 252158 102264
rect 257430 102252 257436 102264
rect 252152 102224 257436 102252
rect 252152 102212 252158 102224
rect 257430 102212 257436 102224
rect 257488 102212 257494 102264
rect 269758 102212 269764 102264
rect 269816 102252 269822 102264
rect 306742 102252 306748 102264
rect 269816 102224 306748 102252
rect 269816 102212 269822 102224
rect 306742 102212 306748 102224
rect 306800 102212 306806 102264
rect 204898 102144 204904 102196
rect 204956 102184 204962 102196
rect 213914 102184 213920 102196
rect 204956 102156 213920 102184
rect 204956 102144 204962 102156
rect 213914 102144 213920 102156
rect 213972 102144 213978 102196
rect 257338 102144 257344 102196
rect 257396 102184 257402 102196
rect 306926 102184 306932 102196
rect 257396 102156 306932 102184
rect 257396 102144 257402 102156
rect 306926 102144 306932 102156
rect 306984 102144 306990 102196
rect 252462 102076 252468 102128
rect 252520 102116 252526 102128
rect 293494 102116 293500 102128
rect 252520 102088 293500 102116
rect 252520 102076 252526 102088
rect 293494 102076 293500 102088
rect 293552 102076 293558 102128
rect 252370 102008 252376 102060
rect 252428 102048 252434 102060
rect 286318 102048 286324 102060
rect 252428 102020 286324 102048
rect 252428 102008 252434 102020
rect 286318 102008 286324 102020
rect 286376 102008 286382 102060
rect 303062 100852 303068 100904
rect 303120 100892 303126 100904
rect 307570 100892 307576 100904
rect 303120 100864 307576 100892
rect 303120 100852 303126 100864
rect 307570 100852 307576 100864
rect 307628 100852 307634 100904
rect 207842 100784 207848 100836
rect 207900 100824 207906 100836
rect 214006 100824 214012 100836
rect 207900 100796 214012 100824
rect 207900 100784 207906 100796
rect 214006 100784 214012 100796
rect 214064 100784 214070 100836
rect 293586 100784 293592 100836
rect 293644 100824 293650 100836
rect 307662 100824 307668 100836
rect 293644 100796 307668 100824
rect 293644 100784 293650 100796
rect 307662 100784 307668 100796
rect 307720 100784 307726 100836
rect 172054 100716 172060 100768
rect 172112 100756 172118 100768
rect 213914 100756 213920 100768
rect 172112 100728 213920 100756
rect 172112 100716 172118 100728
rect 213914 100716 213920 100728
rect 213972 100716 213978 100768
rect 286410 100716 286416 100768
rect 286468 100756 286474 100768
rect 307478 100756 307484 100768
rect 286468 100728 307484 100756
rect 286468 100716 286474 100728
rect 307478 100716 307484 100728
rect 307536 100716 307542 100768
rect 252094 100648 252100 100700
rect 252152 100688 252158 100700
rect 304442 100688 304448 100700
rect 252152 100660 304448 100688
rect 252152 100648 252158 100660
rect 304442 100648 304448 100660
rect 304500 100648 304506 100700
rect 395338 100648 395344 100700
rect 395396 100688 395402 100700
rect 580166 100688 580172 100700
rect 395396 100660 580172 100688
rect 395396 100648 395402 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 252462 100580 252468 100632
rect 252520 100620 252526 100632
rect 292114 100620 292120 100632
rect 252520 100592 292120 100620
rect 252520 100580 252526 100592
rect 292114 100580 292120 100592
rect 292172 100580 292178 100632
rect 251174 100104 251180 100156
rect 251232 100144 251238 100156
rect 253290 100144 253296 100156
rect 251232 100116 253296 100144
rect 251232 100104 251238 100116
rect 253290 100104 253296 100116
rect 253348 100104 253354 100156
rect 173434 99424 173440 99476
rect 173492 99464 173498 99476
rect 213914 99464 213920 99476
rect 173492 99436 213920 99464
rect 173492 99424 173498 99436
rect 213914 99424 213920 99436
rect 213972 99424 213978 99476
rect 304626 99424 304632 99476
rect 304684 99464 304690 99476
rect 307478 99464 307484 99476
rect 304684 99436 307484 99464
rect 304684 99424 304690 99436
rect 307478 99424 307484 99436
rect 307536 99424 307542 99476
rect 167914 99356 167920 99408
rect 167972 99396 167978 99408
rect 214006 99396 214012 99408
rect 167972 99368 214012 99396
rect 167972 99356 167978 99368
rect 214006 99356 214012 99368
rect 214064 99356 214070 99408
rect 289262 99356 289268 99408
rect 289320 99396 289326 99408
rect 307662 99396 307668 99408
rect 289320 99368 307668 99396
rect 289320 99356 289326 99368
rect 307662 99356 307668 99368
rect 307720 99356 307726 99408
rect 252186 99288 252192 99340
rect 252244 99328 252250 99340
rect 269942 99328 269948 99340
rect 252244 99300 269948 99328
rect 252244 99288 252250 99300
rect 269942 99288 269948 99300
rect 270000 99288 270006 99340
rect 252278 99152 252284 99204
rect 252336 99192 252342 99204
rect 256050 99192 256056 99204
rect 252336 99164 256056 99192
rect 252336 99152 252342 99164
rect 256050 99152 256056 99164
rect 256108 99152 256114 99204
rect 251174 98608 251180 98660
rect 251232 98648 251238 98660
rect 254578 98648 254584 98660
rect 251232 98620 254584 98648
rect 251232 98608 251238 98620
rect 254578 98608 254584 98620
rect 254636 98608 254642 98660
rect 294782 98132 294788 98184
rect 294840 98172 294846 98184
rect 307662 98172 307668 98184
rect 294840 98144 307668 98172
rect 294840 98132 294846 98144
rect 307662 98132 307668 98144
rect 307720 98132 307726 98184
rect 286318 98064 286324 98116
rect 286376 98104 286382 98116
rect 307478 98104 307484 98116
rect 286376 98076 307484 98104
rect 286376 98064 286382 98076
rect 307478 98064 307484 98076
rect 307536 98064 307542 98116
rect 167822 97996 167828 98048
rect 167880 98036 167886 98048
rect 213914 98036 213920 98048
rect 167880 98008 213920 98036
rect 167880 97996 167886 98008
rect 213914 97996 213920 98008
rect 213972 97996 213978 98048
rect 260098 97996 260104 98048
rect 260156 98036 260162 98048
rect 307570 98036 307576 98048
rect 260156 98008 307576 98036
rect 260156 97996 260162 98008
rect 307570 97996 307576 98008
rect 307628 97996 307634 98048
rect 252462 97860 252468 97912
rect 252520 97900 252526 97912
rect 263042 97900 263048 97912
rect 252520 97872 263048 97900
rect 252520 97860 252526 97872
rect 263042 97860 263048 97872
rect 263100 97860 263106 97912
rect 249518 97520 249524 97572
rect 249576 97560 249582 97572
rect 255958 97560 255964 97572
rect 249576 97532 255964 97560
rect 249576 97520 249582 97532
rect 255958 97520 255964 97532
rect 256016 97520 256022 97572
rect 166534 97248 166540 97300
rect 166592 97288 166598 97300
rect 214558 97288 214564 97300
rect 166592 97260 214564 97288
rect 166592 97248 166598 97260
rect 214558 97248 214564 97260
rect 214616 97248 214622 97300
rect 292114 96704 292120 96756
rect 292172 96744 292178 96756
rect 306742 96744 306748 96756
rect 292172 96716 306748 96744
rect 292172 96704 292178 96716
rect 306742 96704 306748 96716
rect 306800 96704 306806 96756
rect 164878 96636 164884 96688
rect 164936 96676 164942 96688
rect 213914 96676 213920 96688
rect 164936 96648 213920 96676
rect 164936 96636 164942 96648
rect 213914 96636 213920 96648
rect 213972 96636 213978 96688
rect 256050 96636 256056 96688
rect 256108 96676 256114 96688
rect 307478 96676 307484 96688
rect 256108 96648 307484 96676
rect 256108 96636 256114 96648
rect 307478 96636 307484 96648
rect 307536 96636 307542 96688
rect 278038 96568 278044 96620
rect 278096 96608 278102 96620
rect 321462 96608 321468 96620
rect 278096 96580 321468 96608
rect 278096 96568 278102 96580
rect 321462 96568 321468 96580
rect 321520 96568 321526 96620
rect 250438 95208 250444 95260
rect 250496 95248 250502 95260
rect 307662 95248 307668 95260
rect 250496 95220 307668 95248
rect 250496 95208 250502 95220
rect 307662 95208 307668 95220
rect 307720 95208 307726 95260
rect 196710 95140 196716 95192
rect 196768 95180 196774 95192
rect 324314 95180 324320 95192
rect 196768 95152 324320 95180
rect 196768 95140 196774 95152
rect 324314 95140 324320 95152
rect 324372 95140 324378 95192
rect 308582 95072 308588 95124
rect 308640 95112 308646 95124
rect 321554 95112 321560 95124
rect 308640 95084 321560 95112
rect 308640 95072 308646 95084
rect 321554 95072 321560 95084
rect 321612 95072 321618 95124
rect 309778 95004 309784 95056
rect 309836 95044 309842 95056
rect 324406 95044 324412 95056
rect 309836 95016 324412 95044
rect 309836 95004 309842 95016
rect 324406 95004 324412 95016
rect 324464 95004 324470 95056
rect 308398 94936 308404 94988
rect 308456 94976 308462 94988
rect 321738 94976 321744 94988
rect 308456 94948 321744 94976
rect 308456 94936 308462 94948
rect 321738 94936 321744 94948
rect 321796 94936 321802 94988
rect 239398 94460 239404 94512
rect 239456 94500 239462 94512
rect 248414 94500 248420 94512
rect 239456 94472 248420 94500
rect 239456 94460 239462 94472
rect 248414 94460 248420 94472
rect 248472 94460 248478 94512
rect 134334 94120 134340 94172
rect 134392 94160 134398 94172
rect 170490 94160 170496 94172
rect 134392 94132 170496 94160
rect 134392 94120 134398 94132
rect 170490 94120 170496 94132
rect 170548 94120 170554 94172
rect 117958 94052 117964 94104
rect 118016 94092 118022 94104
rect 171870 94092 171876 94104
rect 118016 94064 171876 94092
rect 118016 94052 118022 94064
rect 171870 94052 171876 94064
rect 171928 94052 171934 94104
rect 105446 93984 105452 94036
rect 105504 94024 105510 94036
rect 178954 94024 178960 94036
rect 105504 93996 178960 94024
rect 105504 93984 105510 93996
rect 178954 93984 178960 93996
rect 179012 93984 179018 94036
rect 129366 93916 129372 93968
rect 129424 93956 129430 93968
rect 210418 93956 210424 93968
rect 129424 93928 210424 93956
rect 129424 93916 129430 93928
rect 210418 93916 210424 93928
rect 210476 93916 210482 93968
rect 119522 93848 119528 93900
rect 119580 93888 119586 93900
rect 207658 93888 207664 93900
rect 119580 93860 207664 93888
rect 119580 93848 119586 93860
rect 207658 93848 207664 93860
rect 207716 93848 207722 93900
rect 67358 93780 67364 93832
rect 67416 93820 67422 93832
rect 209038 93820 209044 93832
rect 67416 93792 209044 93820
rect 67416 93780 67422 93792
rect 209038 93780 209044 93792
rect 209096 93780 209102 93832
rect 188338 93712 188344 93764
rect 188396 93752 188402 93764
rect 324498 93752 324504 93764
rect 188396 93724 324504 93752
rect 188396 93712 188402 93724
rect 324498 93712 324504 93724
rect 324556 93712 324562 93764
rect 151722 93372 151728 93424
rect 151780 93412 151786 93424
rect 178678 93412 178684 93424
rect 151780 93384 178684 93412
rect 151780 93372 151786 93384
rect 178678 93372 178684 93384
rect 178736 93372 178742 93424
rect 130746 93304 130752 93356
rect 130804 93344 130810 93356
rect 173158 93344 173164 93356
rect 130804 93316 173164 93344
rect 130804 93304 130810 93316
rect 173158 93304 173164 93316
rect 173216 93304 173222 93356
rect 115842 93236 115848 93288
rect 115900 93276 115906 93288
rect 167638 93276 167644 93288
rect 115900 93248 167644 93276
rect 115900 93236 115906 93248
rect 167638 93236 167644 93248
rect 167696 93236 167702 93288
rect 110690 93168 110696 93220
rect 110748 93208 110754 93220
rect 169110 93208 169116 93220
rect 110748 93180 169116 93208
rect 110748 93168 110754 93180
rect 169110 93168 169116 93180
rect 169168 93168 169174 93220
rect 125502 93100 125508 93152
rect 125560 93140 125566 93152
rect 214834 93140 214840 93152
rect 125560 93112 214840 93140
rect 125560 93100 125566 93112
rect 214834 93100 214840 93112
rect 214892 93100 214898 93152
rect 115474 92420 115480 92472
rect 115532 92460 115538 92472
rect 203518 92460 203524 92472
rect 115532 92432 203524 92460
rect 115532 92420 115538 92432
rect 203518 92420 203524 92432
rect 203576 92420 203582 92472
rect 116762 92352 116768 92404
rect 116820 92392 116826 92404
rect 176102 92392 176108 92404
rect 116820 92364 176108 92392
rect 116820 92352 116826 92364
rect 176102 92352 176108 92364
rect 176160 92352 176166 92404
rect 85666 92284 85672 92336
rect 85724 92324 85730 92336
rect 125502 92324 125508 92336
rect 85724 92296 125508 92324
rect 85724 92284 85730 92296
rect 125502 92284 125508 92296
rect 125560 92284 125566 92336
rect 151538 92284 151544 92336
rect 151596 92324 151602 92336
rect 206278 92324 206284 92336
rect 151596 92296 206284 92324
rect 151596 92284 151602 92296
rect 206278 92284 206284 92296
rect 206336 92284 206342 92336
rect 152090 92216 152096 92268
rect 152148 92256 152154 92268
rect 202138 92256 202144 92268
rect 152148 92228 202144 92256
rect 152148 92216 152154 92228
rect 202138 92216 202144 92228
rect 202196 92216 202202 92268
rect 119706 92148 119712 92200
rect 119764 92188 119770 92200
rect 166534 92188 166540 92200
rect 119764 92160 166540 92188
rect 119764 92148 119770 92160
rect 166534 92148 166540 92160
rect 166592 92148 166598 92200
rect 125778 92080 125784 92132
rect 125836 92120 125842 92132
rect 171778 92120 171784 92132
rect 125836 92092 171784 92120
rect 125836 92080 125842 92092
rect 171778 92080 171784 92092
rect 171836 92080 171842 92132
rect 180058 91740 180064 91792
rect 180116 91780 180122 91792
rect 307294 91780 307300 91792
rect 180116 91752 307300 91780
rect 180116 91740 180122 91752
rect 307294 91740 307300 91752
rect 307352 91740 307358 91792
rect 91646 91060 91652 91112
rect 91704 91100 91710 91112
rect 108298 91100 108304 91112
rect 91704 91072 108304 91100
rect 91704 91060 91710 91072
rect 108298 91060 108304 91072
rect 108356 91060 108362 91112
rect 114186 90992 114192 91044
rect 114244 91032 114250 91044
rect 207750 91032 207756 91044
rect 114244 91004 207756 91032
rect 114244 90992 114250 91004
rect 207750 90992 207756 91004
rect 207808 90992 207814 91044
rect 107746 90924 107752 90976
rect 107804 90964 107810 90976
rect 189810 90964 189816 90976
rect 107804 90936 189816 90964
rect 107804 90924 107810 90936
rect 189810 90924 189816 90936
rect 189868 90924 189874 90976
rect 151446 90856 151452 90908
rect 151504 90896 151510 90908
rect 215938 90896 215944 90908
rect 151504 90868 215944 90896
rect 151504 90856 151510 90868
rect 215938 90856 215944 90868
rect 215996 90856 216002 90908
rect 122466 90788 122472 90840
rect 122524 90828 122530 90840
rect 166258 90828 166264 90840
rect 122524 90800 166264 90828
rect 122524 90788 122530 90800
rect 166258 90788 166264 90800
rect 166316 90788 166322 90840
rect 125502 90720 125508 90772
rect 125560 90760 125566 90772
rect 166350 90760 166356 90772
rect 125560 90732 166356 90760
rect 125560 90720 125566 90732
rect 166350 90720 166356 90732
rect 166408 90720 166414 90772
rect 207658 90312 207664 90364
rect 207716 90352 207722 90364
rect 307110 90352 307116 90364
rect 207716 90324 307116 90352
rect 207716 90312 207722 90324
rect 307110 90312 307116 90324
rect 307168 90312 307174 90364
rect 90542 89632 90548 89684
rect 90600 89672 90606 89684
rect 212074 89672 212080 89684
rect 90600 89644 212080 89672
rect 90600 89632 90606 89644
rect 212074 89632 212080 89644
rect 212132 89632 212138 89684
rect 99742 89564 99748 89616
rect 99800 89604 99806 89616
rect 199378 89604 199384 89616
rect 99800 89576 199384 89604
rect 99800 89564 99806 89576
rect 199378 89564 199384 89576
rect 199436 89564 199442 89616
rect 89346 89496 89352 89548
rect 89404 89536 89410 89548
rect 167914 89536 167920 89548
rect 89404 89508 167920 89536
rect 89404 89496 89410 89508
rect 167914 89496 167920 89508
rect 167972 89496 167978 89548
rect 103146 89428 103152 89480
rect 103204 89468 103210 89480
rect 171962 89468 171968 89480
rect 103204 89440 171968 89468
rect 103204 89428 103210 89440
rect 171962 89428 171968 89440
rect 172020 89428 172026 89480
rect 117130 89360 117136 89412
rect 117188 89400 117194 89412
rect 185578 89400 185584 89412
rect 117188 89372 185584 89400
rect 117188 89360 117194 89372
rect 185578 89360 185584 89372
rect 185636 89360 185642 89412
rect 136450 89292 136456 89344
rect 136508 89332 136514 89344
rect 170398 89332 170404 89344
rect 136508 89304 170404 89332
rect 136508 89292 136514 89304
rect 170398 89292 170404 89304
rect 170456 89292 170462 89344
rect 67266 88272 67272 88324
rect 67324 88312 67330 88324
rect 214742 88312 214748 88324
rect 67324 88284 214748 88312
rect 67324 88272 67330 88284
rect 214742 88272 214748 88284
rect 214800 88272 214806 88324
rect 115290 88204 115296 88256
rect 115348 88244 115354 88256
rect 196618 88244 196624 88256
rect 115348 88216 196624 88244
rect 115348 88204 115354 88216
rect 196618 88204 196624 88216
rect 196676 88204 196682 88256
rect 111978 88136 111984 88188
rect 112036 88176 112042 88188
rect 174630 88176 174636 88188
rect 112036 88148 174636 88176
rect 112036 88136 112042 88148
rect 174630 88136 174636 88148
rect 174688 88136 174694 88188
rect 109218 88068 109224 88120
rect 109276 88108 109282 88120
rect 169294 88108 169300 88120
rect 109276 88080 169300 88108
rect 109276 88068 109282 88080
rect 169294 88068 169300 88080
rect 169352 88068 169358 88120
rect 133138 88000 133144 88052
rect 133196 88040 133202 88052
rect 181438 88040 181444 88052
rect 133196 88012 181444 88040
rect 133196 88000 133202 88012
rect 181438 88000 181444 88012
rect 181496 88000 181502 88052
rect 126514 87932 126520 87984
rect 126572 87972 126578 87984
rect 169202 87972 169208 87984
rect 126572 87944 169208 87972
rect 126572 87932 126578 87944
rect 169202 87932 169208 87944
rect 169260 87932 169266 87984
rect 75362 86912 75368 86964
rect 75420 86952 75426 86964
rect 214558 86952 214564 86964
rect 75420 86924 214564 86952
rect 75420 86912 75426 86924
rect 214558 86912 214564 86924
rect 214616 86912 214622 86964
rect 88058 86844 88064 86896
rect 88116 86884 88122 86896
rect 173434 86884 173440 86896
rect 88116 86856 173440 86884
rect 88116 86844 88122 86856
rect 173434 86844 173440 86856
rect 173492 86844 173498 86896
rect 109770 86776 109776 86828
rect 109828 86816 109834 86828
rect 192478 86816 192484 86828
rect 109828 86788 192484 86816
rect 109828 86776 109834 86788
rect 192478 86776 192484 86788
rect 192536 86776 192542 86828
rect 112346 86708 112352 86760
rect 112404 86748 112410 86760
rect 166442 86748 166448 86760
rect 112404 86720 166448 86748
rect 112404 86708 112410 86720
rect 166442 86708 166448 86720
rect 166500 86708 166506 86760
rect 124122 86640 124128 86692
rect 124180 86680 124186 86692
rect 170582 86680 170588 86692
rect 124180 86652 170588 86680
rect 124180 86640 124186 86652
rect 170582 86640 170588 86652
rect 170640 86640 170646 86692
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 44818 85524 44824 85536
rect 3200 85496 44824 85524
rect 3200 85484 3206 85496
rect 44818 85484 44824 85496
rect 44876 85484 44882 85536
rect 111610 85484 111616 85536
rect 111668 85524 111674 85536
rect 210602 85524 210608 85536
rect 111668 85496 210608 85524
rect 111668 85484 111674 85496
rect 210602 85484 210608 85496
rect 210660 85484 210666 85536
rect 66070 85416 66076 85468
rect 66128 85456 66134 85468
rect 164878 85456 164884 85468
rect 66128 85428 164884 85456
rect 66128 85416 66134 85428
rect 164878 85416 164884 85428
rect 164936 85416 164942 85468
rect 104342 85348 104348 85400
rect 104400 85388 104406 85400
rect 184198 85388 184204 85400
rect 104400 85360 184204 85388
rect 104400 85348 104406 85360
rect 184198 85348 184204 85360
rect 184256 85348 184262 85400
rect 100570 85280 100576 85332
rect 100628 85320 100634 85332
rect 170674 85320 170680 85332
rect 100628 85292 170680 85320
rect 100628 85280 100634 85292
rect 170674 85280 170680 85292
rect 170732 85280 170738 85332
rect 122834 85212 122840 85264
rect 122892 85252 122898 85264
rect 173342 85252 173348 85264
rect 122892 85224 173348 85252
rect 122892 85212 122898 85224
rect 173342 85212 173348 85224
rect 173400 85212 173406 85264
rect 132034 85144 132040 85196
rect 132092 85184 132098 85196
rect 176010 85184 176016 85196
rect 132092 85156 176016 85184
rect 132092 85144 132098 85156
rect 176010 85144 176016 85156
rect 176068 85144 176074 85196
rect 63402 84124 63408 84176
rect 63460 84164 63466 84176
rect 216030 84164 216036 84176
rect 63460 84136 216036 84164
rect 63460 84124 63466 84136
rect 216030 84124 216036 84136
rect 216088 84124 216094 84176
rect 107470 84056 107476 84108
rect 107528 84096 107534 84108
rect 211982 84096 211988 84108
rect 107528 84068 211988 84096
rect 107528 84056 107534 84068
rect 211982 84056 211988 84068
rect 212040 84056 212046 84108
rect 101858 83988 101864 84040
rect 101916 84028 101922 84040
rect 197998 84028 198004 84040
rect 101916 84000 198004 84028
rect 101916 83988 101922 84000
rect 197998 83988 198004 84000
rect 198056 83988 198062 84040
rect 118602 83920 118608 83972
rect 118660 83960 118666 83972
rect 180242 83960 180248 83972
rect 118660 83932 180248 83960
rect 118660 83920 118666 83932
rect 180242 83920 180248 83932
rect 180300 83920 180306 83972
rect 67450 82764 67456 82816
rect 67508 82804 67514 82816
rect 204898 82804 204904 82816
rect 67508 82776 204904 82804
rect 67508 82764 67514 82776
rect 204898 82764 204904 82776
rect 204956 82764 204962 82816
rect 99098 82696 99104 82748
rect 99156 82736 99162 82748
rect 202230 82736 202236 82748
rect 99156 82708 202236 82736
rect 99156 82696 99162 82708
rect 202230 82696 202236 82708
rect 202288 82696 202294 82748
rect 110322 82628 110328 82680
rect 110380 82668 110386 82680
rect 213178 82668 213184 82680
rect 110380 82640 213184 82668
rect 110380 82628 110386 82640
rect 213178 82628 213184 82640
rect 213236 82628 213242 82680
rect 121362 82560 121368 82612
rect 121420 82600 121426 82612
rect 174722 82600 174728 82612
rect 121420 82572 174728 82600
rect 121420 82560 121426 82572
rect 174722 82560 174728 82572
rect 174780 82560 174786 82612
rect 126882 82492 126888 82544
rect 126940 82532 126946 82544
rect 169018 82532 169024 82544
rect 126940 82504 169024 82532
rect 126940 82492 126946 82504
rect 169018 82492 169024 82504
rect 169076 82492 169082 82544
rect 108298 81336 108304 81388
rect 108356 81376 108362 81388
rect 214650 81376 214656 81388
rect 108356 81348 214656 81376
rect 108356 81336 108362 81348
rect 214650 81336 214656 81348
rect 214708 81336 214714 81388
rect 97810 81268 97816 81320
rect 97868 81308 97874 81320
rect 178770 81308 178776 81320
rect 97868 81280 178776 81308
rect 97868 81268 97874 81280
rect 178770 81268 178776 81280
rect 178828 81268 178834 81320
rect 86862 81200 86868 81252
rect 86920 81240 86926 81252
rect 167822 81240 167828 81252
rect 86920 81212 167828 81240
rect 86920 81200 86926 81212
rect 167822 81200 167828 81212
rect 167880 81200 167886 81252
rect 93762 81132 93768 81184
rect 93820 81172 93826 81184
rect 167730 81172 167736 81184
rect 93820 81144 167736 81172
rect 93820 81132 93826 81144
rect 167730 81132 167736 81144
rect 167788 81132 167794 81184
rect 125410 81064 125416 81116
rect 125468 81104 125474 81116
rect 193858 81104 193864 81116
rect 125468 81076 193864 81104
rect 125468 81064 125474 81076
rect 193858 81064 193864 81076
rect 193916 81064 193922 81116
rect 67542 79976 67548 80028
rect 67600 80016 67606 80028
rect 207842 80016 207848 80028
rect 67600 79988 207848 80016
rect 67600 79976 67606 79988
rect 207842 79976 207848 79988
rect 207900 79976 207906 80028
rect 114462 79908 114468 79960
rect 114520 79948 114526 79960
rect 210510 79948 210516 79960
rect 114520 79920 210516 79948
rect 114520 79908 114526 79920
rect 210510 79908 210516 79920
rect 210568 79908 210574 79960
rect 103422 79840 103428 79892
rect 103480 79880 103486 79892
rect 189718 79880 189724 79892
rect 103480 79852 189724 79880
rect 103480 79840 103486 79852
rect 189718 79840 189724 79852
rect 189776 79840 189782 79892
rect 95050 79772 95056 79824
rect 95108 79812 95114 79824
rect 174814 79812 174820 79824
rect 95108 79784 174820 79812
rect 95108 79772 95114 79784
rect 174814 79772 174820 79784
rect 174872 79772 174878 79824
rect 97902 78616 97908 78668
rect 97960 78656 97966 78668
rect 206370 78656 206376 78668
rect 97960 78628 206376 78656
rect 97960 78616 97966 78628
rect 206370 78616 206376 78628
rect 206428 78616 206434 78668
rect 122742 78548 122748 78600
rect 122800 78588 122806 78600
rect 211798 78588 211804 78600
rect 122800 78560 211804 78588
rect 122800 78548 122806 78560
rect 211798 78548 211804 78560
rect 211856 78548 211862 78600
rect 99282 78480 99288 78532
rect 99340 78520 99346 78532
rect 177298 78520 177304 78532
rect 99340 78492 177304 78520
rect 99340 78480 99346 78492
rect 177298 78480 177304 78492
rect 177356 78480 177362 78532
rect 99190 78412 99196 78464
rect 99248 78452 99254 78464
rect 173250 78452 173256 78464
rect 99248 78424 173256 78452
rect 99248 78412 99254 78424
rect 173250 78412 173256 78424
rect 173308 78412 173314 78464
rect 85482 77188 85488 77240
rect 85540 77228 85546 77240
rect 172054 77228 172060 77240
rect 85540 77200 172060 77228
rect 85540 77188 85546 77200
rect 172054 77188 172060 77200
rect 172112 77188 172118 77240
rect 77294 76576 77300 76628
rect 77352 76616 77358 76628
rect 290642 76616 290648 76628
rect 77352 76588 290648 76616
rect 77352 76576 77358 76588
rect 290642 76576 290648 76588
rect 290700 76576 290706 76628
rect 89714 76508 89720 76560
rect 89772 76548 89778 76560
rect 306006 76548 306012 76560
rect 89772 76520 306012 76548
rect 89772 76508 89778 76520
rect 306006 76508 306012 76520
rect 306064 76508 306070 76560
rect 95142 75828 95148 75880
rect 95200 75868 95206 75880
rect 203610 75868 203616 75880
rect 95200 75840 203616 75868
rect 95200 75828 95206 75840
rect 203610 75828 203616 75840
rect 203668 75828 203674 75880
rect 102042 75760 102048 75812
rect 102100 75800 102106 75812
rect 177390 75800 177396 75812
rect 102100 75772 177396 75800
rect 102100 75760 102106 75772
rect 177390 75760 177396 75772
rect 177448 75760 177454 75812
rect 107654 75148 107660 75200
rect 107712 75188 107718 75200
rect 303154 75188 303160 75200
rect 107712 75160 303160 75188
rect 107712 75148 107718 75160
rect 303154 75148 303160 75160
rect 303212 75148 303218 75200
rect 103514 73856 103520 73908
rect 103572 73896 103578 73908
rect 304534 73896 304540 73908
rect 103572 73868 304540 73896
rect 103572 73856 103578 73868
rect 304534 73856 304540 73868
rect 304592 73856 304598 73908
rect 9674 73788 9680 73840
rect 9732 73828 9738 73840
rect 294690 73828 294696 73840
rect 9732 73800 294696 73828
rect 9732 73788 9738 73800
rect 294690 73788 294696 73800
rect 294748 73788 294754 73840
rect 122834 72496 122840 72548
rect 122892 72536 122898 72548
rect 289354 72536 289360 72548
rect 122892 72508 289360 72536
rect 122892 72496 122898 72508
rect 289354 72496 289360 72508
rect 289412 72496 289418 72548
rect 53834 72428 53840 72480
rect 53892 72468 53898 72480
rect 305822 72468 305828 72480
rect 53892 72440 305828 72468
rect 53892 72428 53898 72440
rect 305822 72428 305828 72440
rect 305880 72428 305886 72480
rect 62114 71068 62120 71120
rect 62172 71108 62178 71120
rect 293402 71108 293408 71120
rect 62172 71080 293408 71108
rect 62172 71068 62178 71080
rect 293402 71068 293408 71080
rect 293460 71068 293466 71120
rect 68278 71000 68284 71052
rect 68336 71040 68342 71052
rect 307202 71040 307208 71052
rect 68336 71012 307208 71040
rect 68336 71000 68342 71012
rect 307202 71000 307208 71012
rect 307260 71000 307266 71052
rect 66254 69640 66260 69692
rect 66312 69680 66318 69692
rect 299014 69680 299020 69692
rect 66312 69652 299020 69680
rect 66312 69640 66318 69652
rect 299014 69640 299020 69652
rect 299072 69640 299078 69692
rect 57974 68348 57980 68400
rect 58032 68388 58038 68400
rect 287974 68388 287980 68400
rect 58032 68360 287980 68388
rect 58032 68348 58038 68360
rect 287974 68348 287980 68360
rect 288032 68348 288038 68400
rect 20714 68280 20720 68332
rect 20772 68320 20778 68332
rect 304626 68320 304632 68332
rect 20772 68292 304632 68320
rect 20772 68280 20778 68292
rect 304626 68280 304632 68292
rect 304684 68280 304690 68332
rect 71774 66920 71780 66972
rect 71832 66960 71838 66972
rect 269850 66960 269856 66972
rect 71832 66932 269856 66960
rect 71832 66920 71838 66932
rect 269850 66920 269856 66932
rect 269908 66920 269914 66972
rect 26234 66852 26240 66904
rect 26292 66892 26298 66904
rect 293586 66892 293592 66904
rect 26292 66864 293592 66892
rect 26292 66852 26298 66864
rect 293586 66852 293592 66864
rect 293644 66852 293650 66904
rect 82814 65492 82820 65544
rect 82872 65532 82878 65544
rect 282362 65532 282368 65544
rect 82872 65504 282368 65532
rect 82872 65492 82878 65504
rect 282362 65492 282368 65504
rect 282420 65492 282426 65544
rect 33134 64132 33140 64184
rect 33192 64172 33198 64184
rect 286410 64172 286416 64184
rect 33192 64144 286416 64172
rect 33192 64132 33198 64144
rect 286410 64132 286416 64144
rect 286468 64132 286474 64184
rect 80054 62840 80060 62892
rect 80112 62880 80118 62892
rect 266998 62880 267004 62892
rect 80112 62852 267004 62880
rect 80112 62840 80118 62852
rect 266998 62840 267004 62852
rect 267056 62840 267062 62892
rect 35894 62772 35900 62824
rect 35952 62812 35958 62824
rect 303062 62812 303068 62824
rect 35952 62784 303068 62812
rect 35952 62772 35958 62784
rect 303062 62772 303068 62784
rect 303120 62772 303126 62824
rect 93854 61344 93860 61396
rect 93912 61384 93918 61396
rect 268378 61384 268384 61396
rect 93912 61356 268384 61384
rect 93912 61344 93918 61356
rect 268378 61344 268384 61356
rect 268436 61344 268442 61396
rect 175918 60664 175924 60716
rect 175976 60704 175982 60716
rect 580166 60704 580172 60716
rect 175976 60676 580172 60704
rect 175976 60664 175982 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 118694 59984 118700 60036
rect 118752 60024 118758 60036
rect 300302 60024 300308 60036
rect 118752 59996 300308 60024
rect 118752 59984 118758 59996
rect 300302 59984 300308 59996
rect 300360 59984 300366 60036
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 48958 59344 48964 59356
rect 3108 59316 48964 59344
rect 3108 59304 3114 59316
rect 48958 59304 48964 59316
rect 49016 59304 49022 59356
rect 110414 58692 110420 58744
rect 110472 58732 110478 58744
rect 301774 58732 301780 58744
rect 110472 58704 301780 58732
rect 110472 58692 110478 58704
rect 301774 58692 301780 58704
rect 301832 58692 301838 58744
rect 48314 58624 48320 58676
rect 48372 58664 48378 58676
rect 292022 58664 292028 58676
rect 48372 58636 292028 58664
rect 48372 58624 48378 58636
rect 292022 58624 292028 58636
rect 292080 58624 292086 58676
rect 81434 57196 81440 57248
rect 81492 57236 81498 57248
rect 283742 57236 283748 57248
rect 81492 57208 283748 57236
rect 81492 57196 81498 57208
rect 283742 57196 283748 57208
rect 283800 57196 283806 57248
rect 40034 55904 40040 55956
rect 40092 55944 40098 55956
rect 257338 55944 257344 55956
rect 40092 55916 257344 55944
rect 40092 55904 40098 55916
rect 257338 55904 257344 55916
rect 257396 55904 257402 55956
rect 55214 55836 55220 55888
rect 55272 55876 55278 55888
rect 300394 55876 300400 55888
rect 55272 55848 300400 55876
rect 55272 55836 55278 55848
rect 300394 55836 300400 55848
rect 300452 55836 300458 55888
rect 92474 54544 92480 54596
rect 92532 54584 92538 54596
rect 271230 54584 271236 54596
rect 92532 54556 271236 54584
rect 92532 54544 92538 54556
rect 271230 54544 271236 54556
rect 271288 54544 271294 54596
rect 15194 54476 15200 54528
rect 15252 54516 15258 54528
rect 292114 54516 292120 54528
rect 15252 54488 292120 54516
rect 15252 54476 15258 54488
rect 292114 54476 292120 54488
rect 292172 54476 292178 54528
rect 99374 53116 99380 53168
rect 99432 53156 99438 53168
rect 284938 53156 284944 53168
rect 99432 53128 284944 53156
rect 99432 53116 99438 53128
rect 284938 53116 284944 53128
rect 284996 53116 285002 53168
rect 24854 53048 24860 53100
rect 24912 53088 24918 53100
rect 294782 53088 294788 53100
rect 24912 53060 294788 53088
rect 24912 53048 24918 53060
rect 294782 53048 294788 53060
rect 294840 53048 294846 53100
rect 12434 51688 12440 51740
rect 12492 51728 12498 51740
rect 279602 51728 279608 51740
rect 12492 51700 279608 51728
rect 12492 51688 12498 51700
rect 279602 51688 279608 51700
rect 279660 51688 279666 51740
rect 84194 50396 84200 50448
rect 84252 50436 84258 50448
rect 287882 50436 287888 50448
rect 84252 50408 287888 50436
rect 84252 50396 84258 50408
rect 287882 50396 287888 50408
rect 287940 50396 287946 50448
rect 27614 50328 27620 50380
rect 27672 50368 27678 50380
rect 272518 50368 272524 50380
rect 27672 50340 272524 50368
rect 27672 50328 27678 50340
rect 272518 50328 272524 50340
rect 272576 50328 272582 50380
rect 86954 49036 86960 49088
rect 87012 49076 87018 49088
rect 297542 49076 297548 49088
rect 87012 49048 297548 49076
rect 87012 49036 87018 49048
rect 297542 49036 297548 49048
rect 297600 49036 297606 49088
rect 23474 48968 23480 49020
rect 23532 49008 23538 49020
rect 285030 49008 285036 49020
rect 23532 48980 285036 49008
rect 23532 48968 23538 48980
rect 285030 48968 285036 48980
rect 285088 48968 285094 49020
rect 88334 47608 88340 47660
rect 88392 47648 88398 47660
rect 302878 47648 302884 47660
rect 88392 47620 302884 47648
rect 88392 47608 88398 47620
rect 302878 47608 302884 47620
rect 302936 47608 302942 47660
rect 17954 47540 17960 47592
rect 18012 47580 18018 47592
rect 291930 47580 291936 47592
rect 18012 47552 291936 47580
rect 18012 47540 18018 47552
rect 291930 47540 291936 47552
rect 291988 47540 291994 47592
rect 106274 46180 106280 46232
rect 106332 46220 106338 46232
rect 282270 46220 282276 46232
rect 106332 46192 282276 46220
rect 106332 46180 106338 46192
rect 282270 46180 282276 46192
rect 282328 46180 282334 46232
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 43438 45540 43444 45552
rect 3476 45512 43444 45540
rect 3476 45500 3482 45512
rect 43438 45500 43444 45512
rect 43496 45500 43502 45552
rect 102134 44888 102140 44940
rect 102192 44928 102198 44940
rect 302970 44928 302976 44940
rect 102192 44900 302976 44928
rect 102192 44888 102198 44900
rect 302970 44888 302976 44900
rect 303028 44888 303034 44940
rect 63494 44820 63500 44872
rect 63552 44860 63558 44872
rect 279510 44860 279516 44872
rect 63552 44832 279516 44860
rect 63552 44820 63558 44832
rect 279510 44820 279516 44832
rect 279568 44820 279574 44872
rect 56594 43392 56600 43444
rect 56652 43432 56658 43444
rect 291838 43432 291844 43444
rect 56652 43404 291844 43432
rect 56652 43392 56658 43404
rect 291838 43392 291844 43404
rect 291896 43392 291902 43444
rect 85574 42100 85580 42152
rect 85632 42140 85638 42152
rect 275278 42140 275284 42152
rect 85632 42112 275284 42140
rect 85632 42100 85638 42112
rect 275278 42100 275284 42112
rect 275336 42100 275342 42152
rect 97994 42032 98000 42084
rect 98052 42072 98058 42084
rect 300210 42072 300216 42084
rect 98052 42044 300216 42072
rect 98052 42032 98058 42044
rect 300210 42032 300216 42044
rect 300268 42032 300274 42084
rect 91094 40740 91100 40792
rect 91152 40780 91158 40792
rect 293310 40780 293316 40792
rect 91152 40752 293316 40780
rect 91152 40740 91158 40752
rect 293310 40740 293316 40752
rect 293368 40740 293374 40792
rect 19334 40672 19340 40724
rect 19392 40712 19398 40724
rect 295978 40712 295984 40724
rect 19392 40684 295984 40712
rect 19392 40672 19398 40684
rect 295978 40672 295984 40684
rect 296036 40672 296042 40724
rect 95234 39380 95240 39432
rect 95292 39420 95298 39432
rect 297358 39420 297364 39432
rect 95292 39392 297364 39420
rect 95292 39380 95298 39392
rect 297358 39380 297364 39392
rect 297416 39380 297422 39432
rect 31754 39312 31760 39364
rect 31812 39352 31818 39364
rect 294598 39352 294604 39364
rect 31812 39324 294604 39352
rect 31812 39312 31818 39324
rect 294598 39312 294604 39324
rect 294656 39312 294662 39364
rect 77386 37952 77392 38004
rect 77444 37992 77450 38004
rect 301682 37992 301688 38004
rect 77444 37964 301688 37992
rect 77444 37952 77450 37964
rect 301682 37952 301688 37964
rect 301740 37952 301746 38004
rect 38654 37884 38660 37936
rect 38712 37924 38718 37936
rect 265618 37924 265624 37936
rect 38712 37896 265624 37924
rect 38712 37884 38718 37896
rect 265618 37884 265624 37896
rect 265676 37884 265682 37936
rect 73154 36592 73160 36644
rect 73212 36632 73218 36644
rect 296162 36632 296168 36644
rect 73212 36604 296168 36632
rect 73212 36592 73218 36604
rect 296162 36592 296168 36604
rect 296220 36592 296226 36644
rect 42794 36524 42800 36576
rect 42852 36564 42858 36576
rect 276658 36564 276664 36576
rect 42852 36536 276664 36564
rect 42852 36524 42858 36536
rect 276658 36524 276664 36536
rect 276716 36524 276722 36576
rect 69014 35232 69020 35284
rect 69072 35272 69078 35284
rect 305730 35272 305736 35284
rect 69072 35244 305736 35272
rect 69072 35232 69078 35244
rect 305730 35232 305736 35244
rect 305788 35232 305794 35284
rect 16574 35164 16580 35216
rect 16632 35204 16638 35216
rect 289262 35204 289268 35216
rect 16632 35176 289268 35204
rect 16632 35164 16638 35176
rect 289262 35164 289268 35176
rect 289320 35164 289326 35216
rect 113174 33804 113180 33856
rect 113232 33844 113238 33856
rect 298738 33844 298744 33856
rect 113232 33816 298744 33844
rect 113232 33804 113238 33816
rect 298738 33804 298744 33816
rect 298796 33804 298802 33856
rect 3234 33736 3240 33788
rect 3292 33776 3298 33788
rect 46198 33776 46204 33788
rect 3292 33748 46204 33776
rect 3292 33736 3298 33748
rect 46198 33736 46204 33748
rect 46256 33736 46262 33788
rect 52454 33736 52460 33788
rect 52512 33776 52518 33788
rect 296070 33776 296076 33788
rect 52512 33748 296076 33776
rect 52512 33736 52518 33748
rect 296070 33736 296076 33748
rect 296128 33736 296134 33788
rect 27706 32376 27712 32428
rect 27764 32416 27770 32428
rect 298830 32416 298836 32428
rect 27764 32388 298836 32416
rect 27764 32376 27770 32388
rect 298830 32376 298836 32388
rect 298888 32376 298894 32428
rect 85666 31084 85672 31136
rect 85724 31124 85730 31136
rect 304350 31124 304356 31136
rect 85724 31096 304356 31124
rect 85724 31084 85730 31096
rect 304350 31084 304356 31096
rect 304408 31084 304414 31136
rect 44174 31016 44180 31068
rect 44232 31056 44238 31068
rect 298922 31056 298928 31068
rect 44232 31028 298928 31056
rect 44232 31016 44238 31028
rect 298922 31016 298928 31028
rect 298980 31016 298986 31068
rect 118786 29656 118792 29708
rect 118844 29696 118850 29708
rect 297450 29696 297456 29708
rect 118844 29668 297456 29696
rect 118844 29656 118850 29668
rect 297450 29656 297456 29668
rect 297508 29656 297514 29708
rect 37274 29588 37280 29640
rect 37332 29628 37338 29640
rect 264330 29628 264336 29640
rect 37332 29600 264336 29628
rect 37332 29588 37338 29600
rect 264330 29588 264336 29600
rect 264388 29588 264394 29640
rect 114554 28296 114560 28348
rect 114612 28336 114618 28348
rect 296254 28336 296260 28348
rect 114612 28308 296260 28336
rect 114612 28296 114618 28308
rect 296254 28296 296260 28308
rect 296312 28296 296318 28348
rect 44266 28228 44272 28280
rect 44324 28268 44330 28280
rect 265710 28268 265716 28280
rect 44324 28240 265716 28268
rect 44324 28228 44330 28240
rect 265710 28228 265716 28240
rect 265768 28228 265774 28280
rect 121454 26936 121460 26988
rect 121512 26976 121518 26988
rect 300118 26976 300124 26988
rect 121512 26948 300124 26976
rect 121512 26936 121518 26948
rect 300118 26936 300124 26948
rect 300176 26936 300182 26988
rect 52546 26868 52552 26920
rect 52604 26908 52610 26920
rect 290550 26908 290556 26920
rect 52604 26880 290556 26908
rect 52604 26868 52610 26880
rect 290550 26868 290556 26880
rect 290608 26868 290614 26920
rect 100754 25576 100760 25628
rect 100812 25616 100818 25628
rect 278222 25616 278228 25628
rect 100812 25588 278228 25616
rect 100812 25576 100818 25588
rect 278222 25576 278228 25588
rect 278280 25576 278286 25628
rect 60734 25508 60740 25560
rect 60792 25548 60798 25560
rect 287790 25548 287796 25560
rect 60792 25520 287796 25548
rect 60792 25508 60798 25520
rect 287790 25508 287796 25520
rect 287848 25508 287854 25560
rect 93946 24148 93952 24200
rect 94004 24188 94010 24200
rect 301590 24188 301596 24200
rect 94004 24160 301596 24188
rect 94004 24148 94010 24160
rect 301590 24148 301596 24160
rect 301648 24148 301654 24200
rect 13814 24080 13820 24132
rect 13872 24120 13878 24132
rect 271138 24120 271144 24132
rect 13872 24092 271144 24120
rect 13872 24080 13878 24092
rect 271138 24080 271144 24092
rect 271196 24080 271202 24132
rect 75914 22720 75920 22772
rect 75972 22760 75978 22772
rect 283650 22760 283656 22772
rect 75972 22732 283656 22760
rect 75972 22720 75978 22732
rect 283650 22720 283656 22732
rect 283708 22720 283714 22772
rect 78674 21428 78680 21480
rect 78732 21468 78738 21480
rect 301498 21468 301504 21480
rect 78732 21440 301504 21468
rect 78732 21428 78738 21440
rect 301498 21428 301504 21440
rect 301556 21428 301562 21480
rect 35986 21360 35992 21412
rect 36044 21400 36050 21412
rect 273990 21400 273996 21412
rect 36044 21372 273996 21400
rect 36044 21360 36050 21372
rect 273990 21360 273996 21372
rect 274048 21360 274054 21412
rect 3510 20612 3516 20664
rect 3568 20652 3574 20664
rect 32398 20652 32404 20664
rect 3568 20624 32404 20652
rect 3568 20612 3574 20624
rect 32398 20612 32404 20624
rect 32456 20612 32462 20664
rect 3418 19932 3424 19984
rect 3476 19972 3482 19984
rect 57238 19972 57244 19984
rect 3476 19944 57244 19972
rect 3476 19932 3482 19944
rect 57238 19932 57244 19944
rect 57296 19932 57302 19984
rect 115934 19932 115940 19984
rect 115992 19972 115998 19984
rect 304258 19972 304264 19984
rect 115992 19944 304264 19972
rect 115992 19932 115998 19944
rect 304258 19932 304264 19944
rect 304316 19932 304322 19984
rect 69106 18640 69112 18692
rect 69164 18680 69170 18692
rect 289170 18680 289176 18692
rect 69164 18652 289176 18680
rect 69164 18640 69170 18652
rect 289170 18640 289176 18652
rect 289228 18640 289234 18692
rect 45554 18572 45560 18624
rect 45612 18612 45618 18624
rect 279418 18612 279424 18624
rect 45612 18584 279424 18612
rect 45612 18572 45618 18584
rect 279418 18572 279424 18584
rect 279476 18572 279482 18624
rect 64874 17280 64880 17332
rect 64932 17320 64938 17332
rect 305638 17320 305644 17332
rect 64932 17292 305644 17320
rect 64932 17280 64938 17292
rect 305638 17280 305644 17292
rect 305696 17280 305702 17332
rect 11146 17212 11152 17264
rect 11204 17252 11210 17264
rect 256050 17252 256056 17264
rect 11204 17224 256056 17252
rect 11204 17212 11210 17224
rect 256050 17212 256056 17224
rect 256108 17212 256114 17264
rect 61562 15920 61568 15972
rect 61620 15960 61626 15972
rect 280890 15960 280896 15972
rect 61620 15932 280896 15960
rect 61620 15920 61626 15932
rect 280890 15920 280896 15932
rect 280948 15920 280954 15972
rect 20162 15852 20168 15904
rect 20220 15892 20226 15904
rect 260098 15892 260104 15904
rect 20220 15864 260104 15892
rect 20220 15852 20226 15864
rect 260098 15852 260104 15864
rect 260156 15852 260162 15904
rect 105722 14424 105728 14476
rect 105780 14464 105786 14476
rect 283558 14464 283564 14476
rect 105780 14436 283564 14464
rect 105780 14424 105786 14436
rect 283558 14424 283564 14436
rect 283616 14424 283622 14476
rect 124674 13132 124680 13184
rect 124732 13172 124738 13184
rect 280798 13172 280804 13184
rect 124732 13144 280804 13172
rect 124732 13132 124738 13144
rect 280798 13132 280804 13144
rect 280856 13132 280862 13184
rect 47394 13064 47400 13116
rect 47452 13104 47458 13116
rect 269758 13104 269764 13116
rect 47452 13076 269764 13104
rect 47452 13064 47458 13076
rect 269758 13064 269764 13076
rect 269816 13064 269822 13116
rect 117314 11772 117320 11824
rect 117372 11812 117378 11824
rect 278130 11812 278136 11824
rect 117372 11784 278136 11812
rect 117372 11772 117378 11784
rect 278130 11772 278136 11784
rect 278188 11772 278194 11824
rect 7650 11704 7656 11756
rect 7708 11744 7714 11756
rect 286318 11744 286324 11756
rect 7708 11716 286324 11744
rect 7708 11704 7714 11716
rect 286318 11704 286324 11716
rect 286376 11704 286382 11756
rect 110506 10344 110512 10396
rect 110564 10384 110570 10396
rect 264238 10384 264244 10396
rect 110564 10356 264244 10384
rect 110564 10344 110570 10356
rect 264238 10344 264244 10356
rect 264296 10344 264302 10396
rect 2866 10276 2872 10328
rect 2924 10316 2930 10328
rect 289078 10316 289084 10328
rect 2924 10288 289084 10316
rect 2924 10276 2930 10288
rect 289078 10276 289084 10288
rect 289136 10276 289142 10328
rect 7466 9596 7472 9648
rect 7524 9636 7530 9648
rect 8202 9636 8208 9648
rect 7524 9608 8208 9636
rect 7524 9596 7530 9608
rect 8202 9596 8208 9608
rect 8260 9636 8266 9648
rect 251174 9636 251180 9648
rect 8260 9608 251180 9636
rect 8260 9596 8266 9608
rect 251174 9596 251180 9608
rect 251232 9596 251238 9648
rect 74994 8916 75000 8968
rect 75052 8956 75058 8968
rect 293218 8956 293224 8968
rect 75052 8928 293224 8956
rect 75052 8916 75058 8928
rect 293218 8916 293224 8928
rect 293276 8916 293282 8968
rect 1670 8304 1676 8356
rect 1728 8344 1734 8356
rect 7466 8344 7472 8356
rect 1728 8316 7472 8344
rect 1728 8304 1734 8316
rect 7466 8304 7472 8316
rect 7524 8304 7530 8356
rect 63494 8236 63500 8288
rect 63552 8276 63558 8288
rect 64782 8276 64788 8288
rect 63552 8248 64788 8276
rect 63552 8236 63558 8248
rect 64782 8236 64788 8248
rect 64840 8276 64846 8288
rect 248414 8276 248420 8288
rect 64840 8248 248420 8276
rect 64840 8236 64846 8248
rect 248414 8236 248420 8248
rect 248472 8236 248478 8288
rect 566 7556 572 7608
rect 624 7596 630 7608
rect 63494 7596 63500 7608
rect 624 7568 63500 7596
rect 624 7556 630 7568
rect 63494 7556 63500 7568
rect 63552 7556 63558 7608
rect 71498 7556 71504 7608
rect 71556 7596 71562 7608
rect 287698 7596 287704 7608
rect 71556 7568 287704 7596
rect 71556 7556 71562 7568
rect 287698 7556 287704 7568
rect 287756 7556 287762 7608
rect 31294 6128 31300 6180
rect 31352 6168 31358 6180
rect 282178 6168 282184 6180
rect 31352 6140 282184 6168
rect 31352 6128 31358 6140
rect 282178 6128 282184 6140
rect 282236 6128 282242 6180
rect 97442 4836 97448 4888
rect 97500 4876 97506 4888
rect 261478 4876 261484 4888
rect 97500 4848 261484 4876
rect 97500 4836 97506 4848
rect 261478 4836 261484 4848
rect 261536 4836 261542 4888
rect 6454 4768 6460 4820
rect 6512 4808 6518 4820
rect 307018 4808 307024 4820
rect 6512 4780 307024 4808
rect 6512 4768 6518 4780
rect 307018 4768 307024 4780
rect 307076 4768 307082 4820
rect 235810 3952 235816 4004
rect 235868 3992 235874 4004
rect 239398 3992 239404 4004
rect 235868 3964 239404 3992
rect 235868 3952 235874 3964
rect 239398 3952 239404 3964
rect 239456 3952 239462 4004
rect 103486 3692 112576 3720
rect 41874 3544 41880 3596
rect 41932 3584 41938 3596
rect 68278 3584 68284 3596
rect 41932 3556 68284 3584
rect 41932 3544 41938 3556
rect 68278 3544 68284 3556
rect 68336 3544 68342 3596
rect 68388 3556 74534 3584
rect 2774 3476 2780 3528
rect 2832 3516 2838 3528
rect 3694 3516 3700 3528
rect 2832 3488 3700 3516
rect 2832 3476 2838 3488
rect 3694 3476 3700 3488
rect 3752 3476 3758 3528
rect 11054 3476 11060 3528
rect 11112 3516 11118 3528
rect 11974 3516 11980 3528
rect 11112 3488 11980 3516
rect 11112 3476 11118 3488
rect 11974 3476 11980 3488
rect 12032 3476 12038 3528
rect 27614 3476 27620 3528
rect 27672 3516 27678 3528
rect 28534 3516 28540 3528
rect 27672 3488 28540 3516
rect 27672 3476 27678 3488
rect 28534 3476 28540 3488
rect 28592 3476 28598 3528
rect 35894 3476 35900 3528
rect 35952 3516 35958 3528
rect 36814 3516 36820 3528
rect 35952 3488 36820 3516
rect 35952 3476 35958 3488
rect 36814 3476 36820 3488
rect 36872 3476 36878 3528
rect 67910 3476 67916 3528
rect 67968 3516 67974 3528
rect 68388 3516 68416 3556
rect 67968 3488 68416 3516
rect 67968 3476 67974 3488
rect 69014 3476 69020 3528
rect 69072 3516 69078 3528
rect 69934 3516 69940 3528
rect 69072 3488 69940 3516
rect 69072 3476 69078 3488
rect 69934 3476 69940 3488
rect 69992 3476 69998 3528
rect 74506 3516 74534 3556
rect 77294 3544 77300 3596
rect 77352 3584 77358 3596
rect 78214 3584 78220 3596
rect 77352 3556 78220 3584
rect 77352 3544 77358 3556
rect 78214 3544 78220 3556
rect 78272 3544 78278 3596
rect 93854 3544 93860 3596
rect 93912 3584 93918 3596
rect 94774 3584 94780 3596
rect 93912 3556 94780 3584
rect 93912 3544 93918 3556
rect 94774 3544 94780 3556
rect 94832 3544 94838 3596
rect 103330 3544 103336 3596
rect 103388 3584 103394 3596
rect 103486 3584 103514 3692
rect 112438 3584 112444 3596
rect 103388 3556 103514 3584
rect 108040 3556 112444 3584
rect 103388 3544 103394 3556
rect 108040 3516 108068 3556
rect 112438 3544 112444 3556
rect 112496 3544 112502 3596
rect 112548 3584 112576 3692
rect 112806 3612 112812 3664
rect 112864 3652 112870 3664
rect 180058 3652 180064 3664
rect 112864 3624 180064 3652
rect 112864 3612 112870 3624
rect 180058 3612 180064 3624
rect 180116 3612 180122 3664
rect 207658 3584 207664 3596
rect 112548 3556 207664 3584
rect 207658 3544 207664 3556
rect 207716 3544 207722 3596
rect 74506 3488 108068 3516
rect 110414 3476 110420 3528
rect 110472 3516 110478 3528
rect 111610 3516 111616 3528
rect 110472 3488 111616 3516
rect 110472 3476 110478 3488
rect 111610 3476 111616 3488
rect 111668 3476 111674 3528
rect 118694 3476 118700 3528
rect 118752 3516 118758 3528
rect 119890 3516 119896 3528
rect 118752 3488 119896 3516
rect 118752 3476 118758 3488
rect 119890 3476 119896 3488
rect 119948 3476 119954 3528
rect 121086 3476 121092 3528
rect 121144 3516 121150 3528
rect 273898 3516 273904 3528
rect 121144 3488 273904 3516
rect 121144 3476 121150 3488
rect 273898 3476 273904 3488
rect 273956 3476 273962 3528
rect 51350 3408 51356 3460
rect 51408 3448 51414 3460
rect 253198 3448 253204 3460
rect 51408 3420 253204 3448
rect 51408 3408 51414 3420
rect 253198 3408 253204 3420
rect 253256 3408 253262 3460
rect 109310 2116 109316 2168
rect 109368 2156 109374 2168
rect 290458 2156 290464 2168
rect 109368 2128 290464 2156
rect 109368 2116 109374 2128
rect 290458 2116 290464 2128
rect 290516 2116 290522 2168
rect 5258 2048 5264 2100
rect 5316 2088 5322 2100
rect 250438 2088 250444 2100
rect 5316 2060 250444 2088
rect 5316 2048 5322 2060
rect 250438 2048 250444 2060
rect 250496 2048 250502 2100
<< via1 >>
rect 201500 703060 201552 703112
rect 202788 703060 202840 703112
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 84292 702992 84344 703044
rect 348792 702992 348844 703044
rect 107660 702924 107712 702976
rect 413652 702924 413704 702976
rect 129004 702856 129056 702908
rect 462320 702856 462372 702908
rect 49608 702788 49660 702840
rect 397460 702788 397512 702840
rect 63408 702720 63460 702772
rect 429844 702720 429896 702772
rect 106280 702652 106332 702704
rect 478512 702652 478564 702704
rect 124864 702584 124916 702636
rect 527180 702584 527232 702636
rect 134524 702516 134576 702568
rect 559656 702516 559708 702568
rect 80704 702448 80756 702500
rect 580908 702448 580960 702500
rect 55128 700408 55180 700460
rect 105452 700408 105504 700460
rect 149704 700408 149756 700460
rect 235172 700408 235224 700460
rect 57888 700340 57940 700392
rect 170312 700340 170364 700392
rect 269764 700340 269816 700392
rect 332508 700340 332560 700392
rect 8116 700272 8168 700324
rect 8944 700272 8996 700324
rect 24308 700272 24360 700324
rect 82084 700272 82136 700324
rect 135904 700272 135956 700324
rect 364984 700272 365036 700324
rect 214564 699660 214616 699712
rect 218980 699660 219032 699712
rect 264244 699660 264296 699712
rect 267648 699660 267700 699712
rect 59268 697552 59320 697604
rect 137836 697552 137888 697604
rect 53748 696192 53800 696244
rect 300124 696192 300176 696244
rect 144184 683136 144236 683188
rect 580172 683136 580224 683188
rect 3516 670692 3568 670744
rect 26884 670692 26936 670744
rect 148324 670692 148376 670744
rect 580172 670692 580224 670744
rect 3516 656888 3568 656940
rect 39304 656888 39356 656940
rect 3516 632068 3568 632120
rect 21364 632068 21416 632120
rect 126244 630640 126296 630692
rect 580172 630640 580224 630692
rect 3516 618264 3568 618316
rect 46204 618264 46256 618316
rect 130384 616836 130436 616888
rect 580172 616836 580224 616888
rect 2780 605888 2832 605940
rect 4804 605888 4856 605940
rect 3332 579640 3384 579692
rect 116584 579640 116636 579692
rect 142804 576852 142856 576904
rect 580172 576852 580224 576904
rect 3240 565836 3292 565888
rect 64144 565836 64196 565888
rect 102784 563048 102836 563100
rect 579804 563048 579856 563100
rect 3332 553392 3384 553444
rect 18604 553392 18656 553444
rect 2964 527144 3016 527196
rect 36544 527144 36596 527196
rect 140044 524424 140096 524476
rect 580172 524424 580224 524476
rect 3332 500964 3384 501016
rect 100024 500964 100076 501016
rect 129096 484372 129148 484424
rect 580172 484372 580224 484424
rect 3056 474716 3108 474768
rect 111064 474716 111116 474768
rect 138664 470568 138716 470620
rect 580172 470568 580224 470620
rect 3332 462340 3384 462392
rect 31024 462340 31076 462392
rect 59176 456764 59228 456816
rect 580172 456764 580224 456816
rect 3332 448536 3384 448588
rect 25504 448536 25556 448588
rect 123484 430584 123536 430636
rect 579896 430584 579948 430636
rect 3332 423308 3384 423360
rect 7564 423308 7616 423360
rect 93124 418140 93176 418192
rect 580172 418140 580224 418192
rect 3332 409844 3384 409896
rect 17224 409844 17276 409896
rect 67548 404336 67600 404388
rect 580172 404336 580224 404388
rect 3332 397468 3384 397520
rect 43444 397468 43496 397520
rect 124956 378156 125008 378208
rect 580172 378156 580224 378208
rect 3332 371220 3384 371272
rect 50344 371220 50396 371272
rect 130476 364352 130528 364404
rect 579620 364352 579672 364404
rect 3332 357416 3384 357468
rect 13084 357416 13136 357468
rect 80796 351908 80848 351960
rect 580172 351908 580224 351960
rect 3332 345040 3384 345092
rect 117964 345040 118016 345092
rect 13084 338716 13136 338768
rect 98000 338716 98052 338768
rect 88340 334568 88392 334620
rect 103796 334568 103848 334620
rect 3424 326340 3476 326392
rect 120172 326340 120224 326392
rect 123576 324300 123628 324352
rect 580172 324300 580224 324352
rect 68928 323552 68980 323604
rect 269764 323552 269816 323604
rect 111064 322192 111116 322244
rect 121460 322192 121512 322244
rect 91100 319404 91152 319456
rect 148324 319404 148376 319456
rect 3332 318792 3384 318844
rect 22100 318792 22152 318844
rect 22100 318044 22152 318096
rect 115940 318044 115992 318096
rect 93952 317500 94004 317552
rect 102784 317500 102836 317552
rect 77300 315256 77352 315308
rect 93124 315256 93176 315308
rect 3516 313896 3568 313948
rect 120080 313896 120132 313948
rect 125140 313896 125192 313948
rect 282920 313896 282972 313948
rect 4804 312536 4856 312588
rect 94136 312536 94188 312588
rect 100024 312536 100076 312588
rect 121552 312536 121604 312588
rect 126336 311856 126388 311908
rect 580172 311856 580224 311908
rect 69112 311108 69164 311160
rect 153200 311108 153252 311160
rect 39304 309748 39356 309800
rect 121644 309748 121696 309800
rect 71780 308388 71832 308440
rect 114560 308388 114612 308440
rect 98092 307776 98144 307828
rect 283564 307776 283616 307828
rect 69020 307028 69072 307080
rect 580264 307028 580316 307080
rect 75920 306348 75972 306400
rect 342260 306348 342312 306400
rect 123668 305600 123720 305652
rect 201500 305600 201552 305652
rect 3424 305056 3476 305108
rect 119804 305056 119856 305108
rect 112444 304988 112496 305040
rect 281540 304988 281592 305040
rect 102140 303764 102192 303816
rect 185584 303764 185636 303816
rect 102416 303696 102468 303748
rect 224224 303696 224276 303748
rect 90272 303628 90324 303680
rect 278780 303628 278832 303680
rect 82084 303560 82136 303612
rect 84476 303560 84528 303612
rect 79232 302268 79284 302320
rect 189724 302268 189776 302320
rect 112168 302200 112220 302252
rect 273260 302200 273312 302252
rect 117964 301520 118016 301572
rect 119160 301520 119212 301572
rect 25504 301452 25556 301504
rect 70952 301452 71004 301504
rect 73528 301452 73580 301504
rect 80796 301452 80848 301504
rect 67456 300908 67508 300960
rect 152464 300908 152516 300960
rect 86408 300840 86460 300892
rect 319444 300840 319496 300892
rect 110420 299684 110472 299736
rect 184204 299684 184256 299736
rect 87696 299616 87748 299668
rect 225604 299616 225656 299668
rect 68744 299548 68796 299600
rect 308404 299548 308456 299600
rect 71780 299480 71832 299532
rect 343640 299480 343692 299532
rect 7564 298732 7616 298784
rect 72608 298732 72660 298784
rect 89996 298460 90048 298512
rect 166264 298460 166316 298512
rect 93216 298392 93268 298444
rect 174544 298392 174596 298444
rect 74540 298324 74592 298376
rect 192484 298324 192536 298376
rect 75184 298256 75236 298308
rect 274640 298256 274692 298308
rect 81624 298188 81676 298240
rect 333980 298188 334032 298240
rect 106096 298120 106148 298172
rect 582564 298120 582616 298172
rect 114468 297032 114520 297084
rect 160744 297032 160796 297084
rect 86132 296964 86184 297016
rect 210424 296964 210476 297016
rect 70032 296896 70084 296948
rect 248420 296896 248472 296948
rect 89352 296828 89404 296880
rect 339500 296828 339552 296880
rect 88708 296760 88760 296812
rect 340880 296760 340932 296812
rect 70676 296692 70728 296744
rect 325792 296692 325844 296744
rect 111248 295672 111300 295724
rect 157984 295672 158036 295724
rect 77116 295604 77168 295656
rect 126428 295604 126480 295656
rect 82268 295536 82320 295588
rect 178684 295536 178736 295588
rect 84200 295468 84252 295520
rect 196624 295468 196676 295520
rect 68560 295400 68612 295452
rect 278044 295400 278096 295452
rect 109960 295332 110012 295384
rect 347044 295332 347096 295384
rect 87420 294652 87472 294704
rect 112444 294652 112496 294704
rect 73252 294584 73304 294636
rect 111800 294584 111852 294636
rect 113824 294380 113876 294432
rect 118424 294380 118476 294432
rect 106740 294312 106792 294364
rect 170404 294312 170456 294364
rect 91928 294244 91980 294296
rect 215944 294244 215996 294296
rect 82912 294176 82964 294228
rect 255320 294176 255372 294228
rect 32404 294108 32456 294160
rect 69480 294040 69532 294092
rect 92572 294040 92624 294092
rect 117688 294108 117740 294160
rect 308496 294108 308548 294160
rect 118332 294040 118384 294092
rect 118424 294040 118476 294092
rect 345020 294040 345072 294092
rect 39304 293972 39356 294024
rect 77760 293972 77812 294024
rect 80704 293972 80756 294024
rect 84292 293972 84344 294024
rect 85212 293972 85264 294024
rect 93952 293972 94004 294024
rect 94780 293972 94832 294024
rect 111892 293972 111944 294024
rect 350540 293972 350592 294024
rect 78772 293904 78824 293956
rect 93860 292884 93912 292936
rect 120264 292884 120316 292936
rect 2780 292816 2832 292868
rect 4804 292816 4856 292868
rect 83556 292816 83608 292868
rect 220084 292816 220136 292868
rect 100944 292748 100996 292800
rect 263600 292748 263652 292800
rect 103520 292680 103572 292732
rect 318064 292680 318116 292732
rect 48964 292612 49016 292664
rect 97080 292612 97132 292664
rect 97724 292612 97776 292664
rect 320180 292612 320232 292664
rect 8208 292544 8260 292596
rect 96436 292544 96488 292596
rect 109316 292544 109368 292596
rect 336740 292544 336792 292596
rect 115848 291864 115900 291916
rect 117228 291864 117280 291916
rect 119068 291864 119120 291916
rect 119896 291864 119948 291916
rect 3424 291796 3476 291848
rect 69480 291796 69532 291848
rect 148324 291320 148376 291372
rect 345112 291252 345164 291304
rect 69756 291184 69808 291236
rect 582656 291184 582708 291236
rect 121644 289892 121696 289944
rect 246304 289892 246356 289944
rect 25504 289824 25556 289876
rect 67640 289824 67692 289876
rect 121736 289824 121788 289876
rect 269120 289824 269172 289876
rect 121644 289756 121696 289808
rect 124956 289756 125008 289808
rect 68560 289484 68612 289536
rect 68928 289484 68980 289536
rect 120264 289076 120316 289128
rect 202144 289076 202196 289128
rect 66076 288396 66128 288448
rect 68192 288396 68244 288448
rect 121644 288396 121696 288448
rect 313924 288396 313976 288448
rect 55036 287036 55088 287088
rect 67640 287036 67692 287088
rect 121644 286968 121696 287020
rect 123668 286968 123720 287020
rect 26884 286900 26936 286952
rect 67640 286900 67692 286952
rect 121828 286288 121880 286340
rect 327080 286288 327132 286340
rect 60648 285676 60700 285728
rect 67732 285676 67784 285728
rect 121552 285676 121604 285728
rect 193128 285676 193180 285728
rect 121644 285608 121696 285660
rect 138664 285608 138716 285660
rect 52368 284316 52420 284368
rect 67640 284316 67692 284368
rect 121552 284316 121604 284368
rect 335360 284316 335412 284368
rect 121552 284112 121604 284164
rect 124864 284112 124916 284164
rect 121552 282888 121604 282940
rect 307024 282888 307076 282940
rect 193128 282140 193180 282192
rect 580264 282140 580316 282192
rect 121552 281528 121604 281580
rect 242164 281528 242216 281580
rect 121552 280236 121604 280288
rect 238024 280236 238076 280288
rect 46848 280168 46900 280220
rect 67640 280168 67692 280220
rect 121644 280168 121696 280220
rect 342352 280168 342404 280220
rect 121552 278808 121604 278860
rect 206284 278808 206336 278860
rect 57244 278740 57296 278792
rect 67640 278740 67692 278792
rect 121644 278740 121696 278792
rect 318156 278740 318208 278792
rect 56508 277448 56560 277500
rect 67640 277448 67692 277500
rect 121644 277448 121696 277500
rect 328460 277448 328512 277500
rect 50896 277380 50948 277432
rect 67732 277380 67784 277432
rect 121552 277380 121604 277432
rect 347780 277380 347832 277432
rect 53656 276088 53708 276140
rect 67732 276088 67784 276140
rect 121644 276088 121696 276140
rect 247684 276088 247736 276140
rect 45468 276020 45520 276072
rect 67640 276020 67692 276072
rect 121552 276020 121604 276072
rect 331220 276020 331272 276072
rect 122196 275272 122248 275324
rect 392584 275272 392636 275324
rect 61936 274728 61988 274780
rect 67640 274728 67692 274780
rect 48228 274660 48280 274712
rect 67732 274660 67784 274712
rect 121552 274660 121604 274712
rect 253940 274660 253992 274712
rect 46204 274592 46256 274644
rect 67640 274592 67692 274644
rect 121644 274592 121696 274644
rect 126336 274592 126388 274644
rect 66168 273232 66220 273284
rect 68008 273232 68060 273284
rect 121552 273232 121604 273284
rect 211804 273232 211856 273284
rect 121644 273164 121696 273216
rect 126980 273164 127032 273216
rect 121736 272484 121788 272536
rect 395344 272484 395396 272536
rect 64512 271940 64564 271992
rect 67640 271940 67692 271992
rect 57704 271872 57756 271924
rect 67824 271872 67876 271924
rect 57888 271804 57940 271856
rect 67732 271804 67784 271856
rect 54944 270512 54996 270564
rect 67640 270512 67692 270564
rect 121552 270512 121604 270564
rect 249800 270512 249852 270564
rect 121644 269152 121696 269204
rect 207664 269152 207716 269204
rect 60556 269084 60608 269136
rect 67640 269084 67692 269136
rect 121552 269084 121604 269136
rect 239404 269084 239456 269136
rect 46204 267724 46256 267776
rect 67640 267724 67692 267776
rect 121552 267724 121604 267776
rect 311164 267724 311216 267776
rect 8944 267656 8996 267708
rect 67732 267656 67784 267708
rect 64144 267588 64196 267640
rect 67640 267588 67692 267640
rect 122104 266976 122156 267028
rect 255412 266976 255464 267028
rect 121460 266364 121512 266416
rect 345112 266364 345164 266416
rect 21364 266296 21416 266348
rect 67640 266296 67692 266348
rect 57796 265616 57848 265668
rect 68376 265616 68428 265668
rect 121460 265004 121512 265056
rect 308588 265004 308640 265056
rect 121552 264936 121604 264988
rect 349160 264936 349212 264988
rect 121460 264868 121512 264920
rect 129096 264868 129148 264920
rect 56416 263644 56468 263696
rect 67640 263644 67692 263696
rect 8944 263576 8996 263628
rect 67732 263576 67784 263628
rect 18604 263508 18656 263560
rect 67640 263508 67692 263560
rect 121460 262828 121512 262880
rect 254032 262828 254084 262880
rect 64604 262216 64656 262268
rect 67640 262216 67692 262268
rect 121460 262216 121512 262268
rect 327172 262216 327224 262268
rect 53472 260856 53524 260908
rect 67732 260856 67784 260908
rect 121460 260856 121512 260908
rect 342444 260856 342496 260908
rect 36544 260788 36596 260840
rect 67640 260788 67692 260840
rect 62028 259428 62080 259480
rect 67640 259428 67692 259480
rect 121460 259428 121512 259480
rect 267740 259428 267792 259480
rect 126428 259360 126480 259412
rect 579620 259360 579672 259412
rect 121460 259292 121512 259344
rect 149704 259292 149756 259344
rect 60464 258680 60516 258732
rect 67824 258680 67876 258732
rect 63316 258136 63368 258188
rect 67640 258136 67692 258188
rect 59084 258068 59136 258120
rect 67732 258068 67784 258120
rect 122196 257320 122248 257372
rect 332876 257320 332928 257372
rect 121460 257116 121512 257168
rect 123576 257116 123628 257168
rect 53564 256776 53616 256828
rect 67640 256776 67692 256828
rect 14464 256708 14516 256760
rect 67732 256708 67784 256760
rect 121644 256708 121696 256760
rect 232504 256708 232556 256760
rect 121552 256640 121604 256692
rect 130384 256640 130436 256692
rect 121460 256436 121512 256488
rect 123484 256436 123536 256488
rect 61752 255348 61804 255400
rect 67640 255348 67692 255400
rect 50988 255280 51040 255332
rect 67732 255280 67784 255332
rect 63408 255212 63460 255264
rect 67640 255212 67692 255264
rect 121460 253988 121512 254040
rect 198004 253988 198056 254040
rect 3148 253920 3200 253972
rect 13084 253920 13136 253972
rect 121552 253920 121604 253972
rect 323676 253920 323728 253972
rect 121644 253172 121696 253224
rect 144184 253172 144236 253224
rect 65892 252628 65944 252680
rect 68100 252628 68152 252680
rect 121552 252628 121604 252680
rect 233884 252628 233936 252680
rect 44824 252560 44876 252612
rect 67640 252560 67692 252612
rect 121460 252560 121512 252612
rect 347872 252560 347924 252612
rect 119804 251812 119856 251864
rect 142804 251812 142856 251864
rect 121460 251200 121512 251252
rect 346492 251200 346544 251252
rect 122104 250452 122156 250504
rect 331312 250452 331364 250504
rect 64696 249840 64748 249892
rect 67640 249840 67692 249892
rect 63132 249772 63184 249824
rect 67732 249772 67784 249824
rect 121552 249772 121604 249824
rect 203524 249772 203576 249824
rect 59268 249704 59320 249756
rect 67640 249704 67692 249756
rect 121460 249704 121512 249756
rect 140044 249704 140096 249756
rect 166264 249024 166316 249076
rect 305644 249024 305696 249076
rect 58992 248412 59044 248464
rect 67640 248412 67692 248464
rect 121460 248412 121512 248464
rect 309784 248412 309836 248464
rect 247684 247664 247736 247716
rect 580448 247664 580500 247716
rect 61844 247120 61896 247172
rect 67640 247120 67692 247172
rect 59268 247052 59320 247104
rect 67732 247052 67784 247104
rect 121460 247052 121512 247104
rect 229744 247052 229796 247104
rect 49608 246984 49660 247036
rect 67640 246984 67692 247036
rect 121552 245624 121604 245676
rect 270500 245624 270552 245676
rect 17224 245556 17276 245608
rect 67640 245556 67692 245608
rect 121460 245556 121512 245608
rect 129004 245556 129056 245608
rect 63408 244264 63460 244316
rect 67640 244264 67692 244316
rect 121552 244264 121604 244316
rect 323584 244264 323636 244316
rect 4804 244196 4856 244248
rect 67732 244196 67784 244248
rect 121460 243720 121512 243772
rect 125140 243720 125192 243772
rect 340972 243516 341024 243568
rect 579896 243516 579948 243568
rect 65984 242904 66036 242956
rect 67824 242904 67876 242956
rect 121552 242904 121604 242956
rect 311256 242904 311308 242956
rect 53748 242836 53800 242888
rect 67640 242836 67692 242888
rect 121460 242836 121512 242888
rect 340972 242836 341024 242888
rect 121552 242768 121604 242820
rect 134524 242768 134576 242820
rect 63224 241476 63276 241528
rect 67732 241476 67784 241528
rect 59176 241408 59228 241460
rect 67640 241408 67692 241460
rect 119804 240184 119856 240236
rect 121552 240184 121604 240236
rect 328552 240184 328604 240236
rect 3056 240116 3108 240168
rect 16580 240116 16632 240168
rect 65892 239912 65944 239964
rect 71044 239912 71096 239964
rect 118976 239912 119028 239964
rect 119896 240116 119948 240168
rect 330116 240116 330168 240168
rect 70584 239368 70636 239420
rect 86224 239368 86276 239420
rect 117044 238824 117096 238876
rect 126244 238824 126296 238876
rect 40040 238756 40092 238808
rect 95792 238756 95844 238808
rect 115112 238756 115164 238808
rect 582472 238756 582524 238808
rect 3516 238688 3568 238740
rect 86776 238688 86828 238740
rect 113824 238688 113876 238740
rect 494060 238688 494112 238740
rect 72608 238620 72660 238672
rect 130476 238620 130528 238672
rect 50344 238552 50396 238604
rect 99012 238552 99064 238604
rect 55128 238484 55180 238536
rect 89352 238484 89404 238536
rect 98368 238484 98420 238536
rect 135904 238552 135956 238604
rect 95148 238144 95200 238196
rect 106924 238144 106976 238196
rect 105452 238076 105504 238128
rect 188344 238076 188396 238128
rect 74540 238008 74592 238060
rect 338120 238008 338172 238060
rect 79048 237600 79100 237652
rect 80704 237600 80756 237652
rect 71320 237396 71372 237448
rect 75184 237396 75236 237448
rect 43444 237328 43496 237380
rect 82268 237328 82320 237380
rect 91928 237328 91980 237380
rect 582748 237328 582800 237380
rect 16580 237260 16632 237312
rect 103520 237260 103572 237312
rect 31024 237192 31076 237244
rect 114468 237192 114520 237244
rect 97724 236648 97776 236700
rect 340972 236648 341024 236700
rect 106740 235900 106792 235952
rect 264244 235900 264296 235952
rect 13084 235832 13136 235884
rect 112536 235832 112588 235884
rect 63408 235356 63460 235408
rect 280160 235356 280212 235408
rect 108028 235288 108080 235340
rect 327356 235288 327408 235340
rect 64788 235220 64840 235272
rect 121460 235220 121512 235272
rect 60464 233928 60516 233980
rect 192576 233928 192628 233980
rect 84292 233860 84344 233912
rect 85488 233860 85540 233912
rect 95240 233860 95292 233912
rect 96436 233860 96488 233912
rect 99380 233860 99432 233912
rect 100300 233860 100352 233912
rect 103612 233860 103664 233912
rect 104808 233860 104860 233912
rect 104900 233860 104952 233912
rect 106096 233860 106148 233912
rect 110420 233860 110472 233912
rect 111248 233860 111300 233912
rect 117688 233860 117740 233912
rect 582472 233860 582524 233912
rect 75828 233180 75880 233232
rect 582380 233180 582432 233232
rect 73160 232976 73212 233028
rect 73896 232976 73948 233028
rect 67364 232500 67416 232552
rect 324412 232500 324464 232552
rect 114560 232160 114612 232212
rect 115756 232160 115808 232212
rect 84108 231820 84160 231872
rect 84844 231820 84896 231872
rect 81624 231752 81676 231804
rect 214564 231752 214616 231804
rect 93216 231072 93268 231124
rect 331404 231072 331456 231124
rect 100760 231004 100812 231056
rect 101588 231004 101640 231056
rect 82912 229848 82964 229900
rect 175924 229848 175976 229900
rect 88064 229780 88116 229832
rect 252560 229780 252612 229832
rect 80060 229712 80112 229764
rect 80980 229712 81032 229764
rect 86132 229712 86184 229764
rect 582380 229712 582432 229764
rect 106832 229032 106884 229084
rect 542360 229032 542412 229084
rect 69112 228352 69164 228404
rect 321652 228352 321704 228404
rect 61752 227060 61804 227112
rect 276020 227060 276072 227112
rect 99656 226992 99708 227044
rect 343732 226992 343784 227044
rect 80336 225632 80388 225684
rect 315304 225632 315356 225684
rect 50896 225564 50948 225616
rect 309876 225564 309928 225616
rect 64512 224204 64564 224256
rect 214564 224204 214616 224256
rect 13084 223048 13136 223100
rect 110604 223048 110656 223100
rect 94504 222980 94556 223032
rect 287704 222980 287756 223032
rect 108672 222912 108724 222964
rect 329932 222912 329984 222964
rect 45468 222844 45520 222896
rect 312544 222844 312596 222896
rect 4804 221416 4856 221468
rect 83556 221416 83608 221468
rect 102876 221416 102928 221468
rect 252652 221416 252704 221468
rect 74908 220192 74960 220244
rect 254124 220192 254176 220244
rect 80704 220124 80756 220176
rect 263692 220124 263744 220176
rect 71044 220056 71096 220108
rect 334256 220056 334308 220108
rect 63224 218764 63276 218816
rect 228364 218764 228416 218816
rect 48228 218696 48280 218748
rect 346584 218696 346636 218748
rect 61936 217404 61988 217456
rect 262220 217404 262272 217456
rect 58992 217336 59044 217388
rect 277400 217336 277452 217388
rect 53472 217268 53524 217320
rect 318248 217268 318300 217320
rect 86224 215976 86276 216028
rect 314016 215976 314068 216028
rect 56416 215908 56468 215960
rect 291844 215908 291896 215960
rect 3516 214956 3568 215008
rect 8944 214956 8996 215008
rect 66076 214616 66128 214668
rect 251180 214616 251232 214668
rect 78680 214548 78732 214600
rect 330024 214548 330076 214600
rect 63316 213324 63368 213376
rect 224316 213324 224368 213376
rect 93860 213256 93912 213308
rect 278872 213256 278924 213308
rect 106924 213188 106976 213240
rect 341064 213188 341116 213240
rect 67548 211828 67600 211880
rect 251272 211828 251324 211880
rect 57704 211760 57756 211812
rect 271880 211760 271932 211812
rect 192576 210468 192628 210520
rect 307116 210468 307168 210520
rect 84292 210400 84344 210452
rect 249892 210400 249944 210452
rect 160744 209108 160796 209160
rect 300124 209108 300176 209160
rect 67456 209040 67508 209092
rect 324596 209040 324648 209092
rect 125048 206932 125100 206984
rect 580172 206932 580224 206984
rect 56508 206252 56560 206304
rect 266452 206252 266504 206304
rect 92480 204960 92532 205012
rect 252744 204960 252796 205012
rect 63132 204892 63184 204944
rect 242256 204892 242308 204944
rect 100852 203668 100904 203720
rect 270592 203668 270644 203720
rect 100760 203600 100812 203652
rect 274732 203600 274784 203652
rect 114560 203532 114612 203584
rect 327264 203532 327316 203584
rect 3056 202784 3108 202836
rect 120172 202784 120224 202836
rect 115940 202240 115992 202292
rect 266360 202240 266412 202292
rect 60556 202172 60608 202224
rect 271972 202172 272024 202224
rect 104900 202104 104952 202156
rect 339592 202104 339644 202156
rect 89812 200880 89864 200932
rect 254216 200880 254268 200932
rect 64604 200812 64656 200864
rect 260840 200812 260892 200864
rect 103704 200744 103756 200796
rect 321560 200744 321612 200796
rect 86960 199588 87012 199640
rect 196716 199588 196768 199640
rect 99380 199520 99432 199572
rect 249984 199520 250036 199572
rect 148324 199452 148376 199504
rect 334164 199452 334216 199504
rect 59268 199384 59320 199436
rect 258172 199384 258224 199436
rect 96620 198024 96672 198076
rect 259552 198024 259604 198076
rect 59084 197956 59136 198008
rect 273352 197956 273404 198008
rect 111800 196664 111852 196716
rect 262312 196664 262364 196716
rect 77392 196596 77444 196648
rect 264980 196596 265032 196648
rect 53656 195372 53708 195424
rect 240784 195372 240836 195424
rect 69020 195304 69072 195356
rect 324504 195304 324556 195356
rect 53564 195236 53616 195288
rect 336832 195236 336884 195288
rect 75184 193808 75236 193860
rect 269212 193808 269264 193860
rect 89720 192516 89772 192568
rect 252836 192516 252888 192568
rect 84200 192448 84252 192500
rect 337016 192448 337068 192500
rect 224224 191224 224276 191276
rect 256700 191224 256752 191276
rect 122104 191156 122156 191208
rect 250076 191156 250128 191208
rect 75920 191088 75972 191140
rect 582748 191088 582800 191140
rect 43444 189728 43496 189780
rect 109040 189728 109092 189780
rect 157984 189728 158036 189780
rect 339776 189728 339828 189780
rect 106188 189048 106240 189100
rect 211896 189048 211948 189100
rect 207664 188436 207716 188488
rect 269304 188436 269356 188488
rect 192484 188368 192536 188420
rect 267924 188368 267976 188420
rect 88432 188300 88484 188352
rect 328644 188300 328696 188352
rect 100668 187756 100720 187808
rect 171784 187756 171836 187808
rect 107568 187688 107620 187740
rect 207756 187688 207808 187740
rect 198004 187008 198056 187060
rect 256792 187008 256844 187060
rect 50988 186940 51040 186992
rect 338212 186940 338264 186992
rect 126796 186396 126848 186448
rect 171968 186396 172020 186448
rect 117228 186328 117280 186380
rect 214656 186328 214708 186380
rect 185584 185716 185636 185768
rect 255504 185716 255556 185768
rect 95240 185648 95292 185700
rect 321836 185648 321888 185700
rect 80060 185580 80112 185632
rect 322940 185580 322992 185632
rect 118608 184900 118660 184952
rect 170588 184900 170640 184952
rect 102140 184152 102192 184204
rect 321284 184152 321336 184204
rect 124128 183540 124180 183592
rect 167828 183540 167880 183592
rect 233884 183132 233936 183184
rect 260932 183132 260984 183184
rect 211804 183064 211856 183116
rect 261116 183064 261168 183116
rect 166264 182996 166316 183048
rect 332784 182996 332836 183048
rect 73160 182928 73212 182980
rect 321928 182928 321980 182980
rect 65984 182860 66036 182912
rect 338396 182860 338448 182912
rect 62028 182792 62080 182844
rect 345204 182792 345256 182844
rect 128176 182248 128228 182300
rect 166448 182248 166500 182300
rect 114376 182180 114428 182232
rect 169208 182180 169260 182232
rect 215944 181636 215996 181688
rect 259644 181636 259696 181688
rect 202144 181568 202196 181620
rect 259460 181568 259512 181620
rect 174544 181500 174596 181552
rect 265072 181500 265124 181552
rect 291844 181500 291896 181552
rect 332692 181500 332744 181552
rect 66168 181432 66220 181484
rect 251456 181432 251508 181484
rect 283564 181432 283616 181484
rect 343824 181432 343876 181484
rect 112168 180956 112220 181008
rect 167736 180956 167788 181008
rect 110696 180888 110748 180940
rect 169116 180888 169168 180940
rect 125048 180820 125100 180872
rect 211804 180820 211856 180872
rect 220084 180276 220136 180328
rect 258448 180276 258500 180328
rect 287704 180276 287756 180328
rect 335544 180276 335596 180328
rect 113364 180208 113416 180260
rect 336924 180208 336976 180260
rect 71780 180140 71832 180192
rect 339684 180140 339736 180192
rect 64696 180072 64748 180124
rect 342536 180072 342588 180124
rect 133144 179528 133196 179580
rect 165068 179528 165120 179580
rect 121184 179460 121236 179512
rect 166356 179460 166408 179512
rect 110052 179392 110104 179444
rect 214748 179392 214800 179444
rect 347044 179324 347096 179376
rect 579988 179324 580040 179376
rect 238024 179052 238076 179104
rect 258356 179052 258408 179104
rect 225604 178916 225656 178968
rect 258264 178916 258316 178968
rect 229744 178848 229796 178900
rect 258080 178848 258132 178900
rect 206284 178780 206336 178832
rect 249064 178780 249116 178832
rect 184204 178712 184256 178764
rect 242808 178712 242860 178764
rect 311164 178712 311216 178764
rect 335452 178712 335504 178764
rect 70400 178644 70452 178696
rect 328736 178644 328788 178696
rect 148232 178304 148284 178356
rect 169024 178304 169076 178356
rect 134708 178236 134760 178288
rect 165436 178236 165488 178288
rect 115848 178168 115900 178220
rect 166264 178168 166316 178220
rect 99104 178100 99156 178152
rect 170496 178100 170548 178152
rect 129464 178032 129516 178084
rect 208400 178032 208452 178084
rect 242808 177624 242860 177676
rect 261024 177624 261076 177676
rect 232504 177556 232556 177608
rect 259736 177556 259788 177608
rect 314016 177556 314068 177608
rect 334072 177556 334124 177608
rect 239404 177488 239456 177540
rect 267832 177488 267884 177540
rect 318064 177488 318116 177540
rect 338304 177488 338356 177540
rect 228364 177420 228416 177472
rect 266544 177420 266596 177472
rect 311256 177420 311308 177472
rect 331496 177420 331548 177472
rect 203524 177352 203576 177404
rect 249248 177352 249300 177404
rect 307024 177352 307076 177404
rect 341156 177352 341208 177404
rect 170404 177284 170456 177336
rect 321376 177284 321428 177336
rect 132040 176944 132092 176996
rect 165528 176944 165580 176996
rect 108120 176876 108172 176928
rect 170680 176876 170732 176928
rect 102048 176808 102100 176860
rect 171876 176808 171928 176860
rect 135720 176740 135772 176792
rect 213920 176740 213972 176792
rect 127072 176672 127124 176724
rect 211988 176672 212040 176724
rect 196624 176604 196676 176656
rect 248052 176604 248104 176656
rect 242164 176536 242216 176588
rect 249156 176604 249208 176656
rect 309876 176604 309928 176656
rect 321468 176604 321520 176656
rect 121920 176196 121972 176248
rect 167920 176196 167972 176248
rect 119436 176128 119488 176180
rect 166540 176128 166592 176180
rect 158904 176060 158956 176112
rect 214564 176060 214616 176112
rect 130752 175992 130804 176044
rect 214104 175992 214156 176044
rect 242256 175992 242308 176044
rect 255596 175992 255648 176044
rect 315304 175992 315356 176044
rect 332600 175992 332652 176044
rect 100760 175924 100812 175976
rect 210516 175924 210568 175976
rect 246304 175924 246356 175976
rect 262496 175924 262548 175976
rect 318248 175924 318300 175976
rect 335636 175924 335688 175976
rect 318156 175584 318208 175636
rect 321468 175584 321520 175636
rect 165436 175176 165488 175228
rect 213920 175176 213972 175228
rect 165068 175108 165120 175160
rect 214012 175108 214064 175160
rect 3240 164160 3292 164212
rect 39304 164160 39356 164212
rect 3424 150356 3476 150408
rect 25504 150356 25556 150408
rect 3240 137912 3292 137964
rect 14464 137912 14516 137964
rect 63408 122816 63460 122868
rect 66076 122816 66128 122868
rect 3424 111732 3476 111784
rect 13084 111732 13136 111784
rect 2780 97724 2832 97776
rect 4804 97724 4856 97776
rect 291844 174020 291896 174072
rect 307668 174020 307720 174072
rect 278228 173952 278280 174004
rect 306748 173952 306800 174004
rect 267004 173884 267056 173936
rect 307576 173884 307628 173936
rect 165528 173816 165580 173868
rect 213920 173816 213972 173868
rect 251824 172660 251876 172712
rect 259460 172660 259512 172712
rect 282184 172660 282236 172712
rect 307300 172660 307352 172712
rect 273996 172592 274048 172644
rect 307668 172592 307720 172644
rect 260288 172524 260340 172576
rect 306932 172524 306984 172576
rect 166448 172456 166500 172508
rect 214012 172456 214064 172508
rect 252008 172456 252060 172508
rect 258080 172456 258132 172508
rect 208400 172388 208452 172440
rect 213920 172388 213972 172440
rect 252468 172388 252520 172440
rect 261116 172388 261168 172440
rect 258080 172320 258132 172372
rect 258264 172320 258316 172372
rect 258264 172184 258316 172236
rect 258448 172184 258500 172236
rect 289268 171232 289320 171284
rect 307484 171232 307536 171284
rect 264336 171164 264388 171216
rect 307576 171164 307628 171216
rect 261760 171096 261812 171148
rect 307668 171096 307720 171148
rect 171968 171028 172020 171080
rect 213920 171028 213972 171080
rect 252100 171028 252152 171080
rect 262220 171028 262272 171080
rect 211988 170960 212040 171012
rect 214012 170960 214064 171012
rect 252468 170892 252520 170944
rect 256976 170892 257028 170944
rect 251824 169940 251876 169992
rect 258172 169940 258224 169992
rect 287888 169872 287940 169924
rect 306932 169872 306984 169924
rect 271328 169804 271380 169856
rect 307484 169804 307536 169856
rect 258816 169736 258868 169788
rect 307668 169736 307720 169788
rect 167828 169668 167880 169720
rect 213920 169668 213972 169720
rect 324320 169668 324372 169720
rect 332600 169668 332652 169720
rect 211804 169600 211856 169652
rect 214012 169600 214064 169652
rect 252008 169192 252060 169244
rect 258080 169192 258132 169244
rect 283564 168512 283616 168564
rect 307300 168512 307352 168564
rect 252468 168444 252520 168496
rect 259552 168444 259604 168496
rect 279608 168444 279660 168496
rect 307484 168444 307536 168496
rect 264244 168376 264296 168428
rect 307668 168376 307720 168428
rect 166356 168308 166408 168360
rect 214012 168308 214064 168360
rect 252100 168308 252152 168360
rect 260932 168308 260984 168360
rect 324412 168308 324464 168360
rect 338396 168308 338448 168360
rect 167920 168240 167972 168292
rect 213920 168240 213972 168292
rect 324320 168240 324372 168292
rect 334256 168240 334308 168292
rect 251916 168172 251968 168224
rect 255320 168172 255372 168224
rect 252468 168036 252520 168088
rect 259644 168036 259696 168088
rect 283656 167152 283708 167204
rect 307668 167152 307720 167204
rect 272524 167084 272576 167136
rect 307484 167084 307536 167136
rect 265900 167016 265952 167068
rect 307576 167016 307628 167068
rect 166540 166948 166592 167000
rect 213920 166948 213972 167000
rect 324320 166948 324372 167000
rect 345296 166948 345348 167000
rect 170588 166880 170640 166932
rect 214012 166880 214064 166932
rect 251824 166880 251876 166932
rect 260840 166880 260892 166932
rect 293224 165724 293276 165776
rect 307300 165724 307352 165776
rect 271144 165656 271196 165708
rect 307668 165656 307720 165708
rect 261668 165588 261720 165640
rect 307484 165588 307536 165640
rect 166264 165520 166316 165572
rect 213920 165520 213972 165572
rect 169208 165452 169260 165504
rect 214012 165452 214064 165504
rect 252468 165452 252520 165504
rect 261024 165452 261076 165504
rect 252376 165384 252428 165436
rect 266452 165384 266504 165436
rect 251364 164976 251416 165028
rect 252836 164976 252888 165028
rect 265808 164432 265860 164484
rect 307668 164432 307720 164484
rect 294788 164364 294840 164416
rect 307576 164364 307628 164416
rect 269856 164296 269908 164348
rect 307484 164296 307536 164348
rect 304356 164228 304408 164280
rect 306564 164228 306616 164280
rect 167736 164160 167788 164212
rect 213920 164160 213972 164212
rect 252468 164160 252520 164212
rect 267924 164160 267976 164212
rect 324412 164160 324464 164212
rect 345204 164160 345256 164212
rect 324320 164092 324372 164144
rect 335636 164092 335688 164144
rect 251364 163072 251416 163124
rect 254032 163072 254084 163124
rect 300124 163004 300176 163056
rect 307484 163004 307536 163056
rect 268384 162936 268436 162988
rect 307668 162936 307720 162988
rect 261576 162868 261628 162920
rect 307300 162868 307352 162920
rect 169116 162800 169168 162852
rect 213920 162800 213972 162852
rect 252468 162800 252520 162852
rect 269304 162800 269356 162852
rect 324320 162800 324372 162852
rect 336740 162800 336792 162852
rect 252100 162732 252152 162784
rect 264980 162732 265032 162784
rect 324412 162732 324464 162784
rect 331496 162732 331548 162784
rect 296076 161576 296128 161628
rect 307484 161576 307536 161628
rect 269764 161508 269816 161560
rect 307300 161508 307352 161560
rect 260196 161440 260248 161492
rect 307668 161440 307720 161492
rect 170680 161372 170732 161424
rect 213920 161372 213972 161424
rect 252468 161372 252520 161424
rect 266360 161372 266412 161424
rect 324688 161372 324740 161424
rect 339776 161372 339828 161424
rect 207756 161304 207808 161356
rect 214012 161304 214064 161356
rect 324320 161304 324372 161356
rect 335360 161304 335412 161356
rect 252008 160828 252060 160880
rect 255412 160828 255464 160880
rect 171876 160692 171928 160744
rect 213920 160692 213972 160744
rect 285036 160692 285088 160744
rect 307208 160692 307260 160744
rect 252100 160284 252152 160336
rect 258264 160284 258316 160336
rect 265716 160148 265768 160200
rect 307668 160148 307720 160200
rect 258724 160080 258776 160132
rect 306564 160080 306616 160132
rect 211896 160012 211948 160064
rect 214472 160012 214524 160064
rect 252468 160012 252520 160064
rect 262496 160012 262548 160064
rect 324320 160012 324372 160064
rect 328736 160012 328788 160064
rect 296260 158856 296312 158908
rect 307668 158856 307720 158908
rect 275284 158788 275336 158840
rect 307484 158788 307536 158840
rect 262956 158720 263008 158772
rect 306932 158720 306984 158772
rect 252376 158652 252428 158704
rect 276020 158652 276072 158704
rect 324412 158652 324464 158704
rect 338304 158652 338356 158704
rect 252468 158584 252520 158636
rect 265072 158584 265124 158636
rect 324320 158584 324372 158636
rect 332876 158584 332928 158636
rect 293592 157496 293644 157548
rect 307484 157496 307536 157548
rect 260104 157428 260156 157480
rect 306932 157428 306984 157480
rect 253204 157360 253256 157412
rect 307300 157360 307352 157412
rect 171784 157292 171836 157344
rect 213920 157292 213972 157344
rect 252376 157292 252428 157344
rect 267740 157292 267792 157344
rect 324320 157292 324372 157344
rect 346400 157292 346452 157344
rect 210516 157224 210568 157276
rect 214012 157224 214064 157276
rect 252468 157224 252520 157276
rect 263600 157224 263652 157276
rect 324412 157224 324464 157276
rect 343732 157224 343784 157276
rect 291936 156068 291988 156120
rect 306748 156068 306800 156120
rect 275376 156000 275428 156052
rect 307668 156000 307720 156052
rect 261484 155932 261536 155984
rect 307576 155932 307628 155984
rect 170496 155864 170548 155916
rect 213920 155864 213972 155916
rect 252376 155864 252428 155916
rect 278780 155864 278832 155916
rect 324320 155864 324372 155916
rect 347780 155864 347832 155916
rect 252468 155796 252520 155848
rect 270592 155796 270644 155848
rect 298836 154708 298888 154760
rect 307576 154708 307628 154760
rect 282368 154640 282420 154692
rect 307668 154640 307720 154692
rect 262864 154572 262916 154624
rect 307484 154572 307536 154624
rect 324320 154504 324372 154556
rect 328644 154504 328696 154556
rect 252376 154436 252428 154488
rect 269212 154436 269264 154488
rect 252468 154368 252520 154420
rect 271972 154368 272024 154420
rect 251180 154096 251232 154148
rect 253940 154096 253992 154148
rect 258908 153824 258960 153876
rect 307392 153824 307444 153876
rect 301596 153280 301648 153332
rect 307668 153280 307720 153332
rect 178684 153212 178736 153264
rect 213920 153212 213972 153264
rect 254676 153212 254728 153264
rect 307484 153212 307536 153264
rect 252468 153144 252520 153196
rect 273260 153144 273312 153196
rect 324320 153144 324372 153196
rect 347872 153144 347924 153196
rect 202144 151920 202196 151972
rect 213920 151920 213972 151972
rect 301504 151920 301556 151972
rect 307668 151920 307720 151972
rect 206284 151852 206336 151904
rect 214012 151852 214064 151904
rect 257344 151852 257396 151904
rect 307484 151852 307536 151904
rect 254768 151784 254820 151836
rect 307668 151784 307720 151836
rect 252468 151716 252520 151768
rect 262312 151716 262364 151768
rect 324320 151716 324372 151768
rect 327356 151716 327408 151768
rect 251272 151444 251324 151496
rect 254216 151444 254268 151496
rect 167644 151036 167696 151088
rect 184848 151036 184900 151088
rect 289176 150560 289228 150612
rect 307484 150560 307536 150612
rect 264428 150492 264480 150544
rect 307668 150492 307720 150544
rect 178868 150424 178920 150476
rect 214012 150424 214064 150476
rect 256148 150424 256200 150476
rect 306932 150424 306984 150476
rect 169024 150356 169076 150408
rect 213920 150356 213972 150408
rect 252284 150356 252336 150408
rect 278872 150356 278924 150408
rect 324320 150356 324372 150408
rect 346584 150356 346636 150408
rect 184848 150288 184900 150340
rect 214012 150288 214064 150340
rect 324412 150288 324464 150340
rect 346492 150288 346544 150340
rect 256056 149676 256108 149728
rect 307024 149676 307076 149728
rect 251732 149268 251784 149320
rect 256792 149268 256844 149320
rect 297640 149132 297692 149184
rect 307668 149132 307720 149184
rect 282460 149064 282512 149116
rect 306932 149064 306984 149116
rect 252468 148996 252520 149048
rect 271880 148996 271932 149048
rect 324320 148996 324372 149048
rect 345112 148996 345164 149048
rect 324412 148928 324464 148980
rect 337016 148928 337068 148980
rect 251272 148860 251324 148912
rect 254124 148860 254176 148912
rect 251916 148724 251968 148776
rect 255504 148724 255556 148776
rect 303068 147772 303120 147824
rect 307576 147772 307628 147824
rect 280896 147704 280948 147756
rect 307668 147704 307720 147756
rect 170404 147636 170456 147688
rect 213920 147636 213972 147688
rect 257528 147636 257580 147688
rect 306932 147636 306984 147688
rect 252468 147568 252520 147620
rect 281540 147568 281592 147620
rect 324320 147568 324372 147620
rect 340880 147568 340932 147620
rect 251732 147500 251784 147552
rect 274732 147500 274784 147552
rect 287980 146888 288032 146940
rect 307116 146888 307168 146940
rect 251732 146820 251784 146872
rect 255596 146820 255648 146872
rect 181444 146344 181496 146396
rect 213920 146344 213972 146396
rect 274088 146344 274140 146396
rect 307668 146344 307720 146396
rect 170496 146276 170548 146328
rect 214012 146276 214064 146328
rect 256240 146276 256292 146328
rect 306748 146276 306800 146328
rect 251916 146208 251968 146260
rect 273352 146208 273404 146260
rect 324412 146208 324464 146260
rect 338212 146208 338264 146260
rect 251732 146140 251784 146192
rect 266544 146140 266596 146192
rect 324320 146140 324372 146192
rect 334164 146140 334216 146192
rect 252100 146072 252152 146124
rect 263692 146072 263744 146124
rect 300492 146072 300544 146124
rect 306656 146072 306708 146124
rect 176016 144984 176068 145036
rect 214012 144984 214064 145036
rect 267096 144984 267148 145036
rect 307668 144984 307720 145036
rect 173164 144916 173216 144968
rect 213920 144916 213972 144968
rect 253480 144916 253532 144968
rect 307576 144916 307628 144968
rect 252376 144848 252428 144900
rect 270500 144848 270552 144900
rect 324320 144848 324372 144900
rect 342536 144848 342588 144900
rect 252468 144780 252520 144832
rect 267832 144780 267884 144832
rect 324412 144780 324464 144832
rect 331220 144780 331272 144832
rect 252100 144168 252152 144220
rect 264244 144168 264296 144220
rect 279700 144168 279752 144220
rect 307392 144168 307444 144220
rect 252468 144032 252520 144084
rect 259736 144032 259788 144084
rect 210424 143624 210476 143676
rect 214012 143624 214064 143676
rect 174544 143556 174596 143608
rect 213920 143556 213972 143608
rect 286416 143556 286468 143608
rect 307668 143556 307720 143608
rect 252468 143488 252520 143540
rect 269120 143488 269172 143540
rect 251916 142808 251968 142860
rect 293224 142808 293276 142860
rect 324320 142672 324372 142724
rect 327080 142672 327132 142724
rect 171784 142196 171836 142248
rect 213920 142196 213972 142248
rect 286324 142196 286376 142248
rect 307668 142196 307720 142248
rect 169024 142128 169076 142180
rect 214012 142128 214064 142180
rect 257436 142128 257488 142180
rect 306748 142128 306800 142180
rect 252468 142060 252520 142112
rect 258356 142060 258408 142112
rect 324320 142060 324372 142112
rect 349160 142060 349212 142112
rect 324504 141992 324556 142044
rect 333980 141992 334032 142044
rect 323676 141652 323728 141704
rect 324412 141652 324464 141704
rect 251824 141380 251876 141432
rect 275284 141380 275336 141432
rect 276756 141380 276808 141432
rect 307208 141380 307260 141432
rect 305920 140836 305972 140888
rect 307484 140836 307536 140888
rect 193864 140768 193916 140820
rect 213920 140768 213972 140820
rect 254584 140768 254636 140820
rect 307668 140768 307720 140820
rect 253388 140020 253440 140072
rect 306564 140020 306616 140072
rect 251364 139884 251416 139936
rect 256700 139884 256752 139936
rect 304448 139544 304500 139596
rect 307392 139544 307444 139596
rect 289084 139476 289136 139528
rect 307576 139476 307628 139528
rect 166264 139408 166316 139460
rect 213920 139408 213972 139460
rect 280804 139408 280856 139460
rect 307668 139408 307720 139460
rect 252468 139340 252520 139392
rect 280160 139340 280212 139392
rect 324320 139340 324372 139392
rect 350540 139340 350592 139392
rect 324504 139272 324556 139324
rect 332784 139272 332836 139324
rect 324964 139204 325016 139256
rect 327172 139204 327224 139256
rect 251548 138660 251600 138712
rect 278228 138660 278280 138712
rect 298744 138116 298796 138168
rect 307668 138116 307720 138168
rect 278136 138048 278188 138100
rect 307576 138048 307628 138100
rect 171876 137980 171928 138032
rect 213920 137980 213972 138032
rect 273904 137980 273956 138032
rect 307484 137980 307536 138032
rect 252468 137912 252520 137964
rect 277400 137912 277452 137964
rect 324320 137912 324372 137964
rect 342444 137912 342496 137964
rect 251364 137844 251416 137896
rect 274640 137844 274692 137896
rect 324504 137844 324556 137896
rect 330024 137844 330076 137896
rect 174820 137232 174872 137284
rect 214564 137232 214616 137284
rect 253296 137232 253348 137284
rect 307300 137232 307352 137284
rect 282276 136688 282328 136740
rect 307484 136688 307536 136740
rect 203524 136620 203576 136672
rect 213920 136620 213972 136672
rect 264244 136620 264296 136672
rect 306932 136620 306984 136672
rect 252468 136552 252520 136604
rect 291844 136552 291896 136604
rect 324504 136552 324556 136604
rect 343640 136552 343692 136604
rect 252376 136484 252428 136536
rect 267004 136484 267056 136536
rect 324320 136484 324372 136536
rect 339684 136484 339736 136536
rect 302884 135464 302936 135516
rect 307576 135464 307628 135516
rect 297364 135396 297416 135448
rect 307668 135396 307720 135448
rect 207756 135328 207808 135380
rect 214012 135328 214064 135380
rect 284944 135328 284996 135380
rect 307392 135328 307444 135380
rect 174636 135260 174688 135312
rect 213920 135260 213972 135312
rect 271236 135260 271288 135312
rect 307484 135260 307536 135312
rect 251640 135192 251692 135244
rect 273996 135192 274048 135244
rect 252468 134580 252520 134632
rect 260288 134580 260340 134632
rect 251548 134512 251600 134564
rect 283656 134512 283708 134564
rect 290648 134036 290700 134088
rect 307668 134036 307720 134088
rect 192484 133968 192536 134020
rect 213920 133968 213972 134020
rect 283748 133968 283800 134020
rect 307576 133968 307628 134020
rect 169116 133900 169168 133952
rect 214012 133900 214064 133952
rect 275284 133900 275336 133952
rect 306748 133900 306800 133952
rect 251456 133832 251508 133884
rect 289268 133832 289320 133884
rect 324320 133832 324372 133884
rect 328552 133832 328604 133884
rect 252468 133764 252520 133816
rect 264336 133764 264388 133816
rect 176108 133152 176160 133204
rect 214104 133152 214156 133204
rect 211896 132880 211948 132932
rect 213920 132880 213972 132932
rect 293224 132540 293276 132592
rect 307668 132540 307720 132592
rect 287704 132472 287756 132524
rect 307484 132472 307536 132524
rect 252284 132404 252336 132456
rect 287888 132404 287940 132456
rect 324504 132404 324556 132456
rect 345020 132404 345072 132456
rect 252008 132336 252060 132388
rect 271328 132336 271380 132388
rect 324320 132336 324372 132388
rect 341156 132336 341208 132388
rect 251364 132268 251416 132320
rect 261760 132268 261812 132320
rect 291844 131248 291896 131300
rect 306748 131248 306800 131300
rect 287796 131180 287848 131232
rect 307668 131180 307720 131232
rect 180156 131112 180208 131164
rect 213920 131112 213972 131164
rect 279516 131112 279568 131164
rect 307484 131112 307536 131164
rect 251732 131044 251784 131096
rect 285036 131044 285088 131096
rect 324320 131044 324372 131096
rect 331312 131044 331364 131096
rect 252008 130976 252060 131028
rect 279608 130976 279660 131028
rect 324412 130976 324464 131028
rect 331404 130976 331456 131028
rect 252468 129888 252520 129940
rect 258816 129888 258868 129940
rect 290556 129888 290608 129940
rect 306748 129888 306800 129940
rect 279424 129820 279476 129872
rect 306932 129820 306984 129872
rect 189724 129752 189776 129804
rect 213920 129752 213972 129804
rect 276664 129752 276716 129804
rect 307668 129752 307720 129804
rect 251732 129684 251784 129736
rect 283564 129684 283616 129736
rect 324320 129684 324372 129736
rect 330116 129684 330168 129736
rect 252100 129616 252152 129668
rect 272524 129616 272576 129668
rect 294604 128460 294656 128512
rect 307668 128460 307720 128512
rect 198004 128392 198056 128444
rect 214012 128392 214064 128444
rect 273996 128392 274048 128444
rect 307576 128392 307628 128444
rect 173256 128324 173308 128376
rect 213920 128324 213972 128376
rect 265624 128324 265676 128376
rect 307484 128324 307536 128376
rect 252008 128256 252060 128308
rect 271144 128256 271196 128308
rect 324320 128256 324372 128308
rect 329932 128256 329984 128308
rect 252468 128188 252520 128240
rect 265900 128188 265952 128240
rect 295984 127100 296036 127152
rect 307668 127100 307720 127152
rect 178776 127032 178828 127084
rect 213920 127032 213972 127084
rect 285036 127032 285088 127084
rect 307576 127032 307628 127084
rect 177304 126964 177356 127016
rect 214012 126964 214064 127016
rect 272524 126964 272576 127016
rect 307484 126964 307536 127016
rect 252100 126896 252152 126948
rect 269856 126896 269908 126948
rect 324320 126896 324372 126948
rect 328460 126896 328512 126948
rect 392584 126896 392636 126948
rect 580172 126896 580224 126948
rect 252468 126828 252520 126880
rect 261668 126828 261720 126880
rect 251272 126216 251324 126268
rect 294788 126216 294840 126268
rect 294696 125740 294748 125792
rect 307668 125740 307720 125792
rect 169208 125672 169260 125724
rect 214012 125672 214064 125724
rect 289360 125672 289412 125724
rect 306748 125672 306800 125724
rect 166356 125604 166408 125656
rect 213920 125604 213972 125656
rect 271144 125604 271196 125656
rect 307484 125604 307536 125656
rect 252468 125536 252520 125588
rect 304356 125536 304408 125588
rect 252376 125468 252428 125520
rect 265808 125468 265860 125520
rect 252284 124856 252336 124908
rect 300124 124856 300176 124908
rect 300308 124312 300360 124364
rect 306748 124312 306800 124364
rect 173348 124244 173400 124296
rect 213920 124244 213972 124296
rect 304264 124244 304316 124296
rect 307484 124244 307536 124296
rect 170588 124176 170640 124228
rect 214012 124176 214064 124228
rect 290464 124176 290516 124228
rect 307668 124176 307720 124228
rect 252468 124108 252520 124160
rect 268384 124108 268436 124160
rect 324320 124108 324372 124160
rect 342352 124108 342404 124160
rect 252008 124040 252060 124092
rect 261576 124040 261628 124092
rect 323584 124040 323636 124092
rect 324504 124040 324556 124092
rect 252100 123428 252152 123480
rect 301596 123428 301648 123480
rect 211804 123360 211856 123412
rect 214012 123360 214064 123412
rect 300216 122952 300268 123004
rect 307668 122952 307720 123004
rect 302976 122884 303028 122936
rect 307576 122884 307628 122936
rect 174728 122816 174780 122868
rect 213920 122816 213972 122868
rect 283564 122816 283616 122868
rect 306564 122816 306616 122868
rect 252468 122748 252520 122800
rect 296076 122748 296128 122800
rect 324688 122748 324740 122800
rect 343824 122748 343876 122800
rect 252376 122680 252428 122732
rect 269764 122680 269816 122732
rect 324320 122680 324372 122732
rect 338120 122680 338172 122732
rect 252468 122000 252520 122052
rect 260196 122000 260248 122052
rect 297548 121592 297600 121644
rect 307668 121592 307720 121644
rect 207664 121524 207716 121576
rect 214012 121524 214064 121576
rect 293316 121524 293368 121576
rect 307576 121524 307628 121576
rect 180248 121456 180300 121508
rect 213920 121456 213972 121508
rect 268384 121456 268436 121508
rect 307484 121456 307536 121508
rect 251916 121388 251968 121440
rect 287980 121388 288032 121440
rect 324412 121388 324464 121440
rect 339500 121388 339552 121440
rect 252468 121320 252520 121372
rect 265716 121320 265768 121372
rect 324320 121320 324372 121372
rect 335544 121320 335596 121372
rect 252376 121252 252428 121304
rect 258724 121252 258776 121304
rect 301688 120232 301740 120284
rect 307668 120232 307720 120284
rect 185584 120164 185636 120216
rect 214012 120164 214064 120216
rect 287888 120164 287940 120216
rect 307484 120164 307536 120216
rect 167644 120096 167696 120148
rect 213920 120096 213972 120148
rect 267004 120096 267056 120148
rect 307576 120096 307628 120148
rect 252468 120028 252520 120080
rect 296260 120028 296312 120080
rect 251364 119960 251416 120012
rect 262956 119960 263008 120012
rect 263048 119348 263100 119400
rect 307208 119348 307260 119400
rect 210516 118804 210568 118856
rect 214104 118804 214156 118856
rect 296168 118804 296220 118856
rect 306748 118804 306800 118856
rect 196624 118736 196676 118788
rect 214012 118736 214064 118788
rect 251180 118736 251232 118788
rect 253204 118736 253256 118788
rect 299020 118736 299072 118788
rect 307668 118736 307720 118788
rect 166448 118668 166500 118720
rect 213920 118668 213972 118720
rect 251824 118600 251876 118652
rect 293592 118600 293644 118652
rect 324412 118600 324464 118652
rect 341064 118600 341116 118652
rect 252468 118532 252520 118584
rect 260104 118532 260156 118584
rect 324320 118532 324372 118584
rect 339592 118532 339644 118584
rect 167736 117920 167788 117972
rect 213276 117920 213328 117972
rect 251640 117920 251692 117972
rect 298836 117920 298888 117972
rect 300400 117444 300452 117496
rect 307576 117444 307628 117496
rect 296076 117376 296128 117428
rect 307668 117376 307720 117428
rect 210608 117308 210660 117360
rect 213920 117308 213972 117360
rect 293408 117308 293460 117360
rect 307484 117308 307536 117360
rect 251916 117240 251968 117292
rect 291936 117240 291988 117292
rect 324412 117240 324464 117292
rect 336924 117240 336976 117292
rect 252376 117172 252428 117224
rect 261484 117172 261536 117224
rect 324320 117172 324372 117224
rect 332692 117172 332744 117224
rect 252468 117104 252520 117156
rect 258908 117104 258960 117156
rect 189816 116016 189868 116068
rect 213920 116016 213972 116068
rect 292028 116016 292080 116068
rect 307668 116016 307720 116068
rect 169300 115948 169352 116000
rect 214012 115948 214064 116000
rect 265716 115948 265768 116000
rect 306748 115948 306800 116000
rect 252468 115880 252520 115932
rect 275376 115880 275428 115932
rect 324320 115880 324372 115932
rect 336832 115880 336884 115932
rect 252376 115812 252428 115864
rect 262864 115812 262916 115864
rect 168196 115200 168248 115252
rect 178868 115200 178920 115252
rect 211988 114588 212040 114640
rect 214012 114588 214064 114640
rect 282184 114588 282236 114640
rect 307668 114588 307720 114640
rect 178960 114520 179012 114572
rect 213920 114520 213972 114572
rect 264336 114520 264388 114572
rect 306748 114520 306800 114572
rect 252468 114452 252520 114504
rect 282368 114452 282420 114504
rect 324320 114452 324372 114504
rect 340972 114452 341024 114504
rect 252376 114384 252428 114436
rect 276756 114384 276808 114436
rect 324412 114384 324464 114436
rect 334072 114384 334124 114436
rect 252100 113704 252152 113756
rect 254676 113704 254728 113756
rect 298836 113296 298888 113348
rect 306748 113296 306800 113348
rect 184204 113228 184256 113280
rect 214012 113228 214064 113280
rect 291936 113228 291988 113280
rect 307576 113228 307628 113280
rect 171968 113160 172020 113212
rect 213920 113160 213972 113212
rect 279608 113160 279660 113212
rect 307668 113160 307720 113212
rect 252468 113092 252520 113144
rect 300492 113092 300544 113144
rect 324320 113092 324372 113144
rect 335452 113092 335504 113144
rect 252376 112412 252428 112464
rect 264428 112412 264480 112464
rect 269396 112412 269448 112464
rect 307024 112412 307076 112464
rect 177396 111868 177448 111920
rect 214012 111868 214064 111920
rect 300124 111868 300176 111920
rect 307576 111868 307628 111920
rect 170680 111800 170732 111852
rect 213920 111800 213972 111852
rect 251548 111800 251600 111852
rect 254768 111800 254820 111852
rect 297456 111800 297508 111852
rect 307668 111800 307720 111852
rect 167920 111732 167972 111784
rect 174820 111732 174872 111784
rect 252468 111732 252520 111784
rect 301504 111732 301556 111784
rect 324320 111732 324372 111784
rect 342260 111732 342312 111784
rect 252284 111664 252336 111716
rect 257344 111664 257396 111716
rect 251732 111052 251784 111104
rect 297640 111052 297692 111104
rect 301780 110576 301832 110628
rect 307576 110576 307628 110628
rect 202236 110508 202288 110560
rect 213920 110508 213972 110560
rect 303160 110508 303212 110560
rect 307668 110508 307720 110560
rect 199384 110440 199436 110492
rect 214012 110440 214064 110492
rect 296260 110440 296312 110492
rect 307484 110440 307536 110492
rect 252468 110372 252520 110424
rect 289176 110372 289228 110424
rect 251272 110304 251324 110356
rect 257528 110304 257580 110356
rect 251916 109284 251968 109336
rect 256148 109284 256200 109336
rect 304540 109148 304592 109200
rect 307484 109148 307536 109200
rect 278228 109080 278280 109132
rect 307576 109080 307628 109132
rect 206376 109012 206428 109064
rect 213920 109012 213972 109064
rect 261484 109012 261536 109064
rect 307668 109012 307720 109064
rect 251364 108944 251416 108996
rect 303068 108944 303120 108996
rect 252468 108876 252520 108928
rect 282460 108876 282512 108928
rect 324320 107992 324372 108044
rect 327264 107992 327316 108044
rect 251180 107856 251232 107908
rect 253480 107856 253532 107908
rect 282368 107856 282420 107908
rect 307668 107856 307720 107908
rect 203616 107720 203668 107772
rect 214012 107720 214064 107772
rect 301596 107720 301648 107772
rect 306748 107720 306800 107772
rect 174820 107652 174872 107704
rect 213920 107652 213972 107704
rect 304356 107652 304408 107704
rect 307576 107652 307628 107704
rect 251364 107584 251416 107636
rect 280896 107584 280948 107636
rect 252468 107516 252520 107568
rect 269396 107516 269448 107568
rect 301504 106428 301556 106480
rect 307484 106428 307536 106480
rect 283656 106360 283708 106412
rect 307576 106360 307628 106412
rect 167736 106292 167788 106344
rect 213920 106292 213972 106344
rect 269856 106292 269908 106344
rect 307668 106292 307720 106344
rect 252008 106224 252060 106276
rect 279700 106224 279752 106276
rect 252284 106156 252336 106208
rect 256240 106156 256292 106208
rect 252008 105544 252060 105596
rect 305828 105544 305880 105596
rect 280896 105000 280948 105052
rect 307668 105000 307720 105052
rect 212080 104932 212132 104984
rect 214012 104932 214064 104984
rect 289176 104932 289228 104984
rect 306564 104932 306616 104984
rect 209044 104864 209096 104916
rect 213920 104864 213972 104916
rect 252468 104796 252520 104848
rect 305920 104796 305972 104848
rect 251548 104116 251600 104168
rect 286416 104116 286468 104168
rect 253204 103640 253256 103692
rect 307668 103640 307720 103692
rect 287980 103572 288032 103624
rect 307576 103572 307628 103624
rect 209136 103504 209188 103556
rect 213920 103504 213972 103556
rect 252468 103436 252520 103488
rect 267096 103436 267148 103488
rect 251180 102756 251232 102808
rect 253388 102756 253440 102808
rect 298928 102280 298980 102332
rect 307484 102280 307536 102332
rect 252100 102212 252152 102264
rect 257436 102212 257488 102264
rect 269764 102212 269816 102264
rect 306748 102212 306800 102264
rect 204904 102144 204956 102196
rect 213920 102144 213972 102196
rect 257344 102144 257396 102196
rect 306932 102144 306984 102196
rect 252468 102076 252520 102128
rect 293500 102076 293552 102128
rect 252376 102008 252428 102060
rect 286324 102008 286376 102060
rect 303068 100852 303120 100904
rect 307576 100852 307628 100904
rect 207848 100784 207900 100836
rect 214012 100784 214064 100836
rect 293592 100784 293644 100836
rect 307668 100784 307720 100836
rect 172060 100716 172112 100768
rect 213920 100716 213972 100768
rect 286416 100716 286468 100768
rect 307484 100716 307536 100768
rect 252100 100648 252152 100700
rect 304448 100648 304500 100700
rect 395344 100648 395396 100700
rect 580172 100648 580224 100700
rect 252468 100580 252520 100632
rect 292120 100580 292172 100632
rect 251180 100104 251232 100156
rect 253296 100104 253348 100156
rect 173440 99424 173492 99476
rect 213920 99424 213972 99476
rect 304632 99424 304684 99476
rect 307484 99424 307536 99476
rect 167920 99356 167972 99408
rect 214012 99356 214064 99408
rect 289268 99356 289320 99408
rect 307668 99356 307720 99408
rect 252192 99288 252244 99340
rect 269948 99288 270000 99340
rect 252284 99152 252336 99204
rect 256056 99152 256108 99204
rect 251180 98608 251232 98660
rect 254584 98608 254636 98660
rect 294788 98132 294840 98184
rect 307668 98132 307720 98184
rect 286324 98064 286376 98116
rect 307484 98064 307536 98116
rect 167828 97996 167880 98048
rect 213920 97996 213972 98048
rect 260104 97996 260156 98048
rect 307576 97996 307628 98048
rect 252468 97860 252520 97912
rect 263048 97860 263100 97912
rect 249524 97520 249576 97572
rect 255964 97520 256016 97572
rect 166540 97248 166592 97300
rect 214564 97248 214616 97300
rect 292120 96704 292172 96756
rect 306748 96704 306800 96756
rect 164884 96636 164936 96688
rect 213920 96636 213972 96688
rect 256056 96636 256108 96688
rect 307484 96636 307536 96688
rect 278044 96568 278096 96620
rect 321468 96568 321520 96620
rect 250444 95208 250496 95260
rect 307668 95208 307720 95260
rect 196716 95140 196768 95192
rect 324320 95140 324372 95192
rect 308588 95072 308640 95124
rect 321560 95072 321612 95124
rect 309784 95004 309836 95056
rect 324412 95004 324464 95056
rect 308404 94936 308456 94988
rect 321744 94936 321796 94988
rect 239404 94460 239456 94512
rect 248420 94460 248472 94512
rect 134340 94120 134392 94172
rect 170496 94120 170548 94172
rect 117964 94052 118016 94104
rect 171876 94052 171928 94104
rect 105452 93984 105504 94036
rect 178960 93984 179012 94036
rect 129372 93916 129424 93968
rect 210424 93916 210476 93968
rect 119528 93848 119580 93900
rect 207664 93848 207716 93900
rect 67364 93780 67416 93832
rect 209044 93780 209096 93832
rect 188344 93712 188396 93764
rect 324504 93712 324556 93764
rect 151728 93372 151780 93424
rect 178684 93372 178736 93424
rect 130752 93304 130804 93356
rect 173164 93304 173216 93356
rect 115848 93236 115900 93288
rect 167644 93236 167696 93288
rect 110696 93168 110748 93220
rect 169116 93168 169168 93220
rect 125508 93100 125560 93152
rect 214840 93100 214892 93152
rect 115480 92420 115532 92472
rect 203524 92420 203576 92472
rect 116768 92352 116820 92404
rect 176108 92352 176160 92404
rect 85672 92284 85724 92336
rect 125508 92284 125560 92336
rect 151544 92284 151596 92336
rect 206284 92284 206336 92336
rect 152096 92216 152148 92268
rect 202144 92216 202196 92268
rect 119712 92148 119764 92200
rect 166540 92148 166592 92200
rect 125784 92080 125836 92132
rect 171784 92080 171836 92132
rect 180064 91740 180116 91792
rect 307300 91740 307352 91792
rect 91652 91060 91704 91112
rect 108304 91060 108356 91112
rect 114192 90992 114244 91044
rect 207756 90992 207808 91044
rect 107752 90924 107804 90976
rect 189816 90924 189868 90976
rect 151452 90856 151504 90908
rect 215944 90856 215996 90908
rect 122472 90788 122524 90840
rect 166264 90788 166316 90840
rect 125508 90720 125560 90772
rect 166356 90720 166408 90772
rect 207664 90312 207716 90364
rect 307116 90312 307168 90364
rect 90548 89632 90600 89684
rect 212080 89632 212132 89684
rect 99748 89564 99800 89616
rect 199384 89564 199436 89616
rect 89352 89496 89404 89548
rect 167920 89496 167972 89548
rect 103152 89428 103204 89480
rect 171968 89428 172020 89480
rect 117136 89360 117188 89412
rect 185584 89360 185636 89412
rect 136456 89292 136508 89344
rect 170404 89292 170456 89344
rect 67272 88272 67324 88324
rect 214748 88272 214800 88324
rect 115296 88204 115348 88256
rect 196624 88204 196676 88256
rect 111984 88136 112036 88188
rect 174636 88136 174688 88188
rect 109224 88068 109276 88120
rect 169300 88068 169352 88120
rect 133144 88000 133196 88052
rect 181444 88000 181496 88052
rect 126520 87932 126572 87984
rect 169208 87932 169260 87984
rect 75368 86912 75420 86964
rect 214564 86912 214616 86964
rect 88064 86844 88116 86896
rect 173440 86844 173492 86896
rect 109776 86776 109828 86828
rect 192484 86776 192536 86828
rect 112352 86708 112404 86760
rect 166448 86708 166500 86760
rect 124128 86640 124180 86692
rect 170588 86640 170640 86692
rect 3148 85484 3200 85536
rect 44824 85484 44876 85536
rect 111616 85484 111668 85536
rect 210608 85484 210660 85536
rect 66076 85416 66128 85468
rect 164884 85416 164936 85468
rect 104348 85348 104400 85400
rect 184204 85348 184256 85400
rect 100576 85280 100628 85332
rect 170680 85280 170732 85332
rect 122840 85212 122892 85264
rect 173348 85212 173400 85264
rect 132040 85144 132092 85196
rect 176016 85144 176068 85196
rect 63408 84124 63460 84176
rect 216036 84124 216088 84176
rect 107476 84056 107528 84108
rect 211988 84056 212040 84108
rect 101864 83988 101916 84040
rect 198004 83988 198056 84040
rect 118608 83920 118660 83972
rect 180248 83920 180300 83972
rect 67456 82764 67508 82816
rect 204904 82764 204956 82816
rect 99104 82696 99156 82748
rect 202236 82696 202288 82748
rect 110328 82628 110380 82680
rect 213184 82628 213236 82680
rect 121368 82560 121420 82612
rect 174728 82560 174780 82612
rect 126888 82492 126940 82544
rect 169024 82492 169076 82544
rect 108304 81336 108356 81388
rect 214656 81336 214708 81388
rect 97816 81268 97868 81320
rect 178776 81268 178828 81320
rect 86868 81200 86920 81252
rect 167828 81200 167880 81252
rect 93768 81132 93820 81184
rect 167736 81132 167788 81184
rect 125416 81064 125468 81116
rect 193864 81064 193916 81116
rect 67548 79976 67600 80028
rect 207848 79976 207900 80028
rect 114468 79908 114520 79960
rect 210516 79908 210568 79960
rect 103428 79840 103480 79892
rect 189724 79840 189776 79892
rect 95056 79772 95108 79824
rect 174820 79772 174872 79824
rect 97908 78616 97960 78668
rect 206376 78616 206428 78668
rect 122748 78548 122800 78600
rect 211804 78548 211856 78600
rect 99288 78480 99340 78532
rect 177304 78480 177356 78532
rect 99196 78412 99248 78464
rect 173256 78412 173308 78464
rect 85488 77188 85540 77240
rect 172060 77188 172112 77240
rect 77300 76576 77352 76628
rect 290648 76576 290700 76628
rect 89720 76508 89772 76560
rect 306012 76508 306064 76560
rect 95148 75828 95200 75880
rect 203616 75828 203668 75880
rect 102048 75760 102100 75812
rect 177396 75760 177448 75812
rect 107660 75148 107712 75200
rect 303160 75148 303212 75200
rect 103520 73856 103572 73908
rect 304540 73856 304592 73908
rect 9680 73788 9732 73840
rect 294696 73788 294748 73840
rect 122840 72496 122892 72548
rect 289360 72496 289412 72548
rect 53840 72428 53892 72480
rect 305828 72428 305880 72480
rect 62120 71068 62172 71120
rect 293408 71068 293460 71120
rect 68284 71000 68336 71052
rect 307208 71000 307260 71052
rect 66260 69640 66312 69692
rect 299020 69640 299072 69692
rect 57980 68348 58032 68400
rect 287980 68348 288032 68400
rect 20720 68280 20772 68332
rect 304632 68280 304684 68332
rect 71780 66920 71832 66972
rect 269856 66920 269908 66972
rect 26240 66852 26292 66904
rect 293592 66852 293644 66904
rect 82820 65492 82872 65544
rect 282368 65492 282420 65544
rect 33140 64132 33192 64184
rect 286416 64132 286468 64184
rect 80060 62840 80112 62892
rect 267004 62840 267056 62892
rect 35900 62772 35952 62824
rect 303068 62772 303120 62824
rect 93860 61344 93912 61396
rect 268384 61344 268436 61396
rect 175924 60664 175976 60716
rect 580172 60664 580224 60716
rect 118700 59984 118752 60036
rect 300308 59984 300360 60036
rect 3056 59304 3108 59356
rect 48964 59304 49016 59356
rect 110420 58692 110472 58744
rect 301780 58692 301832 58744
rect 48320 58624 48372 58676
rect 292028 58624 292080 58676
rect 81440 57196 81492 57248
rect 283748 57196 283800 57248
rect 40040 55904 40092 55956
rect 257344 55904 257396 55956
rect 55220 55836 55272 55888
rect 300400 55836 300452 55888
rect 92480 54544 92532 54596
rect 271236 54544 271288 54596
rect 15200 54476 15252 54528
rect 292120 54476 292172 54528
rect 99380 53116 99432 53168
rect 284944 53116 284996 53168
rect 24860 53048 24912 53100
rect 294788 53048 294840 53100
rect 12440 51688 12492 51740
rect 279608 51688 279660 51740
rect 84200 50396 84252 50448
rect 287888 50396 287940 50448
rect 27620 50328 27672 50380
rect 272524 50328 272576 50380
rect 86960 49036 87012 49088
rect 297548 49036 297600 49088
rect 23480 48968 23532 49020
rect 285036 48968 285088 49020
rect 88340 47608 88392 47660
rect 302884 47608 302936 47660
rect 17960 47540 18012 47592
rect 291936 47540 291988 47592
rect 106280 46180 106332 46232
rect 282276 46180 282328 46232
rect 3424 45500 3476 45552
rect 43444 45500 43496 45552
rect 102140 44888 102192 44940
rect 302976 44888 303028 44940
rect 63500 44820 63552 44872
rect 279516 44820 279568 44872
rect 56600 43392 56652 43444
rect 291844 43392 291896 43444
rect 85580 42100 85632 42152
rect 275284 42100 275336 42152
rect 98000 42032 98052 42084
rect 300216 42032 300268 42084
rect 91100 40740 91152 40792
rect 293316 40740 293368 40792
rect 19340 40672 19392 40724
rect 295984 40672 296036 40724
rect 95240 39380 95292 39432
rect 297364 39380 297416 39432
rect 31760 39312 31812 39364
rect 294604 39312 294656 39364
rect 77392 37952 77444 38004
rect 301688 37952 301740 38004
rect 38660 37884 38712 37936
rect 265624 37884 265676 37936
rect 73160 36592 73212 36644
rect 296168 36592 296220 36644
rect 42800 36524 42852 36576
rect 276664 36524 276716 36576
rect 69020 35232 69072 35284
rect 305736 35232 305788 35284
rect 16580 35164 16632 35216
rect 289268 35164 289320 35216
rect 113180 33804 113232 33856
rect 298744 33804 298796 33856
rect 3240 33736 3292 33788
rect 46204 33736 46256 33788
rect 52460 33736 52512 33788
rect 296076 33736 296128 33788
rect 27712 32376 27764 32428
rect 298836 32376 298888 32428
rect 85672 31084 85724 31136
rect 304356 31084 304408 31136
rect 44180 31016 44232 31068
rect 298928 31016 298980 31068
rect 118792 29656 118844 29708
rect 297456 29656 297508 29708
rect 37280 29588 37332 29640
rect 264336 29588 264388 29640
rect 114560 28296 114612 28348
rect 296260 28296 296312 28348
rect 44272 28228 44324 28280
rect 265716 28228 265768 28280
rect 121460 26936 121512 26988
rect 300124 26936 300176 26988
rect 52552 26868 52604 26920
rect 290556 26868 290608 26920
rect 100760 25576 100812 25628
rect 278228 25576 278280 25628
rect 60740 25508 60792 25560
rect 287796 25508 287848 25560
rect 93952 24148 94004 24200
rect 301596 24148 301648 24200
rect 13820 24080 13872 24132
rect 271144 24080 271196 24132
rect 75920 22720 75972 22772
rect 283656 22720 283708 22772
rect 78680 21428 78732 21480
rect 301504 21428 301556 21480
rect 35992 21360 36044 21412
rect 273996 21360 274048 21412
rect 3516 20612 3568 20664
rect 32404 20612 32456 20664
rect 3424 19932 3476 19984
rect 57244 19932 57296 19984
rect 115940 19932 115992 19984
rect 304264 19932 304316 19984
rect 69112 18640 69164 18692
rect 289176 18640 289228 18692
rect 45560 18572 45612 18624
rect 279424 18572 279476 18624
rect 64880 17280 64932 17332
rect 305644 17280 305696 17332
rect 11152 17212 11204 17264
rect 256056 17212 256108 17264
rect 61568 15920 61620 15972
rect 280896 15920 280948 15972
rect 20168 15852 20220 15904
rect 260104 15852 260156 15904
rect 105728 14424 105780 14476
rect 283564 14424 283616 14476
rect 124680 13132 124732 13184
rect 280804 13132 280856 13184
rect 47400 13064 47452 13116
rect 269764 13064 269816 13116
rect 117320 11772 117372 11824
rect 278136 11772 278188 11824
rect 7656 11704 7708 11756
rect 286324 11704 286376 11756
rect 110512 10344 110564 10396
rect 264244 10344 264296 10396
rect 2872 10276 2924 10328
rect 289084 10276 289136 10328
rect 7472 9596 7524 9648
rect 8208 9596 8260 9648
rect 251180 9596 251232 9648
rect 75000 8916 75052 8968
rect 293224 8916 293276 8968
rect 1676 8304 1728 8356
rect 7472 8304 7524 8356
rect 63500 8236 63552 8288
rect 64788 8236 64840 8288
rect 248420 8236 248472 8288
rect 572 7556 624 7608
rect 63500 7556 63552 7608
rect 71504 7556 71556 7608
rect 287704 7556 287756 7608
rect 31300 6128 31352 6180
rect 282184 6128 282236 6180
rect 97448 4836 97500 4888
rect 261484 4836 261536 4888
rect 6460 4768 6512 4820
rect 307024 4768 307076 4820
rect 235816 3952 235868 4004
rect 239404 3952 239456 4004
rect 41880 3544 41932 3596
rect 68284 3544 68336 3596
rect 2780 3476 2832 3528
rect 3700 3476 3752 3528
rect 11060 3476 11112 3528
rect 11980 3476 12032 3528
rect 27620 3476 27672 3528
rect 28540 3476 28592 3528
rect 35900 3476 35952 3528
rect 36820 3476 36872 3528
rect 67916 3476 67968 3528
rect 69020 3476 69072 3528
rect 69940 3476 69992 3528
rect 77300 3544 77352 3596
rect 78220 3544 78272 3596
rect 93860 3544 93912 3596
rect 94780 3544 94832 3596
rect 103336 3544 103388 3596
rect 112444 3544 112496 3596
rect 112812 3612 112864 3664
rect 180064 3612 180116 3664
rect 207664 3544 207716 3596
rect 110420 3476 110472 3528
rect 111616 3476 111668 3528
rect 118700 3476 118752 3528
rect 119896 3476 119948 3528
rect 121092 3476 121144 3528
rect 273904 3476 273956 3528
rect 51356 3408 51408 3460
rect 253204 3408 253256 3460
rect 109316 2116 109368 2168
rect 290464 2116 290516 2168
rect 5264 2048 5316 2100
rect 250444 2048 250496 2100
<< obsm1 >>
rect 68800 95100 164756 174600
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 700330 8156 703520
rect 24320 700330 24348 703520
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 8944 700324 8996 700330
rect 8944 700266 8996 700272
rect 24308 700324 24360 700330
rect 24308 700266 24360 700272
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 2778 606112 2834 606121
rect 2778 606047 2834 606056
rect 2792 605946 2820 606047
rect 2780 605940 2832 605946
rect 2780 605882 2832 605888
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3238 566944 3294 566953
rect 3238 566879 3294 566888
rect 3252 565894 3280 566879
rect 3240 565888 3292 565894
rect 3240 565830 3292 565836
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553450 3372 553823
rect 3332 553444 3384 553450
rect 3332 553386 3384 553392
rect 2962 527912 3018 527921
rect 2962 527847 3018 527856
rect 2976 527202 3004 527847
rect 2964 527196 3016 527202
rect 2964 527138 3016 527144
rect 3330 501800 3386 501809
rect 3330 501735 3386 501744
rect 3344 501022 3372 501735
rect 3332 501016 3384 501022
rect 3332 500958 3384 500964
rect 3054 475688 3110 475697
rect 3054 475623 3110 475632
rect 3068 474774 3096 475623
rect 3056 474768 3108 474774
rect 3056 474710 3108 474716
rect 3330 462632 3386 462641
rect 3330 462567 3386 462576
rect 3344 462398 3372 462567
rect 3332 462392 3384 462398
rect 3332 462334 3384 462340
rect 3330 449576 3386 449585
rect 3330 449511 3386 449520
rect 3344 448594 3372 449511
rect 3332 448588 3384 448594
rect 3332 448530 3384 448536
rect 3330 423600 3386 423609
rect 3330 423535 3386 423544
rect 3344 423366 3372 423535
rect 3332 423360 3384 423366
rect 3332 423302 3384 423308
rect 3330 410544 3386 410553
rect 3330 410479 3386 410488
rect 3344 409902 3372 410479
rect 3332 409896 3384 409902
rect 3332 409838 3384 409844
rect 3332 397520 3384 397526
rect 3330 397488 3332 397497
rect 3384 397488 3386 397497
rect 3330 397423 3386 397432
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 3344 371278 3372 371311
rect 3332 371272 3384 371278
rect 3332 371214 3384 371220
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3344 357474 3372 358391
rect 3332 357468 3384 357474
rect 3332 357410 3384 357416
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 3436 326398 3464 684247
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3514 658200 3570 658209
rect 3514 658135 3570 658144
rect 3528 656946 3556 658135
rect 3516 656940 3568 656946
rect 3516 656882 3568 656888
rect 3516 632120 3568 632126
rect 3514 632088 3516 632097
rect 3568 632088 3570 632097
rect 3514 632023 3570 632032
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3528 618322 3556 619103
rect 3516 618316 3568 618322
rect 3516 618258 3568 618264
rect 4804 605940 4856 605946
rect 4804 605882 4856 605888
rect 3514 514856 3570 514865
rect 3514 514791 3570 514800
rect 3424 326392 3476 326398
rect 3424 326334 3476 326340
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3344 318850 3372 319223
rect 3332 318844 3384 318850
rect 3332 318786 3384 318792
rect 3528 313954 3556 514791
rect 3516 313948 3568 313954
rect 3516 313890 3568 313896
rect 4816 312594 4844 605882
rect 7564 423360 7616 423366
rect 7564 423302 7616 423308
rect 4804 312588 4856 312594
rect 4804 312530 4856 312536
rect 3422 306232 3478 306241
rect 3422 306167 3478 306176
rect 3436 305114 3464 306167
rect 3424 305108 3476 305114
rect 3424 305050 3476 305056
rect 7576 298790 7604 423302
rect 7564 298784 7616 298790
rect 7564 298726 7616 298732
rect 2778 293176 2834 293185
rect 2778 293111 2834 293120
rect 2792 292874 2820 293111
rect 2780 292868 2832 292874
rect 2780 292810 2832 292816
rect 4804 292868 4856 292874
rect 4804 292810 4856 292816
rect 3424 291848 3476 291854
rect 3424 291790 3476 291796
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3160 253978 3188 254079
rect 3148 253972 3200 253978
rect 3148 253914 3200 253920
rect 3054 241088 3110 241097
rect 3054 241023 3110 241032
rect 3068 240174 3096 241023
rect 3056 240168 3108 240174
rect 3056 240110 3108 240116
rect 3056 202836 3108 202842
rect 3056 202778 3108 202784
rect 3068 201929 3096 202778
rect 3054 201920 3110 201929
rect 3054 201855 3110 201864
rect 3436 188873 3464 291790
rect 3514 267200 3570 267209
rect 3514 267135 3570 267144
rect 3528 238746 3556 267135
rect 4816 244254 4844 292810
rect 8208 292596 8260 292602
rect 8208 292538 8260 292544
rect 4804 244248 4856 244254
rect 4804 244190 4856 244196
rect 3516 238740 3568 238746
rect 3516 238682 3568 238688
rect 4804 221468 4856 221474
rect 4804 221410 4856 221416
rect 3516 215008 3568 215014
rect 3514 214976 3516 214985
rect 3568 214976 3570 214985
rect 3514 214911 3570 214920
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 3424 150408 3476 150414
rect 3424 150350 3476 150356
rect 3436 149841 3464 150350
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3240 137964 3292 137970
rect 3240 137906 3292 137912
rect 3252 136785 3280 137906
rect 3238 136776 3294 136785
rect 3238 136711 3294 136720
rect 3424 111784 3476 111790
rect 3424 111726 3476 111732
rect 3436 110673 3464 111726
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 4816 97782 4844 221410
rect 2780 97776 2832 97782
rect 2780 97718 2832 97724
rect 4804 97776 4856 97782
rect 4804 97718 4856 97724
rect 2792 97617 2820 97718
rect 2778 97608 2834 97617
rect 2778 97543 2834 97552
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 2778 61432 2834 61441
rect 2778 61367 2834 61376
rect 1676 8356 1728 8362
rect 1676 8298 1728 8304
rect 572 7608 624 7614
rect 572 7550 624 7556
rect 584 480 612 7550
rect 1688 480 1716 8298
rect 2792 3534 2820 61367
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3240 33788 3292 33794
rect 3240 33730 3292 33736
rect 3252 32473 3280 33730
rect 3238 32464 3294 32473
rect 3238 32399 3294 32408
rect 3516 20664 3568 20670
rect 3516 20606 3568 20612
rect 3424 19984 3476 19990
rect 3424 19926 3476 19932
rect 2872 10328 2924 10334
rect 2872 10270 2924 10276
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2884 480 2912 10270
rect 3436 6497 3464 19926
rect 3528 19417 3556 20606
rect 3514 19408 3570 19417
rect 3514 19343 3570 19352
rect 7656 11756 7708 11762
rect 7656 11698 7708 11704
rect 7472 9648 7524 9654
rect 7472 9590 7524 9596
rect 7484 8362 7512 9590
rect 7472 8356 7524 8362
rect 7472 8298 7524 8304
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 6460 4820 6512 4826
rect 6460 4762 6512 4768
rect 3700 3528 3752 3534
rect 3700 3470 3752 3476
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3712 354 3740 3470
rect 5264 2100 5316 2106
rect 5264 2042 5316 2048
rect 5276 480 5304 2042
rect 6472 480 6500 4762
rect 7668 480 7696 11698
rect 8220 9654 8248 292538
rect 8956 267714 8984 700266
rect 26884 670744 26936 670750
rect 26884 670686 26936 670692
rect 21364 632120 21416 632126
rect 21364 632062 21416 632068
rect 18604 553444 18656 553450
rect 18604 553386 18656 553392
rect 17224 409896 17276 409902
rect 17224 409838 17276 409844
rect 13084 357468 13136 357474
rect 13084 357410 13136 357416
rect 13096 338774 13124 357410
rect 13084 338768 13136 338774
rect 13084 338710 13136 338716
rect 8944 267708 8996 267714
rect 8944 267650 8996 267656
rect 8944 263628 8996 263634
rect 8944 263570 8996 263576
rect 8956 215014 8984 263570
rect 14464 256760 14516 256766
rect 14464 256702 14516 256708
rect 13084 253972 13136 253978
rect 13084 253914 13136 253920
rect 13096 235890 13124 253914
rect 13084 235884 13136 235890
rect 13084 235826 13136 235832
rect 13084 223100 13136 223106
rect 13084 223042 13136 223048
rect 8944 215008 8996 215014
rect 8944 214950 8996 214956
rect 13096 111790 13124 223042
rect 14476 137970 14504 256702
rect 17236 245614 17264 409838
rect 18616 263566 18644 553386
rect 21376 266354 21404 632062
rect 25504 448588 25556 448594
rect 25504 448530 25556 448536
rect 22100 318844 22152 318850
rect 22100 318786 22152 318792
rect 22112 318102 22140 318786
rect 22100 318096 22152 318102
rect 22100 318038 22152 318044
rect 25516 301510 25544 448530
rect 25504 301504 25556 301510
rect 25504 301446 25556 301452
rect 25504 289876 25556 289882
rect 25504 289818 25556 289824
rect 21364 266348 21416 266354
rect 21364 266290 21416 266296
rect 18604 263560 18656 263566
rect 18604 263502 18656 263508
rect 17224 245608 17276 245614
rect 17224 245550 17276 245556
rect 16580 240168 16632 240174
rect 16580 240110 16632 240116
rect 16592 237318 16620 240110
rect 16580 237312 16632 237318
rect 16580 237254 16632 237260
rect 25516 150414 25544 289818
rect 26896 286958 26924 670686
rect 39304 656940 39356 656946
rect 39304 656882 39356 656888
rect 36544 527196 36596 527202
rect 36544 527138 36596 527144
rect 31024 462392 31076 462398
rect 31024 462334 31076 462340
rect 26884 286952 26936 286958
rect 26884 286894 26936 286900
rect 31036 237250 31064 462334
rect 32404 294160 32456 294166
rect 32404 294102 32456 294108
rect 31024 237244 31076 237250
rect 31024 237186 31076 237192
rect 25504 150408 25556 150414
rect 25504 150350 25556 150356
rect 14464 137964 14516 137970
rect 14464 137906 14516 137912
rect 13084 111784 13136 111790
rect 13084 111726 13136 111732
rect 9680 73840 9732 73846
rect 9680 73782 9732 73788
rect 8298 57216 8354 57225
rect 8298 57151 8354 57160
rect 8312 16574 8340 57151
rect 8312 16546 8800 16574
rect 8208 9648 8260 9654
rect 8208 9590 8260 9596
rect 8772 480 8800 16546
rect 4038 354 4150 480
rect 3712 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 73782
rect 20720 68332 20772 68338
rect 20720 68274 20772 68280
rect 15200 54528 15252 54534
rect 15200 54470 15252 54476
rect 12440 51740 12492 51746
rect 12440 51682 12492 51688
rect 11058 22672 11114 22681
rect 11058 22607 11114 22616
rect 11072 3534 11100 22607
rect 11152 17264 11204 17270
rect 11152 17206 11204 17212
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 11164 480 11192 17206
rect 12452 16574 12480 51682
rect 13820 24132 13872 24138
rect 13820 24074 13872 24080
rect 13832 16574 13860 24074
rect 15212 16574 15240 54470
rect 17960 47592 18012 47598
rect 17960 47534 18012 47540
rect 16580 35216 16632 35222
rect 16580 35158 16632 35164
rect 16592 16574 16620 35158
rect 12452 16546 13584 16574
rect 13832 16546 14320 16574
rect 15212 16546 15976 16574
rect 16592 16546 17080 16574
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 11992 354 12020 3470
rect 13556 480 13584 16546
rect 12318 354 12430 480
rect 11992 326 12430 354
rect 12318 -960 12430 326
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 15948 480 15976 16546
rect 17052 480 17080 16546
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 47534
rect 19340 40724 19392 40730
rect 19340 40666 19392 40672
rect 19352 16574 19380 40666
rect 20732 16574 20760 68274
rect 26240 66904 26292 66910
rect 26240 66846 26292 66852
rect 24860 53100 24912 53106
rect 24860 53042 24912 53048
rect 23480 49020 23532 49026
rect 23480 48962 23532 48968
rect 22098 46200 22154 46209
rect 22098 46135 22154 46144
rect 22112 16574 22140 46135
rect 23492 16574 23520 48962
rect 24872 16574 24900 53042
rect 19352 16546 19472 16574
rect 20732 16546 21864 16574
rect 22112 16546 22600 16574
rect 23492 16546 24256 16574
rect 24872 16546 25360 16574
rect 19444 480 19472 16546
rect 20168 15904 20220 15910
rect 20168 15846 20220 15852
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20180 354 20208 15846
rect 21836 480 21864 16546
rect 20598 354 20710 480
rect 20180 326 20710 354
rect 20598 -960 20710 326
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 24228 480 24256 16546
rect 25332 480 25360 16546
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 66846
rect 28998 65512 29054 65521
rect 28998 65447 29054 65456
rect 27620 50380 27672 50386
rect 27620 50322 27672 50328
rect 27632 3534 27660 50322
rect 27712 32428 27764 32434
rect 27712 32370 27764 32376
rect 27620 3528 27672 3534
rect 27620 3470 27672 3476
rect 27724 480 27752 32370
rect 29012 16574 29040 65447
rect 31760 39364 31812 39370
rect 31760 39306 31812 39312
rect 31772 16574 31800 39306
rect 32416 20670 32444 294102
rect 36556 260846 36584 527138
rect 39316 309806 39344 656882
rect 39304 309800 39356 309806
rect 39304 309742 39356 309748
rect 39304 294024 39356 294030
rect 39304 293966 39356 293972
rect 36544 260840 36596 260846
rect 36544 260782 36596 260788
rect 39316 164218 39344 293966
rect 40052 238814 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 84292 703044 84344 703050
rect 84292 702986 84344 702992
rect 49608 702840 49660 702846
rect 49608 702782 49660 702788
rect 46204 618316 46256 618322
rect 46204 618258 46256 618264
rect 43444 397520 43496 397526
rect 43444 397462 43496 397468
rect 40040 238808 40092 238814
rect 40040 238750 40092 238756
rect 43456 237386 43484 397462
rect 45468 276072 45520 276078
rect 45468 276014 45520 276020
rect 44824 252612 44876 252618
rect 44824 252554 44876 252560
rect 43444 237380 43496 237386
rect 43444 237322 43496 237328
rect 43444 189780 43496 189786
rect 43444 189722 43496 189728
rect 39304 164212 39356 164218
rect 39304 164154 39356 164160
rect 34518 69592 34574 69601
rect 34518 69527 34574 69536
rect 33140 64184 33192 64190
rect 33140 64126 33192 64132
rect 32404 20664 32456 20670
rect 32404 20606 32456 20612
rect 33152 16574 33180 64126
rect 29012 16546 30144 16574
rect 31772 16546 31984 16574
rect 33152 16546 33640 16574
rect 28540 3528 28592 3534
rect 28540 3470 28592 3476
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28552 354 28580 3470
rect 30116 480 30144 16546
rect 31300 6180 31352 6186
rect 31300 6122 31352 6128
rect 31312 480 31340 6122
rect 28878 354 28990 480
rect 28552 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 31956 354 31984 16546
rect 33612 480 33640 16546
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 69527
rect 35900 62824 35952 62830
rect 35900 62766 35952 62772
rect 35912 3534 35940 62766
rect 40040 55956 40092 55962
rect 40040 55898 40092 55904
rect 38660 37936 38712 37942
rect 38660 37878 38712 37884
rect 37280 29640 37332 29646
rect 37280 29582 37332 29588
rect 35992 21412 36044 21418
rect 35992 21354 36044 21360
rect 35900 3528 35952 3534
rect 35900 3470 35952 3476
rect 36004 480 36032 21354
rect 37292 16574 37320 29582
rect 38672 16574 38700 37878
rect 40052 16574 40080 55898
rect 43456 45558 43484 189722
rect 44836 85542 44864 252554
rect 45480 222902 45508 276014
rect 46216 274650 46244 618258
rect 48964 292664 49016 292670
rect 48964 292606 49016 292612
rect 46848 280220 46900 280226
rect 46848 280162 46900 280168
rect 46204 274644 46256 274650
rect 46204 274586 46256 274592
rect 46204 267776 46256 267782
rect 46204 267718 46256 267724
rect 45468 222896 45520 222902
rect 45468 222838 45520 222844
rect 44824 85536 44876 85542
rect 44824 85478 44876 85484
rect 43444 45552 43496 45558
rect 43444 45494 43496 45500
rect 42800 36576 42852 36582
rect 42800 36518 42852 36524
rect 37292 16546 38424 16574
rect 38672 16546 39160 16574
rect 40052 16546 40264 16574
rect 36820 3528 36872 3534
rect 36820 3470 36872 3476
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36832 354 36860 3470
rect 38396 480 38424 16546
rect 37158 354 37270 480
rect 36832 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 41880 3596 41932 3602
rect 41880 3538 41932 3544
rect 41892 480 41920 3538
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 42812 354 42840 36518
rect 46216 33794 46244 267718
rect 46860 206281 46888 280162
rect 48228 274712 48280 274718
rect 48228 274654 48280 274660
rect 48240 218754 48268 274654
rect 48228 218748 48280 218754
rect 48228 218690 48280 218696
rect 46846 206272 46902 206281
rect 46846 206207 46902 206216
rect 48976 59362 49004 292606
rect 49620 247042 49648 702782
rect 63408 702772 63460 702778
rect 63408 702714 63460 702720
rect 55128 700460 55180 700466
rect 55128 700402 55180 700408
rect 53748 696244 53800 696250
rect 53748 696186 53800 696192
rect 50344 371272 50396 371278
rect 50344 371214 50396 371220
rect 49608 247036 49660 247042
rect 49608 246978 49660 246984
rect 50356 238610 50384 371214
rect 52368 284368 52420 284374
rect 52368 284310 52420 284316
rect 50896 277432 50948 277438
rect 50896 277374 50948 277380
rect 50344 238604 50396 238610
rect 50344 238546 50396 238552
rect 50908 225622 50936 277374
rect 50988 255332 51040 255338
rect 50988 255274 51040 255280
rect 50896 225616 50948 225622
rect 50896 225558 50948 225564
rect 51000 186998 51028 255274
rect 52380 197985 52408 284310
rect 53656 276140 53708 276146
rect 53656 276082 53708 276088
rect 53472 260908 53524 260914
rect 53472 260850 53524 260856
rect 53484 217326 53512 260850
rect 53564 256828 53616 256834
rect 53564 256770 53616 256776
rect 53472 217320 53524 217326
rect 53472 217262 53524 217268
rect 52366 197976 52422 197985
rect 52366 197911 52422 197920
rect 53576 195294 53604 256770
rect 53668 195430 53696 276082
rect 53760 242894 53788 696186
rect 55036 287088 55088 287094
rect 55036 287030 55088 287036
rect 54944 270564 54996 270570
rect 54944 270506 54996 270512
rect 53748 242888 53800 242894
rect 53748 242830 53800 242836
rect 54956 232529 54984 270506
rect 54942 232520 54998 232529
rect 54942 232455 54998 232464
rect 55048 209001 55076 287030
rect 55140 238542 55168 700402
rect 57888 700392 57940 700398
rect 57888 700334 57940 700340
rect 57244 278792 57296 278798
rect 57244 278734 57296 278740
rect 56508 277500 56560 277506
rect 56508 277442 56560 277448
rect 56416 263696 56468 263702
rect 56416 263638 56468 263644
rect 55128 238536 55180 238542
rect 55128 238478 55180 238484
rect 56428 215966 56456 263638
rect 56416 215960 56468 215966
rect 56416 215902 56468 215908
rect 55034 208992 55090 209001
rect 55034 208927 55090 208936
rect 56520 206310 56548 277442
rect 56508 206304 56560 206310
rect 56508 206246 56560 206252
rect 53656 195424 53708 195430
rect 53656 195366 53708 195372
rect 53564 195288 53616 195294
rect 53564 195230 53616 195236
rect 50988 186992 51040 186998
rect 50988 186934 51040 186940
rect 49698 75168 49754 75177
rect 49698 75103 49754 75112
rect 48964 59356 49016 59362
rect 48964 59298 49016 59304
rect 48320 58676 48372 58682
rect 48320 58618 48372 58624
rect 46204 33788 46256 33794
rect 46204 33730 46256 33736
rect 44180 31068 44232 31074
rect 44180 31010 44232 31016
rect 44192 6914 44220 31010
rect 44272 28280 44324 28286
rect 44272 28222 44324 28228
rect 44284 16574 44312 28222
rect 45560 18624 45612 18630
rect 45560 18566 45612 18572
rect 45572 16574 45600 18566
rect 48332 16574 48360 58618
rect 49712 16574 49740 75103
rect 53840 72480 53892 72486
rect 53840 72422 53892 72428
rect 52460 33788 52512 33794
rect 52460 33730 52512 33736
rect 44284 16546 45048 16574
rect 45572 16546 46704 16574
rect 48332 16546 48544 16574
rect 49712 16546 50200 16574
rect 44192 6886 44312 6914
rect 44284 480 44312 6886
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45020 354 45048 16546
rect 46676 480 46704 16546
rect 47400 13116 47452 13122
rect 47400 13058 47452 13064
rect 45438 354 45550 480
rect 45020 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 13058
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 50172 480 50200 16546
rect 52472 6914 52500 33730
rect 52552 26920 52604 26926
rect 52552 26862 52604 26868
rect 52564 16574 52592 26862
rect 53852 16574 53880 72422
rect 55220 55888 55272 55894
rect 55220 55830 55272 55836
rect 55232 16574 55260 55830
rect 56600 43444 56652 43450
rect 56600 43386 56652 43392
rect 56612 16574 56640 43386
rect 57256 19990 57284 278734
rect 57704 271924 57756 271930
rect 57704 271866 57756 271872
rect 57716 211818 57744 271866
rect 57900 271862 57928 700334
rect 59268 697604 59320 697610
rect 59268 697546 59320 697552
rect 59176 456816 59228 456822
rect 59176 456758 59228 456764
rect 57888 271856 57940 271862
rect 57888 271798 57940 271804
rect 57796 265668 57848 265674
rect 57796 265610 57848 265616
rect 57704 211812 57756 211818
rect 57704 211754 57756 211760
rect 57808 207641 57836 265610
rect 59084 258120 59136 258126
rect 59084 258062 59136 258068
rect 58992 248464 59044 248470
rect 58992 248406 59044 248412
rect 59004 217394 59032 248406
rect 58992 217388 59044 217394
rect 58992 217330 59044 217336
rect 57794 207632 57850 207641
rect 57794 207567 57850 207576
rect 59096 198014 59124 258062
rect 59188 241466 59216 456758
rect 59280 249762 59308 697546
rect 60648 285728 60700 285734
rect 60648 285670 60700 285676
rect 60556 269136 60608 269142
rect 60556 269078 60608 269084
rect 60464 258732 60516 258738
rect 60464 258674 60516 258680
rect 59268 249756 59320 249762
rect 59268 249698 59320 249704
rect 59268 247104 59320 247110
rect 59268 247046 59320 247052
rect 59176 241460 59228 241466
rect 59176 241402 59228 241408
rect 59280 199442 59308 247046
rect 60476 233986 60504 258674
rect 60464 233980 60516 233986
rect 60464 233922 60516 233928
rect 60568 202230 60596 269078
rect 60556 202224 60608 202230
rect 60556 202166 60608 202172
rect 59268 199436 59320 199442
rect 59268 199378 59320 199384
rect 59084 198008 59136 198014
rect 59084 197950 59136 197956
rect 60660 184249 60688 285670
rect 61936 274780 61988 274786
rect 61936 274722 61988 274728
rect 61752 255400 61804 255406
rect 61752 255342 61804 255348
rect 61764 227118 61792 255342
rect 61844 247172 61896 247178
rect 61844 247114 61896 247120
rect 61752 227112 61804 227118
rect 61752 227054 61804 227060
rect 61856 193905 61884 247114
rect 61948 217462 61976 274722
rect 62028 259480 62080 259486
rect 62028 259422 62080 259428
rect 61936 217456 61988 217462
rect 61936 217398 61988 217404
rect 61842 193896 61898 193905
rect 61842 193831 61898 193840
rect 60646 184240 60702 184249
rect 60646 184175 60702 184184
rect 62040 182850 62068 259422
rect 63316 258188 63368 258194
rect 63316 258130 63368 258136
rect 63132 249824 63184 249830
rect 63132 249766 63184 249772
rect 63144 204950 63172 249766
rect 63224 241528 63276 241534
rect 63224 241470 63276 241476
rect 63236 218822 63264 241470
rect 63224 218816 63276 218822
rect 63224 218758 63276 218764
rect 63328 213382 63356 258130
rect 63420 255270 63448 702714
rect 64144 565888 64196 565894
rect 64144 565830 64196 565836
rect 64156 267646 64184 565830
rect 67548 404388 67600 404394
rect 67548 404330 67600 404336
rect 67456 300960 67508 300966
rect 67456 300902 67508 300908
rect 66076 288448 66128 288454
rect 66076 288390 66128 288396
rect 64512 271992 64564 271998
rect 64512 271934 64564 271940
rect 64144 267640 64196 267646
rect 64144 267582 64196 267588
rect 63408 255264 63460 255270
rect 63408 255206 63460 255212
rect 63408 244316 63460 244322
rect 63408 244258 63460 244264
rect 63420 235414 63448 244258
rect 63408 235408 63460 235414
rect 63408 235350 63460 235356
rect 64524 224262 64552 271934
rect 64604 262268 64656 262274
rect 64604 262210 64656 262216
rect 64512 224256 64564 224262
rect 64512 224198 64564 224204
rect 63316 213376 63368 213382
rect 63316 213318 63368 213324
rect 63132 204944 63184 204950
rect 63132 204886 63184 204892
rect 64616 200870 64644 262210
rect 65892 252680 65944 252686
rect 65892 252622 65944 252628
rect 64696 249892 64748 249898
rect 64696 249834 64748 249840
rect 64604 200864 64656 200870
rect 64604 200806 64656 200812
rect 62028 182844 62080 182850
rect 62028 182786 62080 182792
rect 64708 180130 64736 249834
rect 65904 239970 65932 252622
rect 65984 242956 66036 242962
rect 65984 242898 66036 242904
rect 65892 239964 65944 239970
rect 65892 239906 65944 239912
rect 64788 235272 64840 235278
rect 64788 235214 64840 235220
rect 64696 180124 64748 180130
rect 64696 180066 64748 180072
rect 64694 125624 64750 125633
rect 64694 125559 64750 125568
rect 63408 122868 63460 122874
rect 63408 122810 63460 122816
rect 63420 84182 63448 122810
rect 64708 94897 64736 125559
rect 64694 94888 64750 94897
rect 64694 94823 64750 94832
rect 63408 84176 63460 84182
rect 63408 84118 63460 84124
rect 62120 71120 62172 71126
rect 62120 71062 62172 71068
rect 57980 68400 58032 68406
rect 57980 68342 58032 68348
rect 57244 19984 57296 19990
rect 57244 19926 57296 19932
rect 57992 16574 58020 68342
rect 59358 64152 59414 64161
rect 59358 64087 59414 64096
rect 52564 16546 53328 16574
rect 53852 16546 54984 16574
rect 55232 16546 56088 16574
rect 56612 16546 56824 16574
rect 57992 16546 58480 16574
rect 52472 6886 52592 6914
rect 51356 3460 51408 3466
rect 51356 3402 51408 3408
rect 51368 480 51396 3402
rect 52564 480 52592 6886
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53300 354 53328 16546
rect 54956 480 54984 16546
rect 56060 480 56088 16546
rect 53718 354 53830 480
rect 53300 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 58452 480 58480 16546
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 64087
rect 60740 25560 60792 25566
rect 60740 25502 60792 25508
rect 60752 16574 60780 25502
rect 62132 16574 62160 71062
rect 63500 44872 63552 44878
rect 63500 44814 63552 44820
rect 63512 16574 63540 44814
rect 60752 16546 60872 16574
rect 62132 16546 63264 16574
rect 63512 16546 64368 16574
rect 60844 480 60872 16546
rect 61568 15972 61620 15978
rect 61568 15914 61620 15920
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61580 354 61608 15914
rect 63236 480 63264 16546
rect 63500 8288 63552 8294
rect 63500 8230 63552 8236
rect 63512 7614 63540 8230
rect 63500 7608 63552 7614
rect 63500 7550 63552 7556
rect 64340 480 64368 16546
rect 64800 8294 64828 235214
rect 65996 182918 66024 242898
rect 66088 214674 66116 288390
rect 67468 285705 67496 300902
rect 67454 285696 67510 285705
rect 67454 285631 67510 285640
rect 67560 282985 67588 404330
rect 68928 323604 68980 323610
rect 68928 323546 68980 323552
rect 68744 299600 68796 299606
rect 68744 299542 68796 299548
rect 68560 295452 68612 295458
rect 68560 295394 68612 295400
rect 67638 291136 67694 291145
rect 67638 291071 67694 291080
rect 67652 289882 67680 291071
rect 67640 289876 67692 289882
rect 67640 289818 67692 289824
rect 68572 289626 68600 295394
rect 68756 289785 68784 299542
rect 68834 296848 68890 296857
rect 68834 296783 68890 296792
rect 68848 290465 68876 296783
rect 68834 290456 68890 290465
rect 68834 290391 68890 290400
rect 68742 289776 68798 289785
rect 68742 289711 68798 289720
rect 68572 289598 68692 289626
rect 68560 289536 68612 289542
rect 68560 289478 68612 289484
rect 68190 289096 68246 289105
rect 68190 289031 68246 289040
rect 68204 288454 68232 289031
rect 68192 288448 68244 288454
rect 68192 288390 68244 288396
rect 67638 287736 67694 287745
rect 67638 287671 67694 287680
rect 67652 287094 67680 287671
rect 67640 287088 67692 287094
rect 67640 287030 67692 287036
rect 67730 287056 67786 287065
rect 67730 286991 67786 287000
rect 67640 286952 67692 286958
rect 67640 286894 67692 286900
rect 67652 286385 67680 286894
rect 67638 286376 67694 286385
rect 67638 286311 67694 286320
rect 67744 285734 67772 286991
rect 67732 285728 67784 285734
rect 67732 285670 67784 285676
rect 67640 284368 67692 284374
rect 67638 284336 67640 284345
rect 67692 284336 67694 284345
rect 67638 284271 67694 284280
rect 67546 282976 67602 282985
rect 67546 282911 67602 282920
rect 68572 281625 68600 289478
rect 68664 289354 68692 289598
rect 68940 289542 68968 323546
rect 69112 311160 69164 311166
rect 69112 311102 69164 311108
rect 69020 307080 69072 307086
rect 69020 307022 69072 307028
rect 68928 289536 68980 289542
rect 68928 289478 68980 289484
rect 68664 289326 68876 289354
rect 68848 283665 68876 289326
rect 68834 283656 68890 283665
rect 68834 283591 68890 283600
rect 68558 281616 68614 281625
rect 68558 281551 68614 281560
rect 67638 280936 67694 280945
rect 67638 280871 67694 280880
rect 67652 280226 67680 280871
rect 68374 280256 68430 280265
rect 67640 280220 67692 280226
rect 68374 280191 68430 280200
rect 67640 280162 67692 280168
rect 67638 279576 67694 279585
rect 67638 279511 67694 279520
rect 67652 278798 67680 279511
rect 67640 278792 67692 278798
rect 67640 278734 67692 278740
rect 67730 278216 67786 278225
rect 67730 278151 67786 278160
rect 67638 277536 67694 277545
rect 67638 277471 67640 277480
rect 67692 277471 67694 277480
rect 67640 277442 67692 277448
rect 67744 277438 67772 278151
rect 67732 277432 67784 277438
rect 67732 277374 67784 277380
rect 67730 276856 67786 276865
rect 67730 276791 67786 276800
rect 67638 276176 67694 276185
rect 67744 276146 67772 276791
rect 67638 276111 67694 276120
rect 67732 276140 67784 276146
rect 67652 276078 67680 276111
rect 67732 276082 67784 276088
rect 67640 276072 67692 276078
rect 67640 276014 67692 276020
rect 67730 275496 67786 275505
rect 67730 275431 67786 275440
rect 67638 274816 67694 274825
rect 67638 274751 67640 274760
rect 67692 274751 67694 274760
rect 67640 274722 67692 274728
rect 67744 274718 67772 275431
rect 67732 274712 67784 274718
rect 67732 274654 67784 274660
rect 67640 274644 67692 274650
rect 67640 274586 67692 274592
rect 67652 274145 67680 274586
rect 67638 274136 67694 274145
rect 67638 274071 67694 274080
rect 68006 273456 68062 273465
rect 68006 273391 68062 273400
rect 68020 273290 68048 273391
rect 66168 273284 66220 273290
rect 66168 273226 66220 273232
rect 68008 273284 68060 273290
rect 68008 273226 68060 273232
rect 66076 214668 66128 214674
rect 66076 214610 66128 214616
rect 65984 182912 66036 182918
rect 65984 182854 66036 182860
rect 66180 181490 66208 273226
rect 67822 272776 67878 272785
rect 67822 272711 67878 272720
rect 67638 272096 67694 272105
rect 67638 272031 67694 272040
rect 67652 271998 67680 272031
rect 67640 271992 67692 271998
rect 67640 271934 67692 271940
rect 67836 271930 67864 272711
rect 67824 271924 67876 271930
rect 67824 271866 67876 271872
rect 67732 271856 67784 271862
rect 67732 271798 67784 271804
rect 67638 271416 67694 271425
rect 67638 271351 67694 271360
rect 67652 270570 67680 271351
rect 67744 270745 67772 271798
rect 67730 270736 67786 270745
rect 67730 270671 67786 270680
rect 67640 270564 67692 270570
rect 67640 270506 67692 270512
rect 67638 270056 67694 270065
rect 67638 269991 67694 270000
rect 67652 269142 67680 269991
rect 68282 269376 68338 269385
rect 68282 269311 68338 269320
rect 67640 269136 67692 269142
rect 67640 269078 67692 269084
rect 67546 268696 67602 268705
rect 67546 268631 67602 268640
rect 67362 261216 67418 261225
rect 67362 261151 67418 261160
rect 67376 232558 67404 261151
rect 67454 251696 67510 251705
rect 67454 251631 67510 251640
rect 67364 232552 67416 232558
rect 67364 232494 67416 232500
rect 67468 209098 67496 251631
rect 67560 211886 67588 268631
rect 67638 268016 67694 268025
rect 67638 267951 67694 267960
rect 67652 267782 67680 267951
rect 67640 267776 67692 267782
rect 67640 267718 67692 267724
rect 67732 267708 67784 267714
rect 67732 267650 67784 267656
rect 67640 267640 67692 267646
rect 67640 267582 67692 267588
rect 67652 267345 67680 267582
rect 67638 267336 67694 267345
rect 67638 267271 67694 267280
rect 67744 266665 67772 267650
rect 67730 266656 67786 266665
rect 67730 266591 67786 266600
rect 67640 266348 67692 266354
rect 67640 266290 67692 266296
rect 67652 265305 67680 266290
rect 67822 265976 67878 265985
rect 67822 265911 67878 265920
rect 67638 265296 67694 265305
rect 67638 265231 67694 265240
rect 67730 264616 67786 264625
rect 67730 264551 67786 264560
rect 67638 263936 67694 263945
rect 67638 263871 67694 263880
rect 67652 263702 67680 263871
rect 67640 263696 67692 263702
rect 67640 263638 67692 263644
rect 67744 263634 67772 264551
rect 67732 263628 67784 263634
rect 67732 263570 67784 263576
rect 67640 263560 67692 263566
rect 67640 263502 67692 263508
rect 67652 263265 67680 263502
rect 67638 263256 67694 263265
rect 67638 263191 67694 263200
rect 67638 262576 67694 262585
rect 67638 262511 67694 262520
rect 67652 262274 67680 262511
rect 67640 262268 67692 262274
rect 67640 262210 67692 262216
rect 67730 261896 67786 261905
rect 67730 261831 67786 261840
rect 67744 260914 67772 261831
rect 67732 260908 67784 260914
rect 67732 260850 67784 260856
rect 67640 260840 67692 260846
rect 67640 260782 67692 260788
rect 67652 260545 67680 260782
rect 67638 260536 67694 260545
rect 67638 260471 67694 260480
rect 67638 259856 67694 259865
rect 67638 259791 67694 259800
rect 67652 259486 67680 259791
rect 67640 259480 67692 259486
rect 67640 259422 67692 259428
rect 67730 259176 67786 259185
rect 67730 259111 67786 259120
rect 67638 258496 67694 258505
rect 67638 258431 67694 258440
rect 67652 258194 67680 258431
rect 67640 258188 67692 258194
rect 67640 258130 67692 258136
rect 67744 258126 67772 259111
rect 67836 258738 67864 265911
rect 67824 258732 67876 258738
rect 67824 258674 67876 258680
rect 67732 258120 67784 258126
rect 67732 258062 67784 258068
rect 67730 257816 67786 257825
rect 67730 257751 67786 257760
rect 67638 257136 67694 257145
rect 67638 257071 67694 257080
rect 67652 256834 67680 257071
rect 67640 256828 67692 256834
rect 67640 256770 67692 256776
rect 67744 256766 67772 257751
rect 67732 256760 67784 256766
rect 67732 256702 67784 256708
rect 67638 256456 67694 256465
rect 67638 256391 67694 256400
rect 67652 255406 67680 256391
rect 67730 255776 67786 255785
rect 67730 255711 67786 255720
rect 67640 255400 67692 255406
rect 67640 255342 67692 255348
rect 67744 255338 67772 255711
rect 67732 255332 67784 255338
rect 67732 255274 67784 255280
rect 67640 255264 67692 255270
rect 67640 255206 67692 255212
rect 67652 255105 67680 255206
rect 67638 255096 67694 255105
rect 67638 255031 67694 255040
rect 67638 253736 67694 253745
rect 67638 253671 67694 253680
rect 67652 252618 67680 253671
rect 68098 253056 68154 253065
rect 68098 252991 68154 253000
rect 68112 252686 68140 252991
rect 68100 252680 68152 252686
rect 68100 252622 68152 252628
rect 67640 252612 67692 252618
rect 67640 252554 67692 252560
rect 67638 251016 67694 251025
rect 67638 250951 67694 250960
rect 67652 249898 67680 250951
rect 67730 250336 67786 250345
rect 67730 250271 67786 250280
rect 67640 249892 67692 249898
rect 67640 249834 67692 249840
rect 67744 249830 67772 250271
rect 67732 249824 67784 249830
rect 67732 249766 67784 249772
rect 67640 249756 67692 249762
rect 67640 249698 67692 249704
rect 67652 249665 67680 249698
rect 67638 249656 67694 249665
rect 67638 249591 67694 249600
rect 67638 248976 67694 248985
rect 67638 248911 67694 248920
rect 67652 248470 67680 248911
rect 67640 248464 67692 248470
rect 67640 248406 67692 248412
rect 67638 248296 67694 248305
rect 67638 248231 67694 248240
rect 67652 247178 67680 248231
rect 67730 247616 67786 247625
rect 67730 247551 67786 247560
rect 67640 247172 67692 247178
rect 67640 247114 67692 247120
rect 67744 247110 67772 247551
rect 67732 247104 67784 247110
rect 67732 247046 67784 247052
rect 67640 247036 67692 247042
rect 67640 246978 67692 246984
rect 67652 246945 67680 246978
rect 67638 246936 67694 246945
rect 67638 246871 67694 246880
rect 68296 245721 68324 269311
rect 68388 265674 68416 280191
rect 69032 278905 69060 307022
rect 69124 288425 69152 311102
rect 71792 308446 71820 702986
rect 80704 702500 80756 702506
rect 80704 702442 80756 702448
rect 77300 315308 77352 315314
rect 77300 315250 77352 315256
rect 71780 308440 71832 308446
rect 71780 308382 71832 308388
rect 75920 306400 75972 306406
rect 77312 306374 77340 315250
rect 75972 306348 76144 306374
rect 75920 306346 76144 306348
rect 77312 306346 77984 306374
rect 75920 306342 75972 306346
rect 75366 302288 75422 302297
rect 75366 302223 75422 302232
rect 70952 301504 71004 301510
rect 70952 301446 71004 301452
rect 73528 301504 73580 301510
rect 73528 301446 73580 301452
rect 70032 296948 70084 296954
rect 70032 296890 70084 296896
rect 69480 294092 69532 294098
rect 69480 294034 69532 294040
rect 69492 291854 69520 294034
rect 70044 291924 70072 296890
rect 70676 296744 70728 296750
rect 70676 296686 70728 296692
rect 70688 291924 70716 296686
rect 70964 291938 70992 301446
rect 71780 299532 71832 299538
rect 71780 299474 71832 299480
rect 71792 291938 71820 299474
rect 72608 298784 72660 298790
rect 72608 298726 72660 298732
rect 70964 291910 71346 291938
rect 71792 291910 71990 291938
rect 72620 291924 72648 298726
rect 73252 294636 73304 294642
rect 73252 294578 73304 294584
rect 73264 291924 73292 294578
rect 73540 291938 73568 301446
rect 74540 298376 74592 298382
rect 74540 298318 74592 298324
rect 73540 291910 73922 291938
rect 74552 291924 74580 298318
rect 75184 298308 75236 298314
rect 75184 298250 75236 298256
rect 75196 291924 75224 298250
rect 75380 291938 75408 302223
rect 76116 291938 76144 306346
rect 77116 295656 77168 295662
rect 77116 295598 77168 295604
rect 75380 291910 75854 291938
rect 76116 291910 76498 291938
rect 77128 291924 77156 295598
rect 77760 294024 77812 294030
rect 77760 293966 77812 293972
rect 77772 291924 77800 293966
rect 77956 291938 77984 306346
rect 79232 302320 79284 302326
rect 79232 302262 79284 302268
rect 78772 293956 78824 293962
rect 78772 293898 78824 293904
rect 78784 291938 78812 293898
rect 79244 291938 79272 302262
rect 80518 299568 80574 299577
rect 80518 299503 80574 299512
rect 80334 294128 80390 294137
rect 80334 294063 80390 294072
rect 77956 291910 78430 291938
rect 78784 291910 79074 291938
rect 79244 291910 79718 291938
rect 80348 291924 80376 294063
rect 80532 291938 80560 299503
rect 80716 294030 80744 702442
rect 82084 700324 82136 700330
rect 82084 700266 82136 700272
rect 80796 351960 80848 351966
rect 80796 351902 80848 351908
rect 80808 301510 80836 351902
rect 82096 303618 82124 700266
rect 82084 303612 82136 303618
rect 82084 303554 82136 303560
rect 80796 301504 80848 301510
rect 80796 301446 80848 301452
rect 81624 298240 81676 298246
rect 81624 298182 81676 298188
rect 80704 294024 80756 294030
rect 80704 293966 80756 293972
rect 80532 291910 81006 291938
rect 81636 291924 81664 298182
rect 82268 295588 82320 295594
rect 82268 295530 82320 295536
rect 82280 291924 82308 295530
rect 84200 295520 84252 295526
rect 84200 295462 84252 295468
rect 82912 294228 82964 294234
rect 82912 294170 82964 294176
rect 82924 291924 82952 294170
rect 83556 292868 83608 292874
rect 83556 292810 83608 292816
rect 83568 291924 83596 292810
rect 84212 291924 84240 295462
rect 84304 294030 84332 702986
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 88352 334626 88380 702406
rect 105464 700466 105492 703520
rect 107660 702976 107712 702982
rect 107660 702918 107712 702924
rect 106280 702704 106332 702710
rect 106280 702646 106332 702652
rect 105452 700460 105504 700466
rect 105452 700402 105504 700408
rect 102784 563100 102836 563106
rect 102784 563042 102836 563048
rect 100024 501016 100076 501022
rect 100024 500958 100076 500964
rect 93124 418192 93176 418198
rect 93124 418134 93176 418140
rect 88340 334620 88392 334626
rect 88340 334562 88392 334568
rect 91100 319456 91152 319462
rect 91100 319398 91152 319404
rect 90272 303680 90324 303686
rect 90272 303622 90324 303628
rect 84476 303612 84528 303618
rect 84476 303554 84528 303560
rect 84292 294024 84344 294030
rect 84292 293966 84344 293972
rect 84488 291938 84516 303554
rect 86408 300892 86460 300898
rect 86408 300834 86460 300840
rect 86132 297016 86184 297022
rect 86132 296958 86184 296964
rect 85212 294024 85264 294030
rect 85212 293966 85264 293972
rect 85224 291938 85252 293966
rect 84488 291910 84870 291938
rect 85224 291910 85514 291938
rect 86144 291924 86172 296958
rect 86420 291938 86448 300834
rect 87696 299668 87748 299674
rect 87696 299610 87748 299616
rect 87420 294704 87472 294710
rect 87420 294646 87472 294652
rect 86420 291910 86802 291938
rect 87432 291924 87460 294646
rect 87708 291938 87736 299610
rect 89996 298512 90048 298518
rect 89996 298454 90048 298460
rect 89352 296880 89404 296886
rect 89352 296822 89404 296828
rect 88708 296812 88760 296818
rect 88708 296754 88760 296760
rect 87708 291910 88090 291938
rect 88720 291924 88748 296754
rect 89364 291924 89392 296822
rect 90008 291924 90036 298454
rect 90284 291938 90312 303622
rect 91112 291938 91140 319398
rect 93136 315314 93164 418134
rect 98000 338768 98052 338774
rect 98000 338710 98052 338716
rect 93952 317552 94004 317558
rect 93952 317494 94004 317500
rect 93124 315308 93176 315314
rect 93124 315250 93176 315256
rect 93216 298444 93268 298450
rect 93216 298386 93268 298392
rect 91928 294296 91980 294302
rect 91928 294238 91980 294244
rect 90284 291910 90666 291938
rect 91112 291910 91310 291938
rect 91940 291924 91968 294238
rect 92572 294092 92624 294098
rect 92572 294034 92624 294040
rect 92584 291924 92612 294034
rect 93228 291924 93256 298386
rect 93964 294030 93992 317494
rect 94136 312588 94188 312594
rect 94136 312530 94188 312536
rect 93952 294024 94004 294030
rect 93952 293966 94004 293972
rect 93860 292936 93912 292942
rect 93860 292878 93912 292884
rect 93872 291924 93900 292878
rect 94148 291938 94176 312530
rect 95790 294264 95846 294273
rect 95790 294199 95846 294208
rect 94780 294024 94832 294030
rect 94780 293966 94832 293972
rect 94792 291938 94820 293966
rect 94148 291910 94530 291938
rect 94792 291910 95174 291938
rect 95804 291924 95832 294199
rect 97080 292664 97132 292670
rect 97080 292606 97132 292612
rect 97724 292664 97776 292670
rect 97724 292606 97776 292612
rect 96436 292596 96488 292602
rect 96436 292538 96488 292544
rect 96448 291924 96476 292538
rect 97092 291924 97120 292606
rect 97736 291924 97764 292606
rect 98012 291938 98040 338710
rect 100036 312594 100064 500958
rect 102796 317558 102824 563042
rect 103796 334620 103848 334626
rect 103796 334562 103848 334568
rect 102784 317552 102836 317558
rect 102784 317494 102836 317500
rect 100024 312588 100076 312594
rect 100024 312530 100076 312536
rect 98092 307828 98144 307834
rect 98092 307770 98144 307776
rect 98104 306374 98132 307770
rect 103808 306374 103836 334562
rect 106292 306374 106320 702646
rect 107672 306374 107700 702918
rect 129004 702908 129056 702914
rect 129004 702850 129056 702856
rect 124864 702636 124916 702642
rect 124864 702578 124916 702584
rect 116584 579692 116636 579698
rect 116584 579634 116636 579640
rect 111064 474768 111116 474774
rect 111064 474710 111116 474716
rect 111076 322250 111104 474710
rect 111064 322244 111116 322250
rect 111064 322186 111116 322192
rect 115940 318096 115992 318102
rect 115940 318038 115992 318044
rect 114560 308440 114612 308446
rect 114560 308382 114612 308388
rect 114572 306374 114600 308382
rect 115952 306374 115980 318038
rect 98104 306346 98592 306374
rect 103808 306346 104480 306374
rect 106292 306346 107056 306374
rect 107672 306346 108344 306374
rect 114572 306346 114784 306374
rect 115952 306346 116072 306374
rect 98564 291938 98592 306346
rect 102140 303816 102192 303822
rect 102140 303758 102192 303764
rect 99654 295488 99710 295497
rect 99654 295423 99710 295432
rect 98012 291910 98394 291938
rect 98564 291910 99038 291938
rect 99668 291924 99696 295423
rect 100944 292800 100996 292806
rect 100944 292742 100996 292748
rect 100956 291924 100984 292742
rect 101586 292632 101642 292641
rect 101586 292567 101642 292576
rect 101600 291924 101628 292567
rect 102152 291938 102180 303758
rect 102416 303748 102468 303754
rect 102416 303690 102468 303696
rect 102428 291938 102456 303690
rect 103520 292732 103572 292738
rect 103520 292674 103572 292680
rect 102152 291910 102258 291938
rect 102428 291910 102902 291938
rect 103532 291924 103560 292674
rect 104162 292632 104218 292641
rect 104162 292567 104218 292576
rect 104176 291924 104204 292567
rect 104452 291938 104480 306346
rect 106096 298172 106148 298178
rect 106096 298114 106148 298120
rect 105450 292768 105506 292777
rect 105450 292703 105506 292712
rect 104452 291910 104834 291938
rect 105464 291924 105492 292703
rect 106108 291924 106136 298114
rect 106740 294364 106792 294370
rect 106740 294306 106792 294312
rect 106752 291924 106780 294306
rect 107028 291938 107056 306346
rect 108210 291952 108266 291961
rect 107028 291910 107410 291938
rect 108054 291910 108210 291938
rect 108316 291938 108344 306346
rect 112444 305040 112496 305046
rect 112444 304982 112496 304988
rect 112168 302252 112220 302258
rect 112168 302194 112220 302200
rect 110420 299736 110472 299742
rect 110420 299678 110472 299684
rect 109960 295384 110012 295390
rect 109960 295326 110012 295332
rect 109316 292596 109368 292602
rect 109316 292538 109368 292544
rect 108316 291910 108698 291938
rect 109328 291924 109356 292538
rect 109972 291924 110000 295326
rect 110432 291938 110460 299678
rect 111248 295724 111300 295730
rect 111248 295666 111300 295672
rect 110432 291910 110630 291938
rect 111260 291924 111288 295666
rect 111798 295352 111854 295361
rect 111798 295287 111854 295296
rect 111812 294642 111840 295287
rect 111800 294636 111852 294642
rect 111800 294578 111852 294584
rect 111892 294024 111944 294030
rect 111892 293966 111944 293972
rect 111904 291924 111932 293966
rect 112180 291938 112208 302194
rect 112456 294710 112484 304982
rect 114468 297084 114520 297090
rect 114468 297026 114520 297032
rect 112444 294704 112496 294710
rect 112444 294646 112496 294652
rect 113824 294432 113876 294438
rect 113824 294374 113876 294380
rect 113178 293992 113234 294001
rect 113178 293927 113234 293936
rect 112180 291910 112562 291938
rect 113192 291924 113220 293927
rect 113836 291924 113864 294374
rect 114480 291924 114508 297026
rect 114756 291938 114784 306346
rect 116044 291938 116072 306346
rect 116596 293185 116624 579634
rect 123484 430636 123536 430642
rect 123484 430578 123536 430584
rect 117964 345092 118016 345098
rect 117964 345034 118016 345040
rect 117976 301578 118004 345034
rect 120172 326392 120224 326398
rect 120172 326334 120224 326340
rect 120080 313948 120132 313954
rect 120080 313890 120132 313896
rect 119804 305108 119856 305114
rect 119804 305050 119856 305056
rect 117964 301572 118016 301578
rect 117964 301514 118016 301520
rect 119160 301572 119212 301578
rect 119160 301514 119212 301520
rect 118424 294432 118476 294438
rect 118424 294374 118476 294380
rect 117688 294160 117740 294166
rect 117688 294102 117740 294108
rect 116582 293176 116638 293185
rect 116582 293111 116638 293120
rect 114756 291910 115138 291938
rect 115782 291922 115888 291938
rect 115782 291916 115900 291922
rect 115782 291910 115848 291916
rect 108210 291887 108266 291896
rect 116044 291910 116426 291938
rect 117070 291922 117268 291938
rect 117700 291924 117728 294102
rect 118436 294098 118464 294374
rect 118332 294092 118384 294098
rect 118332 294034 118384 294040
rect 118424 294092 118476 294098
rect 118424 294034 118476 294040
rect 118344 291924 118372 294034
rect 119172 291938 119200 301514
rect 119002 291922 119108 291938
rect 117070 291916 117280 291922
rect 117070 291910 117228 291916
rect 115848 291858 115900 291864
rect 119002 291916 119120 291922
rect 119002 291910 119068 291916
rect 117228 291858 117280 291864
rect 119172 291910 119646 291938
rect 119068 291858 119120 291864
rect 69480 291848 69532 291854
rect 69480 291790 69532 291796
rect 69754 291272 69810 291281
rect 69754 291207 69756 291216
rect 69808 291207 69810 291216
rect 69756 291178 69808 291184
rect 69110 288416 69166 288425
rect 69110 288351 69166 288360
rect 119816 286793 119844 305050
rect 119896 291916 119948 291922
rect 119896 291858 119948 291864
rect 119908 290601 119936 291858
rect 119894 290592 119950 290601
rect 119894 290527 119950 290536
rect 119802 286784 119858 286793
rect 119802 286719 119858 286728
rect 69018 278896 69074 278905
rect 69018 278831 69074 278840
rect 68376 265668 68428 265674
rect 68376 265610 68428 265616
rect 119804 251864 119856 251870
rect 119804 251806 119856 251812
rect 69018 246256 69074 246265
rect 69018 246191 69074 246200
rect 68282 245712 68338 245721
rect 68282 245647 68338 245656
rect 67640 245608 67692 245614
rect 67638 245576 67640 245585
rect 67692 245576 67694 245585
rect 67638 245511 67694 245520
rect 67638 244896 67694 244905
rect 67638 244831 67694 244840
rect 67652 244322 67680 244831
rect 67640 244316 67692 244322
rect 67640 244258 67692 244264
rect 67732 244248 67784 244254
rect 67732 244190 67784 244196
rect 67822 244216 67878 244225
rect 67744 243545 67772 244190
rect 67822 244151 67878 244160
rect 67730 243536 67786 243545
rect 67730 243471 67786 243480
rect 67836 242962 67864 244151
rect 67824 242956 67876 242962
rect 67824 242898 67876 242904
rect 67640 242888 67692 242894
rect 67638 242856 67640 242865
rect 67692 242856 67694 242865
rect 67638 242791 67694 242800
rect 67730 242176 67786 242185
rect 67730 242111 67786 242120
rect 67744 241534 67772 242111
rect 67732 241528 67784 241534
rect 67638 241496 67694 241505
rect 67732 241470 67784 241476
rect 67638 241431 67640 241440
rect 67692 241431 67694 241440
rect 67640 241402 67692 241408
rect 67548 211880 67600 211886
rect 67548 211822 67600 211828
rect 67456 209092 67508 209098
rect 67456 209034 67508 209040
rect 69032 195362 69060 246191
rect 119816 240242 119844 251806
rect 120092 247625 120120 313890
rect 120184 261225 120212 326334
rect 121460 322244 121512 322250
rect 121460 322186 121512 322192
rect 120722 293992 120778 294001
rect 120722 293927 120778 293936
rect 120264 292936 120316 292942
rect 120264 292878 120316 292884
rect 120276 289134 120304 292878
rect 120264 289128 120316 289134
rect 120264 289070 120316 289076
rect 120170 261216 120226 261225
rect 120170 261151 120226 261160
rect 120170 251016 120226 251025
rect 120170 250951 120226 250960
rect 120078 247616 120134 247625
rect 120078 247551 120134 247560
rect 119804 240236 119856 240242
rect 119804 240178 119856 240184
rect 119896 240168 119948 240174
rect 69124 240094 70058 240122
rect 119646 240116 119896 240122
rect 119646 240110 119948 240116
rect 69124 228410 69152 240094
rect 70582 239864 70638 239873
rect 70582 239799 70638 239808
rect 70596 239426 70624 239799
rect 70584 239420 70636 239426
rect 70584 239362 70636 239368
rect 69112 228404 69164 228410
rect 69112 228346 69164 228352
rect 70688 219434 70716 240108
rect 71044 239964 71096 239970
rect 71044 239906 71096 239912
rect 71056 220114 71084 239906
rect 71332 237454 71360 240108
rect 71320 237448 71372 237454
rect 71320 237390 71372 237396
rect 71044 220108 71096 220114
rect 71044 220050 71096 220056
rect 71976 219434 72004 240108
rect 72620 238678 72648 240108
rect 72608 238672 72660 238678
rect 72608 238614 72660 238620
rect 73160 233028 73212 233034
rect 73160 232970 73212 232976
rect 70412 219406 70716 219434
rect 71792 219406 72004 219434
rect 69020 195356 69072 195362
rect 69020 195298 69072 195304
rect 66168 181484 66220 181490
rect 66168 181426 66220 181432
rect 70412 178702 70440 219406
rect 71792 180198 71820 219406
rect 73172 182986 73200 232970
rect 73264 186969 73292 240108
rect 73908 233034 73936 240108
rect 74552 238066 74580 240108
rect 75196 238754 75224 240108
rect 74920 238726 75224 238754
rect 74540 238060 74592 238066
rect 74540 238002 74592 238008
rect 73896 233028 73948 233034
rect 73896 232970 73948 232976
rect 74920 220250 74948 238726
rect 75184 237448 75236 237454
rect 75184 237390 75236 237396
rect 74908 220244 74960 220250
rect 74908 220186 74960 220192
rect 75196 193866 75224 237390
rect 75840 233238 75868 240108
rect 76484 238754 76512 240108
rect 75932 238726 76512 238754
rect 75828 233232 75880 233238
rect 75828 233174 75880 233180
rect 75184 193860 75236 193866
rect 75184 193802 75236 193808
rect 75932 191146 75960 238726
rect 77128 224233 77156 240108
rect 77772 238754 77800 240108
rect 77312 238726 77800 238754
rect 77114 224224 77170 224233
rect 77114 224159 77170 224168
rect 75920 191140 75972 191146
rect 75920 191082 75972 191088
rect 77312 189689 77340 238726
rect 78416 219434 78444 240108
rect 79060 237658 79088 240108
rect 79048 237652 79100 237658
rect 79048 237594 79100 237600
rect 79704 219434 79732 240108
rect 80060 229764 80112 229770
rect 80060 229706 80112 229712
rect 77404 219406 78444 219434
rect 78692 219406 79732 219434
rect 77404 196654 77432 219406
rect 78692 214606 78720 219406
rect 78680 214600 78732 214606
rect 78680 214542 78732 214548
rect 77392 196648 77444 196654
rect 77392 196590 77444 196596
rect 77298 189680 77354 189689
rect 77298 189615 77354 189624
rect 73250 186960 73306 186969
rect 73250 186895 73306 186904
rect 80072 185638 80100 229706
rect 80348 225690 80376 240108
rect 80704 237652 80756 237658
rect 80704 237594 80756 237600
rect 80336 225684 80388 225690
rect 80336 225626 80388 225632
rect 80716 220182 80744 237594
rect 80992 229770 81020 240108
rect 81636 231810 81664 240108
rect 82280 237386 82308 240108
rect 82268 237380 82320 237386
rect 82268 237322 82320 237328
rect 81624 231804 81676 231810
rect 81624 231746 81676 231752
rect 82924 229906 82952 240108
rect 82912 229900 82964 229906
rect 82912 229842 82964 229848
rect 80980 229764 81032 229770
rect 80980 229706 81032 229712
rect 83568 221474 83596 240108
rect 84212 238754 84240 240108
rect 84212 238726 84424 238754
rect 84292 233912 84344 233918
rect 84292 233854 84344 233860
rect 84108 231872 84160 231878
rect 84160 231826 84240 231854
rect 84108 231814 84160 231820
rect 83556 221468 83608 221474
rect 83556 221410 83608 221416
rect 80704 220176 80756 220182
rect 80704 220118 80756 220124
rect 84212 192506 84240 231826
rect 84304 210458 84332 233854
rect 84396 221513 84424 238726
rect 84856 231878 84884 240108
rect 85500 233918 85528 240108
rect 85488 233912 85540 233918
rect 85488 233854 85540 233860
rect 84844 231872 84896 231878
rect 84844 231814 84896 231820
rect 86144 229770 86172 240108
rect 86224 239420 86276 239426
rect 86224 239362 86276 239368
rect 86132 229764 86184 229770
rect 86132 229706 86184 229712
rect 84382 221504 84438 221513
rect 84382 221439 84438 221448
rect 86236 216034 86264 239362
rect 86788 238746 86816 240108
rect 86776 238740 86828 238746
rect 86776 238682 86828 238688
rect 87432 219434 87460 240108
rect 88076 229838 88104 240108
rect 88064 229832 88116 229838
rect 88064 229774 88116 229780
rect 88720 219434 88748 240108
rect 89364 238542 89392 240108
rect 90008 238754 90036 240108
rect 89732 238726 90036 238754
rect 89352 238536 89404 238542
rect 89352 238478 89404 238484
rect 86972 219406 87460 219434
rect 88444 219406 88748 219434
rect 86224 216028 86276 216034
rect 86224 215970 86276 215976
rect 84292 210452 84344 210458
rect 84292 210394 84344 210400
rect 86972 199646 87000 219406
rect 86960 199640 87012 199646
rect 86960 199582 87012 199588
rect 84200 192500 84252 192506
rect 84200 192442 84252 192448
rect 88444 188358 88472 219406
rect 89732 192574 89760 238726
rect 90652 219434 90680 240108
rect 91296 238513 91324 240108
rect 91282 238504 91338 238513
rect 91282 238439 91338 238448
rect 91940 237386 91968 240108
rect 91928 237380 91980 237386
rect 91928 237322 91980 237328
rect 92584 219434 92612 240108
rect 93228 231130 93256 240108
rect 93216 231124 93268 231130
rect 93216 231066 93268 231072
rect 89824 219406 90680 219434
rect 92492 219406 92612 219434
rect 89824 200938 89852 219406
rect 92492 205018 92520 219406
rect 93872 213314 93900 240108
rect 94516 223038 94544 240108
rect 95160 238202 95188 240108
rect 95804 238814 95832 240108
rect 95792 238808 95844 238814
rect 95792 238750 95844 238756
rect 95148 238196 95200 238202
rect 95148 238138 95200 238144
rect 96448 233918 96476 240108
rect 95240 233912 95292 233918
rect 95240 233854 95292 233860
rect 96436 233912 96488 233918
rect 96436 233854 96488 233860
rect 94504 223032 94556 223038
rect 94504 222974 94556 222980
rect 93860 213308 93912 213314
rect 93860 213250 93912 213256
rect 92480 205012 92532 205018
rect 92480 204954 92532 204960
rect 89812 200932 89864 200938
rect 89812 200874 89864 200880
rect 89720 192568 89772 192574
rect 89720 192510 89772 192516
rect 88432 188352 88484 188358
rect 88432 188294 88484 188300
rect 95252 185706 95280 233854
rect 97092 219434 97120 240108
rect 97736 236706 97764 240108
rect 98380 238542 98408 240108
rect 99024 238610 99052 240108
rect 99012 238604 99064 238610
rect 99012 238546 99064 238552
rect 98368 238536 98420 238542
rect 98368 238478 98420 238484
rect 97724 236700 97776 236706
rect 97724 236642 97776 236648
rect 99380 233912 99432 233918
rect 99380 233854 99432 233860
rect 96632 219406 97120 219434
rect 96632 198082 96660 219406
rect 99392 199578 99420 233854
rect 99668 227050 99696 240108
rect 100312 233918 100340 240108
rect 100300 233912 100352 233918
rect 100300 233854 100352 233860
rect 100760 231056 100812 231062
rect 100760 230998 100812 231004
rect 99656 227044 99708 227050
rect 99656 226986 99708 226992
rect 100772 203658 100800 230998
rect 100956 219434 100984 240108
rect 101600 231062 101628 240108
rect 102244 238754 102272 240108
rect 102152 238726 102272 238754
rect 101588 231056 101640 231062
rect 101588 230998 101640 231004
rect 100864 219406 100984 219434
rect 100864 203726 100892 219406
rect 100852 203720 100904 203726
rect 100852 203662 100904 203668
rect 100760 203652 100812 203658
rect 100760 203594 100812 203600
rect 99380 199572 99432 199578
rect 99380 199514 99432 199520
rect 96620 198076 96672 198082
rect 96620 198018 96672 198024
rect 100668 187808 100720 187814
rect 100668 187750 100720 187756
rect 95240 185700 95292 185706
rect 95240 185642 95292 185648
rect 80060 185632 80112 185638
rect 80060 185574 80112 185580
rect 73160 182980 73212 182986
rect 73160 182922 73212 182928
rect 71780 180192 71832 180198
rect 71780 180134 71832 180140
rect 97354 179480 97410 179489
rect 97354 179415 97410 179424
rect 70400 178696 70452 178702
rect 70400 178638 70452 178644
rect 97368 176905 97396 179415
rect 99104 178152 99156 178158
rect 99104 178094 99156 178100
rect 97354 176896 97410 176905
rect 97354 176831 97410 176840
rect 99116 176769 99144 178094
rect 100680 177585 100708 187750
rect 102152 184210 102180 238726
rect 102888 221474 102916 240108
rect 103532 237318 103560 240108
rect 103520 237312 103572 237318
rect 103520 237254 103572 237260
rect 103612 233912 103664 233918
rect 103612 233854 103664 233860
rect 102876 221468 102928 221474
rect 102876 221410 102928 221416
rect 103624 204921 103652 233854
rect 104176 219434 104204 240108
rect 104820 233918 104848 240108
rect 105464 238134 105492 240108
rect 105452 238128 105504 238134
rect 105452 238070 105504 238076
rect 106108 233918 106136 240108
rect 106752 235958 106780 240108
rect 107396 238754 107424 240108
rect 106844 238726 107424 238754
rect 106740 235952 106792 235958
rect 106740 235894 106792 235900
rect 104808 233912 104860 233918
rect 104808 233854 104860 233860
rect 104900 233912 104952 233918
rect 104900 233854 104952 233860
rect 106096 233912 106148 233918
rect 106096 233854 106148 233860
rect 103716 219406 104204 219434
rect 103610 204912 103666 204921
rect 103610 204847 103666 204856
rect 103716 200802 103744 219406
rect 104912 202162 104940 233854
rect 106844 229090 106872 238726
rect 106924 238196 106976 238202
rect 106924 238138 106976 238144
rect 106832 229084 106884 229090
rect 106832 229026 106884 229032
rect 106936 213246 106964 238138
rect 108040 235346 108068 240108
rect 108028 235340 108080 235346
rect 108028 235282 108080 235288
rect 108684 222970 108712 240108
rect 108672 222964 108724 222970
rect 108672 222906 108724 222912
rect 109972 219434 110000 240108
rect 110420 233912 110472 233918
rect 110420 233854 110472 233860
rect 109052 219406 110000 219434
rect 106924 213240 106976 213246
rect 106924 213182 106976 213188
rect 104900 202156 104952 202162
rect 104900 202098 104952 202104
rect 103704 200796 103756 200802
rect 103704 200738 103756 200744
rect 109052 189786 109080 219406
rect 110432 214577 110460 233854
rect 110616 223106 110644 240108
rect 111260 233918 111288 240108
rect 111248 233912 111300 233918
rect 111248 233854 111300 233860
rect 110604 223100 110656 223106
rect 110604 223042 110656 223048
rect 111904 219434 111932 240108
rect 112548 235890 112576 240108
rect 113192 238754 113220 240108
rect 113192 238726 113404 238754
rect 113836 238746 113864 240108
rect 112536 235884 112588 235890
rect 112536 235826 112588 235832
rect 111812 219406 111932 219434
rect 110418 214568 110474 214577
rect 110418 214503 110474 214512
rect 111812 196722 111840 219406
rect 111800 196716 111852 196722
rect 111800 196658 111852 196664
rect 109040 189780 109092 189786
rect 109040 189722 109092 189728
rect 106188 189100 106240 189106
rect 106188 189042 106240 189048
rect 102140 184204 102192 184210
rect 102140 184146 102192 184152
rect 106200 177585 106228 189042
rect 107568 187740 107620 187746
rect 107568 187682 107620 187688
rect 107580 177585 107608 187682
rect 112168 181008 112220 181014
rect 112168 180950 112220 180956
rect 110696 180940 110748 180946
rect 110696 180882 110748 180888
rect 110052 179444 110104 179450
rect 110052 179386 110104 179392
rect 100666 177576 100722 177585
rect 100666 177511 100722 177520
rect 106186 177576 106242 177585
rect 106186 177511 106242 177520
rect 107566 177576 107622 177585
rect 107566 177511 107622 177520
rect 108120 176928 108172 176934
rect 108120 176870 108172 176876
rect 102048 176860 102100 176866
rect 102048 176802 102100 176808
rect 102060 176769 102088 176802
rect 108132 176769 108160 176870
rect 110064 176769 110092 179386
rect 110708 177585 110736 180882
rect 112180 177585 112208 180950
rect 113376 180266 113404 238726
rect 113824 238740 113876 238746
rect 113824 238682 113876 238688
rect 114480 237250 114508 240108
rect 115124 238814 115152 240108
rect 115112 238808 115164 238814
rect 115112 238750 115164 238756
rect 114468 237244 114520 237250
rect 114468 237186 114520 237192
rect 115768 232218 115796 240108
rect 114560 232212 114612 232218
rect 114560 232154 114612 232160
rect 115756 232212 115808 232218
rect 115756 232154 115808 232160
rect 114572 203590 114600 232154
rect 116412 219434 116440 240108
rect 117056 238882 117084 240108
rect 117044 238876 117096 238882
rect 117044 238818 117096 238824
rect 117700 233918 117728 240108
rect 118344 238649 118372 240108
rect 118988 239970 119016 240108
rect 119646 240094 119936 240110
rect 118976 239964 119028 239970
rect 118976 239906 119028 239912
rect 118330 238640 118386 238649
rect 118330 238575 118386 238584
rect 117688 233912 117740 233918
rect 117688 233854 117740 233860
rect 115952 219406 116440 219434
rect 114560 203584 114612 203590
rect 114560 203526 114612 203532
rect 115952 202298 115980 219406
rect 120184 202842 120212 250951
rect 120736 246401 120764 293927
rect 121472 267458 121500 322186
rect 121552 312588 121604 312594
rect 121552 312530 121604 312536
rect 121564 285818 121592 312530
rect 121644 309800 121696 309806
rect 121644 309742 121696 309748
rect 121656 291825 121684 309742
rect 121642 291816 121698 291825
rect 121642 291751 121698 291760
rect 121734 291136 121790 291145
rect 121734 291071 121790 291080
rect 121642 290456 121698 290465
rect 121642 290391 121698 290400
rect 121656 289950 121684 290391
rect 121644 289944 121696 289950
rect 121644 289886 121696 289892
rect 121748 289882 121776 291071
rect 121736 289876 121788 289882
rect 121736 289818 121788 289824
rect 121644 289808 121696 289814
rect 121642 289776 121644 289785
rect 121696 289776 121698 289785
rect 121642 289711 121698 289720
rect 121642 289096 121698 289105
rect 121642 289031 121698 289040
rect 121656 288454 121684 289031
rect 121644 288448 121696 288454
rect 121644 288390 121696 288396
rect 121826 288416 121882 288425
rect 121826 288351 121882 288360
rect 121642 287056 121698 287065
rect 121642 286991 121644 287000
rect 121696 286991 121698 287000
rect 121644 286962 121696 286968
rect 121840 286346 121868 288351
rect 122194 287736 122250 287745
rect 122194 287671 122250 287680
rect 121828 286340 121880 286346
rect 121828 286282 121880 286288
rect 121564 285790 121776 285818
rect 121552 285728 121604 285734
rect 121550 285696 121552 285705
rect 121604 285696 121606 285705
rect 121550 285631 121606 285640
rect 121644 285660 121696 285666
rect 121644 285602 121696 285608
rect 121550 285016 121606 285025
rect 121550 284951 121606 284960
rect 121564 284374 121592 284951
rect 121552 284368 121604 284374
rect 121656 284345 121684 285602
rect 121552 284310 121604 284316
rect 121642 284336 121698 284345
rect 121642 284271 121698 284280
rect 121552 284164 121604 284170
rect 121552 284106 121604 284112
rect 121564 283665 121592 284106
rect 121550 283656 121606 283665
rect 121550 283591 121606 283600
rect 121550 282976 121606 282985
rect 121550 282911 121552 282920
rect 121604 282911 121606 282920
rect 121552 282882 121604 282888
rect 121550 282296 121606 282305
rect 121550 282231 121606 282240
rect 121564 281586 121592 282231
rect 121552 281580 121604 281586
rect 121552 281522 121604 281528
rect 121642 280936 121698 280945
rect 121642 280871 121698 280880
rect 121552 280288 121604 280294
rect 121550 280256 121552 280265
rect 121604 280256 121606 280265
rect 121656 280226 121684 280871
rect 121550 280191 121606 280200
rect 121644 280220 121696 280226
rect 121644 280162 121696 280168
rect 121642 279576 121698 279585
rect 121642 279511 121698 279520
rect 121550 278896 121606 278905
rect 121550 278831 121552 278840
rect 121604 278831 121606 278840
rect 121552 278802 121604 278808
rect 121656 278798 121684 279511
rect 121644 278792 121696 278798
rect 121644 278734 121696 278740
rect 121642 278216 121698 278225
rect 121642 278151 121698 278160
rect 121550 277536 121606 277545
rect 121656 277506 121684 278151
rect 121550 277471 121606 277480
rect 121644 277500 121696 277506
rect 121564 277438 121592 277471
rect 121644 277442 121696 277448
rect 121552 277432 121604 277438
rect 121552 277374 121604 277380
rect 121748 277394 121776 285790
rect 122102 281616 122158 281625
rect 122102 281551 122158 281560
rect 121748 277366 121868 277394
rect 121642 276856 121698 276865
rect 121642 276791 121698 276800
rect 121550 276176 121606 276185
rect 121656 276146 121684 276791
rect 121550 276111 121606 276120
rect 121644 276140 121696 276146
rect 121564 276078 121592 276111
rect 121644 276082 121696 276088
rect 121552 276072 121604 276078
rect 121552 276014 121604 276020
rect 121734 275496 121790 275505
rect 121734 275431 121790 275440
rect 121550 274816 121606 274825
rect 121550 274751 121606 274760
rect 121564 274718 121592 274751
rect 121552 274712 121604 274718
rect 121552 274654 121604 274660
rect 121644 274644 121696 274650
rect 121644 274586 121696 274592
rect 121656 274145 121684 274586
rect 121642 274136 121698 274145
rect 121642 274071 121698 274080
rect 121550 273456 121606 273465
rect 121550 273391 121606 273400
rect 121564 273290 121592 273391
rect 121552 273284 121604 273290
rect 121552 273226 121604 273232
rect 121644 273216 121696 273222
rect 121644 273158 121696 273164
rect 121656 272785 121684 273158
rect 121642 272776 121698 272785
rect 121642 272711 121698 272720
rect 121748 272542 121776 275431
rect 121736 272536 121788 272542
rect 121736 272478 121788 272484
rect 121550 271416 121606 271425
rect 121550 271351 121606 271360
rect 121564 270570 121592 271351
rect 121552 270564 121604 270570
rect 121552 270506 121604 270512
rect 121642 270056 121698 270065
rect 121642 269991 121698 270000
rect 121550 269376 121606 269385
rect 121550 269311 121606 269320
rect 121564 269142 121592 269311
rect 121656 269210 121684 269991
rect 121644 269204 121696 269210
rect 121644 269146 121696 269152
rect 121552 269136 121604 269142
rect 121552 269078 121604 269084
rect 121840 268705 121868 277366
rect 121826 268696 121882 268705
rect 121826 268631 121882 268640
rect 121550 268016 121606 268025
rect 121550 267951 121606 267960
rect 121564 267782 121592 267951
rect 121552 267776 121604 267782
rect 121552 267718 121604 267724
rect 121472 267430 121684 267458
rect 121458 267336 121514 267345
rect 121458 267271 121514 267280
rect 121472 266422 121500 267271
rect 121460 266416 121512 266422
rect 121460 266358 121512 266364
rect 121550 265976 121606 265985
rect 121550 265911 121606 265920
rect 121458 265296 121514 265305
rect 121458 265231 121514 265240
rect 121472 265062 121500 265231
rect 121460 265056 121512 265062
rect 121460 264998 121512 265004
rect 121564 264994 121592 265911
rect 121552 264988 121604 264994
rect 121552 264930 121604 264936
rect 121460 264920 121512 264926
rect 121460 264862 121512 264868
rect 121472 264625 121500 264862
rect 121458 264616 121514 264625
rect 121458 264551 121514 264560
rect 121458 263936 121514 263945
rect 121458 263871 121514 263880
rect 121472 262886 121500 263871
rect 121656 263265 121684 267430
rect 122116 267034 122144 281551
rect 122208 275330 122236 287671
rect 122196 275324 122248 275330
rect 122196 275266 122248 275272
rect 122104 267028 122156 267034
rect 122104 266970 122156 266976
rect 122194 266656 122250 266665
rect 122194 266591 122250 266600
rect 121642 263256 121698 263265
rect 121642 263191 121698 263200
rect 121460 262880 121512 262886
rect 121460 262822 121512 262828
rect 121458 262576 121514 262585
rect 121458 262511 121514 262520
rect 121472 262274 121500 262511
rect 121460 262268 121512 262274
rect 121460 262210 121512 262216
rect 121458 261896 121514 261905
rect 121458 261831 121514 261840
rect 121472 260914 121500 261831
rect 121460 260908 121512 260914
rect 121460 260850 121512 260856
rect 121458 259856 121514 259865
rect 121458 259791 121514 259800
rect 121472 259486 121500 259791
rect 121460 259480 121512 259486
rect 121460 259422 121512 259428
rect 121460 259344 121512 259350
rect 121460 259286 121512 259292
rect 121472 258505 121500 259286
rect 122102 259176 122158 259185
rect 122102 259111 122158 259120
rect 121458 258496 121514 258505
rect 121458 258431 121514 258440
rect 121642 257816 121698 257825
rect 121642 257751 121698 257760
rect 121460 257168 121512 257174
rect 121458 257136 121460 257145
rect 121512 257136 121514 257145
rect 121458 257071 121514 257080
rect 121656 256766 121684 257751
rect 121644 256760 121696 256766
rect 121644 256702 121696 256708
rect 121552 256692 121604 256698
rect 121552 256634 121604 256640
rect 121460 256488 121512 256494
rect 121458 256456 121460 256465
rect 121512 256456 121514 256465
rect 121458 256391 121514 256400
rect 121564 255785 121592 256634
rect 121550 255776 121606 255785
rect 121550 255711 121606 255720
rect 121550 255096 121606 255105
rect 121550 255031 121606 255040
rect 121458 254416 121514 254425
rect 121458 254351 121514 254360
rect 121472 254046 121500 254351
rect 121460 254040 121512 254046
rect 121460 253982 121512 253988
rect 121564 253978 121592 255031
rect 121552 253972 121604 253978
rect 121552 253914 121604 253920
rect 121550 253736 121606 253745
rect 121550 253671 121606 253680
rect 121458 253056 121514 253065
rect 121458 252991 121514 253000
rect 121472 252618 121500 252991
rect 121564 252686 121592 253671
rect 121644 253224 121696 253230
rect 121644 253166 121696 253172
rect 121552 252680 121604 252686
rect 121552 252622 121604 252628
rect 121460 252612 121512 252618
rect 121460 252554 121512 252560
rect 121656 252385 121684 253166
rect 121642 252376 121698 252385
rect 121642 252311 121698 252320
rect 121458 251696 121514 251705
rect 121458 251631 121514 251640
rect 121472 251258 121500 251631
rect 121460 251252 121512 251258
rect 121460 251194 121512 251200
rect 122116 250510 122144 259111
rect 122208 257378 122236 266591
rect 122196 257372 122248 257378
rect 122196 257314 122248 257320
rect 123496 256494 123524 430578
rect 123576 324352 123628 324358
rect 123576 324294 123628 324300
rect 123588 257174 123616 324294
rect 123668 305652 123720 305658
rect 123668 305594 123720 305600
rect 123680 287026 123708 305594
rect 123668 287020 123720 287026
rect 123668 286962 123720 286968
rect 124876 284170 124904 702578
rect 126244 630692 126296 630698
rect 126244 630634 126296 630640
rect 124956 378208 125008 378214
rect 124956 378150 125008 378156
rect 124968 289814 124996 378150
rect 125140 313948 125192 313954
rect 125140 313890 125192 313896
rect 125046 292768 125102 292777
rect 125046 292703 125102 292712
rect 124956 289808 125008 289814
rect 124956 289750 125008 289756
rect 124864 284164 124916 284170
rect 124864 284106 124916 284112
rect 123576 257168 123628 257174
rect 123576 257110 123628 257116
rect 123484 256488 123536 256494
rect 123484 256430 123536 256436
rect 122104 250504 122156 250510
rect 122104 250446 122156 250452
rect 121550 250336 121606 250345
rect 121550 250271 121606 250280
rect 121564 249830 121592 250271
rect 121552 249824 121604 249830
rect 121552 249766 121604 249772
rect 121460 249756 121512 249762
rect 121460 249698 121512 249704
rect 121472 249665 121500 249698
rect 121458 249656 121514 249665
rect 121458 249591 121514 249600
rect 121458 248976 121514 248985
rect 121458 248911 121514 248920
rect 121472 248470 121500 248911
rect 121460 248464 121512 248470
rect 121460 248406 121512 248412
rect 121458 248296 121514 248305
rect 121458 248231 121514 248240
rect 121472 247110 121500 248231
rect 121460 247104 121512 247110
rect 121460 247046 121512 247052
rect 121550 246936 121606 246945
rect 121550 246871 121606 246880
rect 120722 246392 120778 246401
rect 120722 246327 120778 246336
rect 121564 245682 121592 246871
rect 121642 246256 121698 246265
rect 121642 246191 121698 246200
rect 121552 245676 121604 245682
rect 121552 245618 121604 245624
rect 121460 245608 121512 245614
rect 121460 245550 121512 245556
rect 121550 245576 121606 245585
rect 121472 244905 121500 245550
rect 121550 245511 121606 245520
rect 121458 244896 121514 244905
rect 121458 244831 121514 244840
rect 121564 244322 121592 245511
rect 121552 244316 121604 244322
rect 121552 244258 121604 244264
rect 121550 244216 121606 244225
rect 121550 244151 121606 244160
rect 121460 243772 121512 243778
rect 121460 243714 121512 243720
rect 121472 243545 121500 243714
rect 121458 243536 121514 243545
rect 121458 243471 121514 243480
rect 121564 242962 121592 244151
rect 121656 243545 121684 246191
rect 121642 243536 121698 243545
rect 121642 243471 121698 243480
rect 121552 242956 121604 242962
rect 121552 242898 121604 242904
rect 121460 242888 121512 242894
rect 121458 242856 121460 242865
rect 121512 242856 121514 242865
rect 121458 242791 121514 242800
rect 121552 242820 121604 242826
rect 121552 242762 121604 242768
rect 121564 242185 121592 242762
rect 121550 242176 121606 242185
rect 121550 242111 121606 242120
rect 121458 241496 121514 241505
rect 121458 241431 121514 241440
rect 121472 235278 121500 241431
rect 122102 240816 122158 240825
rect 122102 240751 122158 240760
rect 121552 240236 121604 240242
rect 121552 240178 121604 240184
rect 121564 240145 121592 240178
rect 121550 240136 121606 240145
rect 121550 240071 121606 240080
rect 121460 235272 121512 235278
rect 121460 235214 121512 235220
rect 120172 202836 120224 202842
rect 120172 202778 120224 202784
rect 115940 202292 115992 202298
rect 115940 202234 115992 202240
rect 122116 191214 122144 240751
rect 125060 206990 125088 292703
rect 125152 243778 125180 313890
rect 125140 243772 125192 243778
rect 125140 243714 125192 243720
rect 126256 238882 126284 630634
rect 126336 311908 126388 311914
rect 126336 311850 126388 311856
rect 126348 274650 126376 311850
rect 126428 295656 126480 295662
rect 126428 295598 126480 295604
rect 126336 274644 126388 274650
rect 126336 274586 126388 274592
rect 126440 259418 126468 295598
rect 126978 293176 127034 293185
rect 126978 293111 127034 293120
rect 126992 273222 127020 293111
rect 126980 273216 127032 273222
rect 126980 273158 127032 273164
rect 126428 259412 126480 259418
rect 126428 259354 126480 259360
rect 129016 245614 129044 702850
rect 134524 702568 134576 702574
rect 134524 702510 134576 702516
rect 130384 616888 130436 616894
rect 130384 616830 130436 616836
rect 129096 484424 129148 484430
rect 129096 484366 129148 484372
rect 129108 264926 129136 484366
rect 129096 264920 129148 264926
rect 129096 264862 129148 264868
rect 130396 256698 130424 616830
rect 130476 364404 130528 364410
rect 130476 364346 130528 364352
rect 130384 256692 130436 256698
rect 130384 256634 130436 256640
rect 129004 245608 129056 245614
rect 129004 245550 129056 245556
rect 126244 238876 126296 238882
rect 126244 238818 126296 238824
rect 130488 238678 130516 364346
rect 134536 242826 134564 702510
rect 135904 700324 135956 700330
rect 135904 700266 135956 700272
rect 134524 242820 134576 242826
rect 134524 242762 134576 242768
rect 130476 238672 130528 238678
rect 130476 238614 130528 238620
rect 135916 238610 135944 700266
rect 137848 697610 137876 703520
rect 154132 702434 154160 703520
rect 153212 702406 154160 702434
rect 149704 700460 149756 700466
rect 149704 700402 149756 700408
rect 137836 697604 137888 697610
rect 137836 697546 137888 697552
rect 144184 683188 144236 683194
rect 144184 683130 144236 683136
rect 142804 576904 142856 576910
rect 142804 576846 142856 576852
rect 140044 524476 140096 524482
rect 140044 524418 140096 524424
rect 138664 470620 138716 470626
rect 138664 470562 138716 470568
rect 138676 285666 138704 470562
rect 138664 285660 138716 285666
rect 138664 285602 138716 285608
rect 140056 249762 140084 524418
rect 142816 251870 142844 576846
rect 144196 253230 144224 683130
rect 148324 670744 148376 670750
rect 148324 670686 148376 670692
rect 148336 319462 148364 670686
rect 148324 319456 148376 319462
rect 148324 319398 148376 319404
rect 148324 291372 148376 291378
rect 148324 291314 148376 291320
rect 144184 253224 144236 253230
rect 144184 253166 144236 253172
rect 142804 251864 142856 251870
rect 142804 251806 142856 251812
rect 140044 249756 140096 249762
rect 140044 249698 140096 249704
rect 135904 238604 135956 238610
rect 135904 238546 135956 238552
rect 125048 206984 125100 206990
rect 125048 206926 125100 206932
rect 148336 199510 148364 291314
rect 149716 259350 149744 700402
rect 153212 311166 153240 702406
rect 170324 700398 170352 703520
rect 202800 703118 202828 703520
rect 201500 703112 201552 703118
rect 201500 703054 201552 703060
rect 202788 703112 202840 703118
rect 202788 703054 202840 703060
rect 170312 700392 170364 700398
rect 170312 700334 170364 700340
rect 153200 311160 153252 311166
rect 153200 311102 153252 311108
rect 201512 305658 201540 703054
rect 218992 699718 219020 703520
rect 235184 700466 235212 703520
rect 235172 700460 235224 700466
rect 235172 700402 235224 700408
rect 267660 699718 267688 703520
rect 283852 702434 283880 703520
rect 282932 702406 283880 702434
rect 269764 700392 269816 700398
rect 269764 700334 269816 700340
rect 214564 699712 214616 699718
rect 214564 699654 214616 699660
rect 218980 699712 219032 699718
rect 218980 699654 219032 699660
rect 264244 699712 264296 699718
rect 264244 699654 264296 699660
rect 267648 699712 267700 699718
rect 267648 699654 267700 699660
rect 201500 305652 201552 305658
rect 201500 305594 201552 305600
rect 185584 303816 185636 303822
rect 185584 303758 185636 303764
rect 152464 300960 152516 300966
rect 152464 300902 152516 300908
rect 149704 259344 149756 259350
rect 149704 259286 149756 259292
rect 148324 199504 148376 199510
rect 148324 199446 148376 199452
rect 152476 196625 152504 300902
rect 184204 299736 184256 299742
rect 184204 299678 184256 299684
rect 166264 298512 166316 298518
rect 166264 298454 166316 298460
rect 160744 297084 160796 297090
rect 160744 297026 160796 297032
rect 157984 295724 158036 295730
rect 157984 295666 158036 295672
rect 152462 196616 152518 196625
rect 152462 196551 152518 196560
rect 122104 191208 122156 191214
rect 122104 191150 122156 191156
rect 157996 189786 158024 295666
rect 160756 209166 160784 297026
rect 166276 249082 166304 298454
rect 174544 298444 174596 298450
rect 174544 298386 174596 298392
rect 170404 294364 170456 294370
rect 170404 294306 170456 294312
rect 166264 249076 166316 249082
rect 166264 249018 166316 249024
rect 166262 236600 166318 236609
rect 166262 236535 166318 236544
rect 160744 209160 160796 209166
rect 160744 209102 160796 209108
rect 157984 189780 158036 189786
rect 157984 189722 158036 189728
rect 126796 186448 126848 186454
rect 126796 186390 126848 186396
rect 117228 186380 117280 186386
rect 117228 186322 117280 186328
rect 114376 182232 114428 182238
rect 114376 182174 114428 182180
rect 113364 180260 113416 180266
rect 113364 180202 113416 180208
rect 114388 177585 114416 182174
rect 115848 178220 115900 178226
rect 115848 178162 115900 178168
rect 110694 177576 110750 177585
rect 110694 177511 110750 177520
rect 112166 177576 112222 177585
rect 112166 177511 112222 177520
rect 114374 177576 114430 177585
rect 114374 177511 114430 177520
rect 115860 176769 115888 178162
rect 117240 177585 117268 186322
rect 118608 184952 118660 184958
rect 118608 184894 118660 184900
rect 118620 177585 118648 184894
rect 124128 183592 124180 183598
rect 124128 183534 124180 183540
rect 121184 179512 121236 179518
rect 121184 179454 121236 179460
rect 117226 177576 117282 177585
rect 117226 177511 117282 177520
rect 118606 177576 118662 177585
rect 118606 177511 118662 177520
rect 121196 177177 121224 179454
rect 124140 177585 124168 183534
rect 125048 180872 125100 180878
rect 125048 180814 125100 180820
rect 125060 177585 125088 180814
rect 126808 177585 126836 186390
rect 166276 183054 166304 236535
rect 167828 183592 167880 183598
rect 167828 183534 167880 183540
rect 166264 183048 166316 183054
rect 166264 182990 166316 182996
rect 128176 182300 128228 182306
rect 128176 182242 128228 182248
rect 166448 182300 166500 182306
rect 166448 182242 166500 182248
rect 124126 177576 124182 177585
rect 124126 177511 124182 177520
rect 125046 177576 125102 177585
rect 125046 177511 125102 177520
rect 126794 177576 126850 177585
rect 126794 177511 126850 177520
rect 121182 177168 121238 177177
rect 121182 177103 121238 177112
rect 128188 176769 128216 182242
rect 133144 179580 133196 179586
rect 133144 179522 133196 179528
rect 165068 179580 165120 179586
rect 165068 179522 165120 179528
rect 129464 178084 129516 178090
rect 129464 178026 129516 178032
rect 129476 176769 129504 178026
rect 133156 177177 133184 179522
rect 148232 178356 148284 178362
rect 148232 178298 148284 178304
rect 134708 178288 134760 178294
rect 134708 178230 134760 178236
rect 133142 177168 133198 177177
rect 133142 177103 133198 177112
rect 132040 176996 132092 177002
rect 132040 176938 132092 176944
rect 132052 176769 132080 176938
rect 134720 176769 134748 178230
rect 135720 176792 135772 176798
rect 99102 176760 99158 176769
rect 99102 176695 99158 176704
rect 102046 176760 102102 176769
rect 102046 176695 102102 176704
rect 108118 176760 108174 176769
rect 108118 176695 108174 176704
rect 110050 176760 110106 176769
rect 110050 176695 110106 176704
rect 115846 176760 115902 176769
rect 115846 176695 115902 176704
rect 127070 176760 127126 176769
rect 127070 176695 127072 176704
rect 127124 176695 127126 176704
rect 128174 176760 128230 176769
rect 128174 176695 128230 176704
rect 129462 176760 129518 176769
rect 129462 176695 129518 176704
rect 132038 176760 132094 176769
rect 132038 176695 132094 176704
rect 134706 176760 134762 176769
rect 134706 176695 134762 176704
rect 135718 176760 135720 176769
rect 148244 176769 148272 178298
rect 135772 176760 135774 176769
rect 135718 176695 135774 176704
rect 148230 176760 148286 176769
rect 148230 176695 148286 176704
rect 127072 176666 127124 176672
rect 121920 176248 121972 176254
rect 121920 176190 121972 176196
rect 119436 176180 119488 176186
rect 119436 176122 119488 176128
rect 100760 175976 100812 175982
rect 100760 175918 100812 175924
rect 100772 175409 100800 175918
rect 100758 175400 100814 175409
rect 100758 175335 100814 175344
rect 119448 175001 119476 176122
rect 121932 175409 121960 176190
rect 158904 176112 158956 176118
rect 158904 176054 158956 176060
rect 130752 176044 130804 176050
rect 130752 175986 130804 175992
rect 130764 175545 130792 175986
rect 158916 175545 158944 176054
rect 130750 175536 130806 175545
rect 130750 175471 130806 175480
rect 158902 175536 158958 175545
rect 158902 175471 158958 175480
rect 121918 175400 121974 175409
rect 121918 175335 121974 175344
rect 165080 175166 165108 179522
rect 166356 179512 166408 179518
rect 166356 179454 166408 179460
rect 165436 178288 165488 178294
rect 165436 178230 165488 178236
rect 165448 175234 165476 178230
rect 166264 178220 166316 178226
rect 166264 178162 166316 178168
rect 165528 176996 165580 177002
rect 165528 176938 165580 176944
rect 165436 175228 165488 175234
rect 165436 175170 165488 175176
rect 165068 175160 165120 175166
rect 165068 175102 165120 175108
rect 119434 174992 119490 175001
rect 119434 174927 119490 174936
rect 67362 129296 67418 129305
rect 67362 129231 67418 129240
rect 64970 126304 65026 126313
rect 64970 126239 65026 126248
rect 64984 125633 65012 126239
rect 64970 125624 65026 125633
rect 64970 125559 65026 125568
rect 66166 125216 66222 125225
rect 66166 125151 66222 125160
rect 66074 123584 66130 123593
rect 66074 123519 66130 123528
rect 66088 122874 66116 123519
rect 66076 122868 66128 122874
rect 66076 122810 66128 122816
rect 66074 102368 66130 102377
rect 66074 102303 66130 102312
rect 66088 85474 66116 102303
rect 66180 91089 66208 125151
rect 67270 100736 67326 100745
rect 67270 100671 67326 100680
rect 66166 91080 66222 91089
rect 66166 91015 66222 91024
rect 67284 88330 67312 100671
rect 67376 93838 67404 129231
rect 67638 128072 67694 128081
rect 67638 128007 67694 128016
rect 67454 122632 67510 122641
rect 67454 122567 67510 122576
rect 67364 93832 67416 93838
rect 67364 93774 67416 93780
rect 67272 88324 67324 88330
rect 67272 88266 67324 88272
rect 66076 85468 66128 85474
rect 66076 85410 66128 85416
rect 67468 82822 67496 122567
rect 67546 120864 67602 120873
rect 67546 120799 67602 120808
rect 67456 82816 67508 82822
rect 67456 82758 67508 82764
rect 67560 80034 67588 120799
rect 67652 93809 67680 128007
rect 165540 173874 165568 176938
rect 165528 173868 165580 173874
rect 165528 173810 165580 173816
rect 166276 165578 166304 178162
rect 166368 168366 166396 179454
rect 166460 172514 166488 182242
rect 167736 181008 167788 181014
rect 167736 180950 167788 180956
rect 166540 176180 166592 176186
rect 166540 176122 166592 176128
rect 166448 172508 166500 172514
rect 166448 172450 166500 172456
rect 166356 168360 166408 168366
rect 166356 168302 166408 168308
rect 166552 167006 166580 176122
rect 167642 171592 167698 171601
rect 167642 171527 167698 171536
rect 166540 167000 166592 167006
rect 166540 166942 166592 166948
rect 166264 165572 166316 165578
rect 166264 165514 166316 165520
rect 167656 151094 167684 171527
rect 167748 164218 167776 180950
rect 167840 169726 167868 183534
rect 169208 182232 169260 182238
rect 169208 182174 169260 182180
rect 169116 180940 169168 180946
rect 169116 180882 169168 180888
rect 169024 178356 169076 178362
rect 169024 178298 169076 178304
rect 167920 176248 167972 176254
rect 167920 176190 167972 176196
rect 167828 169720 167880 169726
rect 167828 169662 167880 169668
rect 167932 168298 167960 176190
rect 167920 168292 167972 168298
rect 167920 168234 167972 168240
rect 167736 164212 167788 164218
rect 167736 164154 167788 164160
rect 167644 151088 167696 151094
rect 167644 151030 167696 151036
rect 169036 150414 169064 178298
rect 169128 162858 169156 180882
rect 169220 165510 169248 182174
rect 170416 177342 170444 294306
rect 171784 187808 171836 187814
rect 171784 187750 171836 187756
rect 170588 184952 170640 184958
rect 170588 184894 170640 184900
rect 170496 178152 170548 178158
rect 170496 178094 170548 178100
rect 170404 177336 170456 177342
rect 170404 177278 170456 177284
rect 169208 165504 169260 165510
rect 169208 165446 169260 165452
rect 169116 162852 169168 162858
rect 169116 162794 169168 162800
rect 170508 155922 170536 178094
rect 170600 166938 170628 184894
rect 170680 176928 170732 176934
rect 170680 176870 170732 176876
rect 170588 166932 170640 166938
rect 170588 166874 170640 166880
rect 170692 161430 170720 176870
rect 170680 161424 170732 161430
rect 170680 161366 170732 161372
rect 171796 157350 171824 187750
rect 171968 186448 172020 186454
rect 171968 186390 172020 186396
rect 171876 176860 171928 176866
rect 171876 176802 171928 176808
rect 171888 160750 171916 176802
rect 171980 171086 172008 186390
rect 174556 181558 174584 298386
rect 178684 295588 178736 295594
rect 178684 295530 178736 295536
rect 175924 229900 175976 229906
rect 175924 229842 175976 229848
rect 174544 181552 174596 181558
rect 174544 181494 174596 181500
rect 171968 171080 172020 171086
rect 171968 171022 172020 171028
rect 171876 160744 171928 160750
rect 171876 160686 171928 160692
rect 171784 157344 171836 157350
rect 171784 157286 171836 157292
rect 170496 155916 170548 155922
rect 170496 155858 170548 155864
rect 169024 150408 169076 150414
rect 169024 150350 169076 150356
rect 170404 147688 170456 147694
rect 170404 147630 170456 147636
rect 169024 142180 169076 142186
rect 169024 142122 169076 142128
rect 166264 139460 166316 139466
rect 166264 139402 166316 139408
rect 164884 96688 164936 96694
rect 164884 96630 164936 96636
rect 105450 94752 105506 94761
rect 105450 94687 105506 94696
rect 117962 94752 118018 94761
rect 117962 94687 118018 94696
rect 119526 94752 119582 94761
rect 119526 94687 119582 94696
rect 129370 94752 129426 94761
rect 129370 94687 129426 94696
rect 134338 94752 134394 94761
rect 134338 94687 134394 94696
rect 105464 94042 105492 94687
rect 117976 94110 118004 94687
rect 117964 94104 118016 94110
rect 117964 94046 118016 94052
rect 105452 94036 105504 94042
rect 105452 93978 105504 93984
rect 119540 93906 119568 94687
rect 129384 93974 129412 94687
rect 134352 94178 134380 94687
rect 134340 94172 134392 94178
rect 134340 94114 134392 94120
rect 129372 93968 129424 93974
rect 129372 93910 129424 93916
rect 119528 93900 119580 93906
rect 119528 93842 119580 93848
rect 67638 93800 67694 93809
rect 67638 93735 67694 93744
rect 130750 93664 130806 93673
rect 130750 93599 130806 93608
rect 151726 93664 151782 93673
rect 151726 93599 151782 93608
rect 110694 93528 110750 93537
rect 110694 93463 110750 93472
rect 115846 93528 115902 93537
rect 115846 93463 115902 93472
rect 110326 93256 110382 93265
rect 110708 93226 110736 93463
rect 115860 93294 115888 93463
rect 130764 93362 130792 93599
rect 151740 93430 151768 93599
rect 151728 93424 151780 93430
rect 151728 93366 151780 93372
rect 130752 93356 130804 93362
rect 130752 93298 130804 93304
rect 115848 93288 115900 93294
rect 115848 93230 115900 93236
rect 128174 93256 128230 93265
rect 110326 93191 110382 93200
rect 110696 93220 110748 93226
rect 85670 92440 85726 92449
rect 85670 92375 85726 92384
rect 91650 92440 91706 92449
rect 91650 92375 91706 92384
rect 107750 92440 107806 92449
rect 107750 92375 107806 92384
rect 85684 92342 85712 92375
rect 85672 92336 85724 92342
rect 85672 92278 85724 92284
rect 89350 91760 89406 91769
rect 89350 91695 89406 91704
rect 90546 91760 90602 91769
rect 90546 91695 90602 91704
rect 75366 91216 75422 91225
rect 75366 91151 75422 91160
rect 85486 91216 85542 91225
rect 85486 91151 85542 91160
rect 86866 91216 86922 91225
rect 86866 91151 86922 91160
rect 88062 91216 88118 91225
rect 88062 91151 88118 91160
rect 75380 86970 75408 91151
rect 75368 86964 75420 86970
rect 75368 86906 75420 86912
rect 67548 80028 67600 80034
rect 67548 79970 67600 79976
rect 85500 77246 85528 91151
rect 86880 81258 86908 91151
rect 88076 86902 88104 91151
rect 89364 89554 89392 91695
rect 90560 89690 90588 91695
rect 91664 91118 91692 92375
rect 99746 91760 99802 91769
rect 99746 91695 99802 91704
rect 99286 91488 99342 91497
rect 99286 91423 99342 91432
rect 95054 91352 95110 91361
rect 95054 91287 95110 91296
rect 97814 91352 97870 91361
rect 97814 91287 97870 91296
rect 99102 91352 99158 91361
rect 99102 91287 99158 91296
rect 93766 91216 93822 91225
rect 93766 91151 93822 91160
rect 91652 91112 91704 91118
rect 91652 91054 91704 91060
rect 90548 89684 90600 89690
rect 90548 89626 90600 89632
rect 89352 89548 89404 89554
rect 89352 89490 89404 89496
rect 88064 86896 88116 86902
rect 88064 86838 88116 86844
rect 86868 81252 86920 81258
rect 86868 81194 86920 81200
rect 93780 81190 93808 91151
rect 93768 81184 93820 81190
rect 93768 81126 93820 81132
rect 95068 79830 95096 91287
rect 95146 91216 95202 91225
rect 95146 91151 95202 91160
rect 96526 91216 96582 91225
rect 96526 91151 96582 91160
rect 95056 79824 95108 79830
rect 95056 79766 95108 79772
rect 85488 77240 85540 77246
rect 85488 77182 85540 77188
rect 77300 76628 77352 76634
rect 77300 76570 77352 76576
rect 68284 71052 68336 71058
rect 68284 70994 68336 71000
rect 66260 69692 66312 69698
rect 66260 69634 66312 69640
rect 64880 17332 64932 17338
rect 64880 17274 64932 17280
rect 64892 16574 64920 17274
rect 66272 16574 66300 69634
rect 64892 16546 65104 16574
rect 66272 16546 66760 16574
rect 64788 8288 64840 8294
rect 64788 8230 64840 8236
rect 61998 354 62110 480
rect 61580 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66732 480 66760 16546
rect 68296 3602 68324 70994
rect 71780 66972 71832 66978
rect 71780 66914 71832 66920
rect 69020 35284 69072 35290
rect 69020 35226 69072 35232
rect 68284 3596 68336 3602
rect 68284 3538 68336 3544
rect 69032 3534 69060 35226
rect 69112 18692 69164 18698
rect 69112 18634 69164 18640
rect 67916 3528 67968 3534
rect 67916 3470 67968 3476
rect 69020 3528 69072 3534
rect 69020 3470 69072 3476
rect 67928 480 67956 3470
rect 69124 480 69152 18634
rect 71792 16574 71820 66914
rect 73160 36644 73212 36650
rect 73160 36586 73212 36592
rect 73172 16574 73200 36586
rect 75920 22772 75972 22778
rect 75920 22714 75972 22720
rect 71792 16546 72648 16574
rect 73172 16546 73384 16574
rect 71504 7608 71556 7614
rect 71504 7550 71556 7556
rect 69940 3528 69992 3534
rect 69940 3470 69992 3476
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 69952 354 69980 3470
rect 71516 480 71544 7550
rect 72620 480 72648 16546
rect 70278 354 70390 480
rect 69952 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 16546
rect 75000 8968 75052 8974
rect 75000 8910 75052 8916
rect 75012 480 75040 8910
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 75932 354 75960 22714
rect 77312 3602 77340 76570
rect 89720 76560 89772 76566
rect 89720 76502 89772 76508
rect 82820 65544 82872 65550
rect 82820 65486 82872 65492
rect 80060 62892 80112 62898
rect 80060 62834 80112 62840
rect 77392 38004 77444 38010
rect 77392 37946 77444 37952
rect 77300 3596 77352 3602
rect 77300 3538 77352 3544
rect 77404 480 77432 37946
rect 78680 21480 78732 21486
rect 78680 21422 78732 21428
rect 78692 16574 78720 21422
rect 80072 16574 80100 62834
rect 81440 57248 81492 57254
rect 81440 57190 81492 57196
rect 81452 16574 81480 57190
rect 82832 16574 82860 65486
rect 84200 50448 84252 50454
rect 84200 50390 84252 50396
rect 78692 16546 79272 16574
rect 80072 16546 80928 16574
rect 81452 16546 81664 16574
rect 82832 16546 83320 16574
rect 78220 3596 78272 3602
rect 78220 3538 78272 3544
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78232 354 78260 3538
rect 78558 354 78670 480
rect 78232 326 78670 354
rect 79244 354 79272 16546
rect 80900 480 80928 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83292 480 83320 16546
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 50390
rect 86960 49088 87012 49094
rect 86960 49030 87012 49036
rect 85580 42152 85632 42158
rect 85580 42094 85632 42100
rect 85592 6914 85620 42094
rect 85672 31136 85724 31142
rect 85672 31078 85724 31084
rect 85684 16574 85712 31078
rect 86972 16574 87000 49030
rect 88340 47660 88392 47666
rect 88340 47602 88392 47608
rect 88352 16574 88380 47602
rect 89732 16574 89760 76502
rect 95160 75886 95188 91151
rect 96540 84153 96568 91151
rect 96526 84144 96582 84153
rect 96526 84079 96582 84088
rect 97828 81326 97856 91287
rect 97906 91216 97962 91225
rect 97906 91151 97962 91160
rect 97816 81320 97868 81326
rect 97816 81262 97868 81268
rect 97920 78674 97948 91151
rect 99116 82754 99144 91287
rect 99194 91216 99250 91225
rect 99194 91151 99250 91160
rect 99104 82748 99156 82754
rect 99104 82690 99156 82696
rect 97908 78668 97960 78674
rect 97908 78610 97960 78616
rect 99208 78470 99236 91151
rect 99300 78538 99328 91423
rect 99760 89622 99788 91695
rect 103150 91624 103206 91633
rect 103150 91559 103206 91568
rect 102046 91488 102102 91497
rect 102046 91423 102102 91432
rect 101862 91352 101918 91361
rect 101862 91287 101918 91296
rect 100574 91216 100630 91225
rect 100574 91151 100630 91160
rect 99748 89616 99800 89622
rect 99748 89558 99800 89564
rect 100588 85338 100616 91151
rect 100576 85332 100628 85338
rect 100576 85274 100628 85280
rect 101876 84046 101904 91287
rect 101954 91216 102010 91225
rect 101954 91151 102010 91160
rect 101864 84040 101916 84046
rect 101864 83982 101916 83988
rect 101968 82793 101996 91151
rect 101954 82784 102010 82793
rect 101954 82719 102010 82728
rect 99288 78532 99340 78538
rect 99288 78474 99340 78480
rect 99196 78464 99248 78470
rect 99196 78406 99248 78412
rect 95148 75880 95200 75886
rect 95148 75822 95200 75828
rect 102060 75818 102088 91423
rect 103164 89486 103192 91559
rect 107566 91352 107622 91361
rect 107566 91287 107622 91296
rect 103426 91216 103482 91225
rect 103426 91151 103482 91160
rect 104346 91216 104402 91225
rect 104346 91151 104402 91160
rect 104622 91216 104678 91225
rect 104622 91151 104678 91160
rect 107474 91216 107530 91225
rect 107474 91151 107530 91160
rect 103152 89480 103204 89486
rect 103152 89422 103204 89428
rect 103440 79898 103468 91151
rect 104360 85406 104388 91151
rect 104636 88233 104664 91151
rect 104622 88224 104678 88233
rect 104622 88159 104678 88168
rect 104348 85400 104400 85406
rect 104348 85342 104400 85348
rect 107488 84114 107516 91151
rect 107476 84108 107528 84114
rect 107476 84050 107528 84056
rect 107580 80073 107608 91287
rect 107764 90982 107792 92375
rect 109222 91216 109278 91225
rect 109222 91151 109278 91160
rect 109774 91216 109830 91225
rect 109774 91151 109830 91160
rect 108304 91112 108356 91118
rect 108304 91054 108356 91060
rect 107752 90976 107804 90982
rect 107752 90918 107804 90924
rect 108316 81394 108344 91054
rect 109236 88126 109264 91151
rect 109224 88120 109276 88126
rect 109224 88062 109276 88068
rect 109788 86834 109816 91151
rect 109776 86828 109828 86834
rect 109776 86770 109828 86776
rect 110340 82686 110368 93191
rect 128174 93191 128230 93200
rect 110696 93162 110748 93168
rect 125508 93152 125560 93158
rect 125508 93094 125560 93100
rect 115480 92472 115532 92478
rect 114190 92440 114246 92449
rect 114190 92375 114246 92384
rect 115478 92440 115480 92449
rect 115532 92440 115534 92449
rect 115478 92375 115534 92384
rect 116766 92440 116822 92449
rect 116766 92375 116768 92384
rect 111614 91216 111670 91225
rect 111614 91151 111670 91160
rect 111982 91216 112038 91225
rect 111982 91151 112038 91160
rect 112350 91216 112406 91225
rect 112350 91151 112406 91160
rect 111628 85542 111656 91151
rect 111996 88194 112024 91151
rect 111984 88188 112036 88194
rect 111984 88130 112036 88136
rect 112364 86766 112392 91151
rect 114204 91050 114232 92375
rect 116820 92375 116822 92384
rect 119710 92440 119766 92449
rect 119710 92375 119766 92384
rect 122470 92440 122526 92449
rect 122470 92375 122526 92384
rect 116768 92346 116820 92352
rect 119724 92206 119752 92375
rect 119712 92200 119764 92206
rect 119712 92142 119764 92148
rect 117134 91760 117190 91769
rect 117134 91695 117190 91704
rect 114466 91216 114522 91225
rect 114466 91151 114522 91160
rect 115294 91216 115350 91225
rect 115294 91151 115350 91160
rect 114192 91044 114244 91050
rect 114192 90986 114244 90992
rect 112352 86760 112404 86766
rect 112352 86702 112404 86708
rect 111616 85536 111668 85542
rect 111616 85478 111668 85484
rect 110328 82680 110380 82686
rect 110328 82622 110380 82628
rect 108304 81388 108356 81394
rect 108304 81330 108356 81336
rect 107566 80064 107622 80073
rect 107566 79999 107622 80008
rect 114480 79966 114508 91151
rect 115308 88262 115336 91151
rect 117148 89418 117176 91695
rect 121274 91352 121330 91361
rect 121274 91287 121330 91296
rect 118606 91216 118662 91225
rect 118606 91151 118662 91160
rect 117136 89412 117188 89418
rect 117136 89354 117188 89360
rect 115296 88256 115348 88262
rect 115296 88198 115348 88204
rect 118620 83978 118648 91151
rect 121288 84017 121316 91287
rect 121366 91216 121422 91225
rect 121366 91151 121422 91160
rect 121274 84008 121330 84017
rect 118608 83972 118660 83978
rect 121274 83943 121330 83952
rect 118608 83914 118660 83920
rect 121380 82618 121408 91151
rect 122484 90846 122512 92375
rect 125520 92342 125548 93094
rect 125782 92440 125838 92449
rect 125782 92375 125838 92384
rect 125508 92336 125560 92342
rect 125508 92278 125560 92284
rect 125506 92168 125562 92177
rect 125796 92138 125824 92375
rect 125506 92103 125562 92112
rect 125784 92132 125836 92138
rect 122838 91488 122894 91497
rect 122838 91423 122894 91432
rect 122746 91216 122802 91225
rect 122746 91151 122802 91160
rect 122472 90840 122524 90846
rect 122472 90782 122524 90788
rect 121368 82612 121420 82618
rect 121368 82554 121420 82560
rect 114468 79960 114520 79966
rect 114468 79902 114520 79908
rect 103428 79892 103480 79898
rect 103428 79834 103480 79840
rect 122760 78606 122788 91151
rect 122852 85270 122880 91423
rect 123574 91216 123630 91225
rect 123574 91151 123630 91160
rect 124126 91216 124182 91225
rect 124126 91151 124182 91160
rect 125414 91216 125470 91225
rect 125414 91151 125470 91160
rect 123588 86873 123616 91151
rect 123574 86864 123630 86873
rect 123574 86799 123630 86808
rect 124140 86698 124168 91151
rect 124128 86692 124180 86698
rect 124128 86634 124180 86640
rect 122840 85264 122892 85270
rect 122840 85206 122892 85212
rect 125428 81122 125456 91151
rect 125520 90778 125548 92103
rect 125784 92074 125836 92080
rect 126518 91216 126574 91225
rect 126518 91151 126574 91160
rect 126886 91216 126942 91225
rect 126886 91151 126942 91160
rect 125508 90772 125560 90778
rect 125508 90714 125560 90720
rect 126532 87990 126560 91151
rect 126520 87984 126572 87990
rect 126520 87926 126572 87932
rect 126900 82550 126928 91151
rect 128188 89729 128216 93191
rect 151542 92440 151598 92449
rect 151542 92375 151598 92384
rect 152094 92440 152150 92449
rect 152094 92375 152150 92384
rect 151556 92342 151584 92375
rect 151544 92336 151596 92342
rect 151544 92278 151596 92284
rect 152108 92274 152136 92375
rect 152096 92268 152148 92274
rect 152096 92210 152148 92216
rect 151450 92168 151506 92177
rect 151450 92103 151506 92112
rect 136454 91488 136510 91497
rect 136454 91423 136510 91432
rect 132038 91216 132094 91225
rect 132038 91151 132094 91160
rect 133142 91216 133198 91225
rect 133142 91151 133198 91160
rect 128174 89720 128230 89729
rect 128174 89655 128230 89664
rect 132052 85202 132080 91151
rect 133156 88058 133184 91151
rect 136468 89350 136496 91423
rect 151464 90914 151492 92103
rect 151452 90908 151504 90914
rect 151452 90850 151504 90856
rect 136456 89344 136508 89350
rect 136456 89286 136508 89292
rect 133144 88052 133196 88058
rect 133144 87994 133196 88000
rect 164896 85474 164924 96630
rect 166276 90846 166304 139402
rect 166356 125656 166408 125662
rect 166356 125598 166408 125604
rect 166264 90840 166316 90846
rect 166264 90782 166316 90788
rect 166368 90778 166396 125598
rect 167644 120148 167696 120154
rect 167644 120090 167696 120096
rect 166448 118720 166500 118726
rect 166448 118662 166500 118668
rect 166356 90772 166408 90778
rect 166356 90714 166408 90720
rect 166460 86766 166488 118662
rect 166540 97300 166592 97306
rect 166540 97242 166592 97248
rect 166552 92206 166580 97242
rect 167656 93294 167684 120090
rect 167736 117972 167788 117978
rect 167736 117914 167788 117920
rect 167748 108769 167776 117914
rect 168196 115252 168248 115258
rect 168196 115194 168248 115200
rect 167920 111784 167972 111790
rect 167918 111752 167920 111761
rect 167972 111752 167974 111761
rect 167918 111687 167974 111696
rect 168208 110129 168236 115194
rect 168194 110120 168250 110129
rect 168194 110055 168250 110064
rect 167734 108760 167790 108769
rect 167734 108695 167790 108704
rect 167736 106344 167788 106350
rect 167736 106286 167788 106292
rect 167644 93288 167696 93294
rect 167644 93230 167696 93236
rect 166540 92200 166592 92206
rect 166540 92142 166592 92148
rect 166448 86760 166500 86766
rect 166448 86702 166500 86708
rect 164884 85468 164936 85474
rect 164884 85410 164936 85416
rect 132040 85196 132092 85202
rect 132040 85138 132092 85144
rect 126888 82544 126940 82550
rect 126888 82486 126940 82492
rect 167748 81190 167776 106286
rect 167920 99408 167972 99414
rect 167920 99350 167972 99356
rect 167828 98048 167880 98054
rect 167828 97990 167880 97996
rect 167840 81258 167868 97990
rect 167932 89554 167960 99350
rect 167920 89548 167972 89554
rect 167920 89490 167972 89496
rect 169036 82550 169064 142122
rect 169116 133952 169168 133958
rect 169116 133894 169168 133900
rect 169128 93226 169156 133894
rect 169208 125724 169260 125730
rect 169208 125666 169260 125672
rect 169116 93220 169168 93226
rect 169116 93162 169168 93168
rect 169220 87990 169248 125666
rect 169300 116000 169352 116006
rect 169300 115942 169352 115948
rect 169312 88126 169340 115942
rect 170416 89350 170444 147630
rect 170496 146328 170548 146334
rect 170496 146270 170548 146276
rect 170508 94178 170536 146270
rect 173164 144968 173216 144974
rect 173164 144910 173216 144916
rect 171784 142248 171836 142254
rect 171784 142190 171836 142196
rect 170588 124228 170640 124234
rect 170588 124170 170640 124176
rect 170496 94172 170548 94178
rect 170496 94114 170548 94120
rect 170404 89344 170456 89350
rect 170404 89286 170456 89292
rect 169300 88120 169352 88126
rect 169300 88062 169352 88068
rect 169208 87984 169260 87990
rect 169208 87926 169260 87932
rect 170600 86698 170628 124170
rect 170680 111852 170732 111858
rect 170680 111794 170732 111800
rect 170588 86692 170640 86698
rect 170588 86634 170640 86640
rect 170692 85338 170720 111794
rect 171796 92138 171824 142190
rect 171876 138032 171928 138038
rect 171876 137974 171928 137980
rect 171888 94110 171916 137974
rect 171968 113212 172020 113218
rect 171968 113154 172020 113160
rect 171876 94104 171928 94110
rect 171876 94046 171928 94052
rect 171784 92132 171836 92138
rect 171784 92074 171836 92080
rect 171980 89486 172008 113154
rect 172060 100768 172112 100774
rect 172060 100710 172112 100716
rect 171968 89480 172020 89486
rect 171968 89422 172020 89428
rect 170680 85332 170732 85338
rect 170680 85274 170732 85280
rect 169024 82544 169076 82550
rect 169024 82486 169076 82492
rect 167828 81252 167880 81258
rect 167828 81194 167880 81200
rect 167736 81184 167788 81190
rect 167736 81126 167788 81132
rect 125416 81116 125468 81122
rect 125416 81058 125468 81064
rect 122748 78600 122800 78606
rect 122748 78542 122800 78548
rect 172072 77246 172100 100710
rect 173176 93362 173204 144910
rect 174544 143608 174596 143614
rect 174544 143550 174596 143556
rect 173256 128376 173308 128382
rect 173256 128318 173308 128324
rect 173164 93356 173216 93362
rect 173164 93298 173216 93304
rect 173268 78470 173296 128318
rect 173348 124296 173400 124302
rect 173348 124238 173400 124244
rect 173360 85270 173388 124238
rect 173440 99476 173492 99482
rect 173440 99418 173492 99424
rect 173452 86902 173480 99418
rect 174556 89729 174584 143550
rect 174820 137284 174872 137290
rect 174820 137226 174872 137232
rect 174636 135312 174688 135318
rect 174636 135254 174688 135260
rect 174542 89720 174598 89729
rect 174542 89655 174598 89664
rect 174648 88194 174676 135254
rect 174728 122868 174780 122874
rect 174728 122810 174780 122816
rect 174636 88188 174688 88194
rect 174636 88130 174688 88136
rect 173440 86896 173492 86902
rect 173440 86838 173492 86844
rect 173348 85264 173400 85270
rect 173348 85206 173400 85212
rect 174740 82618 174768 122810
rect 174832 111790 174860 137226
rect 174820 111784 174872 111790
rect 174820 111726 174872 111732
rect 174820 107704 174872 107710
rect 174820 107646 174872 107652
rect 174728 82612 174780 82618
rect 174728 82554 174780 82560
rect 174832 79830 174860 107646
rect 174820 79824 174872 79830
rect 174820 79766 174872 79772
rect 173256 78464 173308 78470
rect 173256 78406 173308 78412
rect 172060 77240 172112 77246
rect 172060 77182 172112 77188
rect 102048 75812 102100 75818
rect 102048 75754 102100 75760
rect 107660 75200 107712 75206
rect 107660 75142 107712 75148
rect 103520 73908 103572 73914
rect 103520 73850 103572 73856
rect 93860 61396 93912 61402
rect 93860 61338 93912 61344
rect 92480 54596 92532 54602
rect 92480 54538 92532 54544
rect 91100 40792 91152 40798
rect 91100 40734 91152 40740
rect 91112 16574 91140 40734
rect 85684 16546 86448 16574
rect 86972 16546 87552 16574
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 91112 16546 91600 16574
rect 85592 6886 85712 6914
rect 85684 480 85712 6886
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86420 354 86448 16546
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 87524 354 87552 16546
rect 89180 480 89208 16546
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 54538
rect 93872 3602 93900 61338
rect 99380 53168 99432 53174
rect 99380 53110 99432 53116
rect 98000 42084 98052 42090
rect 98000 42026 98052 42032
rect 95240 39432 95292 39438
rect 95240 39374 95292 39380
rect 93952 24200 94004 24206
rect 93952 24142 94004 24148
rect 93860 3596 93912 3602
rect 93860 3538 93912 3544
rect 93964 480 93992 24142
rect 95252 16574 95280 39374
rect 98012 16574 98040 42026
rect 99392 16574 99420 53110
rect 102140 44940 102192 44946
rect 102140 44882 102192 44888
rect 100760 25628 100812 25634
rect 100760 25570 100812 25576
rect 95252 16546 95832 16574
rect 98012 16546 98224 16574
rect 99392 16546 99880 16574
rect 94780 3596 94832 3602
rect 94780 3538 94832 3544
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94792 354 94820 3538
rect 95118 354 95230 480
rect 94792 326 95230 354
rect 95804 354 95832 16546
rect 97448 4888 97500 4894
rect 97448 4830 97500 4836
rect 97460 480 97488 4830
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 25570
rect 102152 16574 102180 44882
rect 103532 16574 103560 73850
rect 106280 46232 106332 46238
rect 106280 46174 106332 46180
rect 106292 16574 106320 46174
rect 107672 16574 107700 75142
rect 122840 72548 122892 72554
rect 122840 72490 122892 72496
rect 118700 60036 118752 60042
rect 118700 59978 118752 59984
rect 110420 58744 110472 58750
rect 110420 58686 110472 58692
rect 102152 16546 102272 16574
rect 103532 16546 104112 16574
rect 106292 16546 106504 16574
rect 107672 16546 108160 16574
rect 102244 480 102272 16546
rect 103336 3596 103388 3602
rect 103336 3538 103388 3544
rect 103348 480 103376 3538
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105728 14476 105780 14482
rect 105728 14418 105780 14424
rect 105740 480 105768 14418
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108132 480 108160 16546
rect 110432 3534 110460 58686
rect 112442 43480 112498 43489
rect 112442 43415 112498 43424
rect 110512 10396 110564 10402
rect 110512 10338 110564 10344
rect 110420 3528 110472 3534
rect 110420 3470 110472 3476
rect 109316 2168 109368 2174
rect 109316 2110 109368 2116
rect 109328 480 109356 2110
rect 110524 480 110552 10338
rect 112456 3602 112484 43415
rect 113180 33856 113232 33862
rect 113180 33798 113232 33804
rect 113192 16574 113220 33798
rect 114560 28348 114612 28354
rect 114560 28290 114612 28296
rect 114572 16574 114600 28290
rect 115940 19984 115992 19990
rect 115940 19926 115992 19932
rect 115952 16574 115980 19926
rect 113192 16546 114048 16574
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 112812 3664 112864 3670
rect 112812 3606 112864 3612
rect 112444 3596 112496 3602
rect 112444 3538 112496 3544
rect 111616 3528 111668 3534
rect 111616 3470 111668 3476
rect 111628 480 111656 3470
rect 112824 480 112852 3606
rect 114020 480 114048 16546
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 117320 11824 117372 11830
rect 117320 11766 117372 11772
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 11766
rect 118712 3534 118740 59978
rect 118792 29708 118844 29714
rect 118792 29650 118844 29656
rect 118700 3528 118752 3534
rect 118700 3470 118752 3476
rect 118804 480 118832 29650
rect 121460 26988 121512 26994
rect 121460 26930 121512 26936
rect 121472 16574 121500 26930
rect 122852 16574 122880 72490
rect 175936 60722 175964 229842
rect 178696 184385 178724 295530
rect 180062 294264 180118 294273
rect 180062 294199 180118 294208
rect 178682 184376 178738 184385
rect 178682 184311 178738 184320
rect 178684 153264 178736 153270
rect 178684 153206 178736 153212
rect 176016 145036 176068 145042
rect 176016 144978 176068 144984
rect 176028 85202 176056 144978
rect 176108 133204 176160 133210
rect 176108 133146 176160 133152
rect 176120 92410 176148 133146
rect 177304 127016 177356 127022
rect 177304 126958 177356 126964
rect 176108 92404 176160 92410
rect 176108 92346 176160 92352
rect 176016 85196 176068 85202
rect 176016 85138 176068 85144
rect 177316 78538 177344 126958
rect 177396 111920 177448 111926
rect 177396 111862 177448 111868
rect 177304 78532 177356 78538
rect 177304 78474 177356 78480
rect 177408 75818 177436 111862
rect 178696 93430 178724 153206
rect 178868 150476 178920 150482
rect 178868 150418 178920 150424
rect 178776 127084 178828 127090
rect 178776 127026 178828 127032
rect 178684 93424 178736 93430
rect 178684 93366 178736 93372
rect 178788 81326 178816 127026
rect 178880 115258 178908 150418
rect 178868 115252 178920 115258
rect 178868 115194 178920 115200
rect 178960 114572 179012 114578
rect 178960 114514 179012 114520
rect 178972 94042 179000 114514
rect 180076 95169 180104 294199
rect 184216 178770 184244 299678
rect 185596 185774 185624 303758
rect 189724 302320 189776 302326
rect 189724 302262 189776 302268
rect 188344 238128 188396 238134
rect 188344 238070 188396 238076
rect 185584 185768 185636 185774
rect 185584 185710 185636 185716
rect 184204 178764 184256 178770
rect 184204 178706 184256 178712
rect 184848 151088 184900 151094
rect 184848 151030 184900 151036
rect 184860 150346 184888 151030
rect 184848 150340 184900 150346
rect 184848 150282 184900 150288
rect 181444 146396 181496 146402
rect 181444 146338 181496 146344
rect 180156 131164 180208 131170
rect 180156 131106 180208 131112
rect 180062 95160 180118 95169
rect 180062 95095 180118 95104
rect 178960 94036 179012 94042
rect 178960 93978 179012 93984
rect 180168 92313 180196 131106
rect 180248 121508 180300 121514
rect 180248 121450 180300 121456
rect 180154 92304 180210 92313
rect 180154 92239 180210 92248
rect 180064 91792 180116 91798
rect 180064 91734 180116 91740
rect 178776 81320 178828 81326
rect 178776 81262 178828 81268
rect 177396 75812 177448 75818
rect 177396 75754 177448 75760
rect 175924 60716 175976 60722
rect 175924 60658 175976 60664
rect 121472 16546 122328 16574
rect 122852 16546 123064 16574
rect 119896 3528 119948 3534
rect 119896 3470 119948 3476
rect 121092 3528 121144 3534
rect 121092 3470 121144 3476
rect 119908 480 119936 3470
rect 121104 480 121132 3470
rect 122300 480 122328 16546
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 124680 13184 124732 13190
rect 124680 13126 124732 13132
rect 124692 480 124720 13126
rect 180076 3670 180104 91734
rect 180260 83978 180288 121450
rect 181456 88058 181484 146338
rect 185584 120216 185636 120222
rect 185584 120158 185636 120164
rect 184204 113280 184256 113286
rect 184204 113222 184256 113228
rect 181444 88052 181496 88058
rect 181444 87994 181496 88000
rect 184216 85406 184244 113222
rect 185596 89418 185624 120158
rect 188356 93770 188384 238070
rect 189736 180033 189764 302262
rect 192484 298376 192536 298382
rect 192484 298318 192536 298324
rect 192496 188426 192524 298318
rect 210424 297016 210476 297022
rect 210424 296958 210476 296964
rect 196624 295520 196676 295526
rect 196624 295462 196676 295468
rect 193128 285728 193180 285734
rect 193128 285670 193180 285676
rect 193140 282198 193168 285670
rect 193128 282192 193180 282198
rect 193128 282134 193180 282140
rect 192576 233980 192628 233986
rect 192576 233922 192628 233928
rect 192588 210526 192616 233922
rect 192576 210520 192628 210526
rect 192576 210462 192628 210468
rect 192484 188420 192536 188426
rect 192484 188362 192536 188368
rect 189722 180024 189778 180033
rect 189722 179959 189778 179968
rect 196636 176662 196664 295462
rect 202144 289128 202196 289134
rect 202144 289070 202196 289076
rect 198004 254040 198056 254046
rect 198004 253982 198056 253988
rect 196716 199640 196768 199646
rect 196716 199582 196768 199588
rect 196624 176656 196676 176662
rect 196624 176598 196676 176604
rect 193864 140820 193916 140826
rect 193864 140762 193916 140768
rect 192484 134020 192536 134026
rect 192484 133962 192536 133968
rect 189724 129804 189776 129810
rect 189724 129746 189776 129752
rect 188344 93764 188396 93770
rect 188344 93706 188396 93712
rect 185584 89412 185636 89418
rect 185584 89354 185636 89360
rect 184204 85400 184256 85406
rect 184204 85342 184256 85348
rect 180248 83972 180300 83978
rect 180248 83914 180300 83920
rect 189736 79898 189764 129746
rect 189816 116068 189868 116074
rect 189816 116010 189868 116016
rect 189828 90982 189856 116010
rect 189816 90976 189868 90982
rect 189816 90918 189868 90924
rect 192496 86834 192524 133962
rect 192484 86828 192536 86834
rect 192484 86770 192536 86776
rect 193876 81122 193904 140762
rect 196624 118788 196676 118794
rect 196624 118730 196676 118736
rect 196636 88262 196664 118730
rect 196728 95198 196756 199582
rect 198016 187066 198044 253982
rect 198004 187060 198056 187066
rect 198004 187002 198056 187008
rect 202156 181626 202184 289070
rect 206284 278860 206336 278866
rect 206284 278802 206336 278808
rect 203524 249824 203576 249830
rect 203524 249766 203576 249772
rect 202144 181620 202196 181626
rect 202144 181562 202196 181568
rect 203536 177410 203564 249766
rect 206296 178838 206324 278802
rect 207664 269204 207716 269210
rect 207664 269146 207716 269152
rect 207676 188494 207704 269146
rect 207664 188488 207716 188494
rect 207664 188430 207716 188436
rect 207756 187740 207808 187746
rect 207756 187682 207808 187688
rect 206284 178832 206336 178838
rect 206284 178774 206336 178780
rect 203524 177404 203576 177410
rect 203524 177346 203576 177352
rect 207768 161362 207796 187682
rect 208400 178084 208452 178090
rect 208400 178026 208452 178032
rect 208412 172446 208440 178026
rect 210436 175953 210464 296958
rect 211804 273284 211856 273290
rect 211804 273226 211856 273232
rect 211816 183122 211844 273226
rect 214576 231810 214604 699654
rect 224224 303748 224276 303754
rect 224224 303690 224276 303696
rect 215944 294296 215996 294302
rect 215944 294238 215996 294244
rect 214564 231804 214616 231810
rect 214564 231746 214616 231752
rect 214564 224256 214616 224262
rect 214564 224198 214616 224204
rect 211896 189100 211948 189106
rect 211896 189042 211948 189048
rect 211804 183116 211856 183122
rect 211804 183058 211856 183064
rect 211804 180872 211856 180878
rect 211804 180814 211856 180820
rect 210516 175976 210568 175982
rect 210422 175944 210478 175953
rect 210516 175918 210568 175924
rect 210422 175879 210478 175888
rect 208400 172440 208452 172446
rect 208400 172382 208452 172388
rect 207756 161356 207808 161362
rect 207756 161298 207808 161304
rect 210528 157282 210556 175918
rect 211816 169658 211844 180814
rect 211804 169652 211856 169658
rect 211804 169594 211856 169600
rect 211908 160070 211936 189042
rect 214576 188329 214604 224198
rect 214562 188320 214618 188329
rect 214562 188255 214618 188264
rect 214656 186380 214708 186386
rect 214656 186322 214708 186328
rect 213920 176792 213972 176798
rect 213920 176734 213972 176740
rect 211988 176724 212040 176730
rect 211988 176666 212040 176672
rect 212000 171018 212028 176666
rect 213932 175681 213960 176734
rect 214564 176112 214616 176118
rect 214564 176054 214616 176060
rect 214104 176044 214156 176050
rect 214104 175986 214156 175992
rect 213918 175672 213974 175681
rect 213918 175607 213974 175616
rect 213920 175228 213972 175234
rect 213920 175170 213972 175176
rect 213932 175001 213960 175170
rect 214012 175160 214064 175166
rect 214012 175102 214064 175108
rect 213918 174992 213974 175001
rect 213918 174927 213974 174936
rect 214024 174321 214052 175102
rect 214010 174312 214066 174321
rect 214010 174247 214066 174256
rect 213920 173868 213972 173874
rect 213920 173810 213972 173816
rect 213932 173641 213960 173810
rect 213918 173632 213974 173641
rect 213918 173567 213974 173576
rect 214116 172961 214144 175986
rect 214102 172952 214158 172961
rect 214102 172887 214158 172896
rect 214012 172508 214064 172514
rect 214012 172450 214064 172456
rect 213920 172440 213972 172446
rect 213920 172382 213972 172388
rect 213932 172281 213960 172382
rect 213918 172272 213974 172281
rect 213918 172207 213974 172216
rect 214024 171601 214052 172450
rect 214010 171592 214066 171601
rect 214010 171527 214066 171536
rect 213920 171080 213972 171086
rect 213920 171022 213972 171028
rect 214010 171048 214066 171057
rect 211988 171012 212040 171018
rect 211988 170954 212040 170960
rect 213932 170377 213960 171022
rect 214010 170983 214012 170992
rect 214064 170983 214066 170992
rect 214012 170954 214064 170960
rect 213918 170368 213974 170377
rect 213918 170303 213974 170312
rect 213920 169720 213972 169726
rect 213920 169662 213972 169668
rect 214010 169688 214066 169697
rect 213932 169017 213960 169662
rect 214010 169623 214012 169632
rect 214064 169623 214066 169632
rect 214012 169594 214064 169600
rect 213918 169008 213974 169017
rect 213918 168943 213974 168952
rect 214012 168360 214064 168366
rect 213918 168328 213974 168337
rect 214012 168302 214064 168308
rect 213918 168263 213920 168272
rect 213972 168263 213974 168272
rect 213920 168234 213972 168240
rect 214024 167657 214052 168302
rect 214010 167648 214066 167657
rect 214010 167583 214066 167592
rect 213920 167000 213972 167006
rect 213918 166968 213920 166977
rect 213972 166968 213974 166977
rect 213918 166903 213974 166912
rect 214012 166932 214064 166938
rect 214012 166874 214064 166880
rect 214024 166433 214052 166874
rect 214010 166424 214066 166433
rect 214010 166359 214066 166368
rect 213920 165572 213972 165578
rect 213920 165514 213972 165520
rect 213932 165073 213960 165514
rect 214012 165504 214064 165510
rect 214012 165446 214064 165452
rect 213918 165064 213974 165073
rect 213918 164999 213974 165008
rect 214024 164393 214052 165446
rect 214010 164384 214066 164393
rect 214010 164319 214066 164328
rect 213920 164212 213972 164218
rect 213920 164154 213972 164160
rect 213932 163033 213960 164154
rect 213918 163024 213974 163033
rect 213918 162959 213974 162968
rect 213920 162852 213972 162858
rect 213920 162794 213972 162800
rect 213932 162353 213960 162794
rect 213918 162344 213974 162353
rect 213918 162279 213974 162288
rect 213920 161424 213972 161430
rect 213920 161366 213972 161372
rect 213932 161129 213960 161366
rect 214012 161356 214064 161362
rect 214012 161298 214064 161304
rect 213918 161120 213974 161129
rect 213918 161055 213974 161064
rect 213920 160744 213972 160750
rect 213920 160686 213972 160692
rect 211896 160064 211948 160070
rect 211896 160006 211948 160012
rect 213932 157729 213960 160686
rect 214024 160449 214052 161298
rect 214010 160440 214066 160449
rect 214010 160375 214066 160384
rect 214472 160064 214524 160070
rect 214472 160006 214524 160012
rect 214484 159769 214512 160006
rect 214470 159760 214526 159769
rect 214470 159695 214526 159704
rect 213918 157720 213974 157729
rect 213918 157655 213974 157664
rect 213920 157344 213972 157350
rect 213920 157286 213972 157292
rect 210516 157276 210568 157282
rect 210516 157218 210568 157224
rect 213932 156505 213960 157286
rect 214012 157276 214064 157282
rect 214012 157218 214064 157224
rect 214024 157185 214052 157218
rect 214010 157176 214066 157185
rect 214010 157111 214066 157120
rect 213918 156496 213974 156505
rect 213918 156431 213974 156440
rect 213920 155916 213972 155922
rect 213920 155858 213972 155864
rect 213932 155825 213960 155858
rect 213918 155816 213974 155825
rect 213918 155751 213974 155760
rect 213918 154456 213974 154465
rect 213918 154391 213974 154400
rect 213932 153270 213960 154391
rect 213920 153264 213972 153270
rect 213920 153206 213972 153212
rect 214010 153096 214066 153105
rect 214010 153031 214066 153040
rect 213918 152552 213974 152561
rect 213918 152487 213974 152496
rect 213932 151978 213960 152487
rect 202144 151972 202196 151978
rect 202144 151914 202196 151920
rect 213920 151972 213972 151978
rect 213920 151914 213972 151920
rect 198004 128444 198056 128450
rect 198004 128386 198056 128392
rect 196716 95192 196768 95198
rect 196716 95134 196768 95140
rect 196624 88256 196676 88262
rect 196624 88198 196676 88204
rect 198016 84046 198044 128386
rect 199384 110492 199436 110498
rect 199384 110434 199436 110440
rect 199396 89622 199424 110434
rect 202156 92274 202184 151914
rect 214024 151910 214052 153031
rect 206284 151904 206336 151910
rect 214012 151904 214064 151910
rect 206284 151846 206336 151852
rect 213274 151872 213330 151881
rect 203524 136672 203576 136678
rect 203524 136614 203576 136620
rect 202236 110560 202288 110566
rect 202236 110502 202288 110508
rect 202144 92268 202196 92274
rect 202144 92210 202196 92216
rect 199384 89616 199436 89622
rect 199384 89558 199436 89564
rect 198004 84040 198056 84046
rect 198004 83982 198056 83988
rect 202248 82754 202276 110502
rect 203536 92478 203564 136614
rect 203616 107772 203668 107778
rect 203616 107714 203668 107720
rect 203524 92472 203576 92478
rect 203524 92414 203576 92420
rect 202236 82748 202288 82754
rect 202236 82690 202288 82696
rect 193864 81116 193916 81122
rect 193864 81058 193916 81064
rect 189724 79892 189776 79898
rect 189724 79834 189776 79840
rect 203628 75886 203656 107714
rect 204904 102196 204956 102202
rect 204904 102138 204956 102144
rect 204916 82822 204944 102138
rect 206296 92342 206324 151846
rect 214012 151846 214064 151852
rect 213274 151807 213330 151816
rect 210424 143676 210476 143682
rect 210424 143618 210476 143624
rect 207756 135380 207808 135386
rect 207756 135322 207808 135328
rect 207664 121576 207716 121582
rect 207664 121518 207716 121524
rect 206376 109064 206428 109070
rect 206376 109006 206428 109012
rect 206284 92336 206336 92342
rect 206284 92278 206336 92284
rect 204904 82816 204956 82822
rect 204904 82758 204956 82764
rect 206388 78674 206416 109006
rect 207676 93906 207704 121518
rect 207664 93900 207716 93906
rect 207664 93842 207716 93848
rect 207768 91050 207796 135322
rect 209044 104916 209096 104922
rect 209044 104858 209096 104864
rect 207848 100836 207900 100842
rect 207848 100778 207900 100784
rect 207756 91044 207808 91050
rect 207756 90986 207808 90992
rect 207664 90364 207716 90370
rect 207664 90306 207716 90312
rect 206376 78668 206428 78674
rect 206376 78610 206428 78616
rect 203616 75880 203668 75886
rect 203616 75822 203668 75828
rect 180064 3664 180116 3670
rect 180064 3606 180116 3612
rect 207676 3602 207704 90306
rect 207860 80034 207888 100778
rect 209056 93838 209084 104858
rect 209136 103556 209188 103562
rect 209136 103498 209188 103504
rect 209148 94897 209176 103498
rect 209134 94888 209190 94897
rect 209134 94823 209190 94832
rect 210436 93974 210464 143618
rect 211896 132932 211948 132938
rect 211896 132874 211948 132880
rect 211804 123412 211856 123418
rect 211804 123354 211856 123360
rect 210516 118856 210568 118862
rect 210516 118798 210568 118804
rect 210424 93968 210476 93974
rect 210424 93910 210476 93916
rect 209044 93832 209096 93838
rect 209044 93774 209096 93780
rect 207848 80028 207900 80034
rect 207848 79970 207900 79976
rect 210528 79966 210556 118798
rect 210608 117360 210660 117366
rect 210608 117302 210660 117308
rect 210620 85542 210648 117302
rect 210608 85536 210660 85542
rect 210608 85478 210660 85484
rect 210516 79960 210568 79966
rect 210516 79902 210568 79908
rect 211816 78606 211844 123354
rect 211908 91633 211936 132874
rect 213288 117978 213316 151807
rect 214010 151192 214066 151201
rect 214010 151127 214066 151136
rect 214024 150482 214052 151127
rect 214012 150476 214064 150482
rect 214012 150418 214064 150424
rect 213920 150408 213972 150414
rect 213920 150350 213972 150356
rect 213932 149841 213960 150350
rect 214012 150340 214064 150346
rect 214012 150282 214064 150288
rect 213918 149832 213974 149841
rect 213918 149767 213974 149776
rect 214024 149161 214052 150282
rect 214010 149152 214066 149161
rect 214010 149087 214066 149096
rect 214576 148481 214604 176054
rect 214668 165753 214696 186322
rect 215956 181694 215984 294238
rect 220084 292868 220136 292874
rect 220084 292810 220136 292816
rect 215944 181688 215996 181694
rect 215944 181630 215996 181636
rect 220096 180334 220124 292810
rect 224236 191282 224264 303690
rect 225604 299668 225656 299674
rect 225604 299610 225656 299616
rect 224316 213376 224368 213382
rect 224316 213318 224368 213324
rect 224224 191276 224276 191282
rect 224224 191218 224276 191224
rect 220084 180328 220136 180334
rect 220084 180270 220136 180276
rect 224328 180169 224356 213318
rect 224314 180160 224370 180169
rect 224314 180095 224370 180104
rect 214748 179444 214800 179450
rect 214748 179386 214800 179392
rect 214654 165744 214710 165753
rect 214654 165679 214710 165688
rect 214760 161809 214788 179386
rect 225616 178974 225644 299610
rect 248420 296948 248472 296954
rect 248420 296890 248472 296896
rect 246304 289944 246356 289950
rect 246304 289886 246356 289892
rect 242164 281580 242216 281586
rect 242164 281522 242216 281528
rect 238024 280288 238076 280294
rect 238024 280230 238076 280236
rect 232504 256760 232556 256766
rect 232504 256702 232556 256708
rect 229744 247104 229796 247110
rect 229744 247046 229796 247052
rect 228364 218816 228416 218822
rect 228364 218758 228416 218764
rect 225604 178968 225656 178974
rect 225604 178910 225656 178916
rect 228376 177478 228404 218758
rect 229756 178906 229784 247046
rect 229744 178900 229796 178906
rect 229744 178842 229796 178848
rect 232516 177614 232544 256702
rect 233884 252680 233936 252686
rect 233884 252622 233936 252628
rect 233896 183190 233924 252622
rect 233884 183184 233936 183190
rect 233884 183126 233936 183132
rect 238036 179110 238064 280230
rect 239404 269136 239456 269142
rect 239404 269078 239456 269084
rect 238024 179104 238076 179110
rect 238024 179046 238076 179052
rect 232504 177608 232556 177614
rect 232504 177550 232556 177556
rect 239416 177546 239444 269078
rect 240784 195424 240836 195430
rect 240784 195366 240836 195372
rect 239404 177540 239456 177546
rect 239404 177482 239456 177488
rect 228364 177472 228416 177478
rect 228364 177414 228416 177420
rect 240796 176089 240824 195366
rect 242176 176594 242204 281522
rect 242256 204944 242308 204950
rect 242256 204886 242308 204892
rect 242164 176588 242216 176594
rect 242164 176530 242216 176536
rect 240782 176080 240838 176089
rect 242268 176050 242296 204886
rect 242808 178764 242860 178770
rect 242808 178706 242860 178712
rect 242820 177682 242848 178706
rect 242808 177676 242860 177682
rect 242808 177618 242860 177624
rect 240782 176015 240838 176024
rect 242256 176044 242308 176050
rect 242256 175986 242308 175992
rect 246316 175982 246344 289886
rect 247684 276140 247736 276146
rect 247684 276082 247736 276088
rect 247696 247722 247724 276082
rect 247684 247716 247736 247722
rect 247684 247658 247736 247664
rect 248432 177585 248460 296890
rect 255320 294228 255372 294234
rect 255320 294170 255372 294176
rect 253940 274712 253992 274718
rect 253940 274654 253992 274660
rect 249800 270564 249852 270570
rect 249800 270506 249852 270512
rect 249064 178832 249116 178838
rect 249064 178774 249116 178780
rect 248418 177576 248474 177585
rect 248418 177511 248474 177520
rect 248052 176656 248104 176662
rect 248052 176598 248104 176604
rect 246304 175976 246356 175982
rect 246304 175918 246356 175924
rect 248064 175817 248092 176598
rect 248050 175808 248106 175817
rect 248050 175743 248106 175752
rect 249076 172802 249104 178774
rect 249248 177404 249300 177410
rect 249248 177346 249300 177352
rect 249156 176656 249208 176662
rect 249156 176598 249208 176604
rect 249168 174729 249196 176598
rect 249260 175273 249288 177346
rect 249246 175264 249302 175273
rect 249246 175199 249302 175208
rect 249154 174720 249210 174729
rect 249154 174655 249210 174664
rect 249154 172816 249210 172825
rect 249076 172774 249154 172802
rect 249154 172751 249210 172760
rect 249812 171873 249840 270506
rect 252560 229832 252612 229838
rect 252560 229774 252612 229780
rect 251180 214668 251232 214674
rect 251180 214610 251232 214616
rect 249892 210452 249944 210458
rect 249892 210394 249944 210400
rect 249798 171864 249854 171873
rect 249798 171799 249854 171808
rect 214746 161800 214802 161809
rect 214746 161735 214802 161744
rect 249904 161474 249932 210394
rect 249984 199572 250036 199578
rect 249984 199514 250036 199520
rect 249812 161446 249932 161474
rect 249812 155417 249840 161446
rect 249798 155408 249854 155417
rect 249798 155343 249854 155352
rect 215942 153776 215998 153785
rect 215942 153711 215998 153720
rect 214654 150512 214710 150521
rect 214654 150447 214710 150456
rect 214562 148472 214618 148481
rect 214562 148407 214618 148416
rect 213918 147928 213974 147937
rect 213918 147863 213974 147872
rect 213932 147694 213960 147863
rect 213920 147688 213972 147694
rect 213920 147630 213972 147636
rect 214010 147248 214066 147257
rect 214010 147183 214066 147192
rect 213918 146568 213974 146577
rect 213918 146503 213974 146512
rect 213932 146402 213960 146503
rect 213920 146396 213972 146402
rect 213920 146338 213972 146344
rect 214024 146334 214052 147183
rect 214012 146328 214064 146334
rect 214012 146270 214064 146276
rect 214010 145888 214066 145897
rect 214010 145823 214066 145832
rect 213918 145208 213974 145217
rect 213918 145143 213974 145152
rect 213932 144974 213960 145143
rect 214024 145042 214052 145823
rect 214012 145036 214064 145042
rect 214012 144978 214064 144984
rect 213920 144968 213972 144974
rect 213920 144910 213972 144916
rect 214010 144528 214066 144537
rect 214010 144463 214066 144472
rect 213918 143848 213974 143857
rect 213918 143783 213974 143792
rect 213932 143614 213960 143783
rect 214024 143682 214052 144463
rect 214012 143676 214064 143682
rect 214012 143618 214064 143624
rect 213920 143608 213972 143614
rect 213920 143550 213972 143556
rect 214010 143304 214066 143313
rect 214010 143239 214066 143248
rect 213918 142624 213974 142633
rect 213918 142559 213974 142568
rect 213932 142254 213960 142559
rect 213920 142248 213972 142254
rect 213920 142190 213972 142196
rect 214024 142186 214052 143239
rect 214012 142180 214064 142186
rect 214668 142154 214696 150447
rect 214012 142122 214064 142128
rect 214576 142126 214696 142154
rect 213918 141944 213974 141953
rect 213918 141879 213974 141888
rect 213932 140826 213960 141879
rect 213920 140820 213972 140826
rect 213920 140762 213972 140768
rect 213918 140584 213974 140593
rect 213918 140519 213974 140528
rect 213932 139466 213960 140519
rect 213920 139460 213972 139466
rect 213920 139402 213972 139408
rect 213918 138680 213974 138689
rect 213918 138615 213974 138624
rect 213932 138038 213960 138615
rect 213920 138032 213972 138038
rect 213920 137974 213972 137980
rect 214102 138000 214158 138009
rect 214102 137935 214158 137944
rect 213918 137320 213974 137329
rect 213918 137255 213974 137264
rect 213932 136678 213960 137255
rect 213920 136672 213972 136678
rect 213920 136614 213972 136620
rect 214010 136640 214066 136649
rect 214010 136575 214066 136584
rect 214024 135386 214052 136575
rect 214012 135380 214064 135386
rect 214012 135322 214064 135328
rect 213920 135312 213972 135318
rect 213918 135280 213920 135289
rect 213972 135280 213974 135289
rect 213918 135215 213974 135224
rect 214010 134600 214066 134609
rect 214010 134535 214066 134544
rect 213920 134020 213972 134026
rect 213920 133962 213972 133968
rect 213932 133929 213960 133962
rect 214024 133958 214052 134535
rect 214012 133952 214064 133958
rect 213918 133920 213974 133929
rect 214012 133894 214064 133900
rect 213918 133855 213974 133864
rect 213918 133376 213974 133385
rect 213918 133311 213974 133320
rect 213932 132938 213960 133311
rect 214116 133210 214144 137935
rect 214576 137290 214604 142126
rect 214654 139224 214710 139233
rect 214654 139159 214710 139168
rect 214564 137284 214616 137290
rect 214564 137226 214616 137232
rect 214104 133204 214156 133210
rect 214104 133146 214156 133152
rect 213920 132932 213972 132938
rect 213920 132874 213972 132880
rect 213918 132016 213974 132025
rect 213918 131951 213974 131960
rect 213932 131170 213960 131951
rect 213920 131164 213972 131170
rect 213920 131106 213972 131112
rect 213918 130656 213974 130665
rect 213918 130591 213974 130600
rect 213932 129810 213960 130591
rect 213920 129804 213972 129810
rect 213920 129746 213972 129752
rect 214010 129296 214066 129305
rect 214010 129231 214066 129240
rect 213918 128752 213974 128761
rect 213918 128687 213974 128696
rect 213932 128382 213960 128687
rect 214024 128450 214052 129231
rect 214012 128444 214064 128450
rect 214012 128386 214064 128392
rect 213920 128376 213972 128382
rect 213920 128318 213972 128324
rect 214010 128072 214066 128081
rect 214010 128007 214066 128016
rect 213918 127392 213974 127401
rect 213918 127327 213974 127336
rect 213932 127090 213960 127327
rect 213920 127084 213972 127090
rect 213920 127026 213972 127032
rect 214024 127022 214052 128007
rect 214012 127016 214064 127022
rect 214012 126958 214064 126964
rect 214010 126712 214066 126721
rect 214010 126647 214066 126656
rect 213918 126032 213974 126041
rect 213918 125967 213974 125976
rect 213932 125662 213960 125967
rect 214024 125730 214052 126647
rect 214012 125724 214064 125730
rect 214012 125666 214064 125672
rect 213920 125656 213972 125662
rect 213920 125598 213972 125604
rect 214010 125352 214066 125361
rect 214010 125287 214066 125296
rect 213918 124672 213974 124681
rect 213918 124607 213974 124616
rect 213932 124302 213960 124607
rect 213920 124296 213972 124302
rect 213920 124238 213972 124244
rect 214024 124234 214052 125287
rect 214012 124228 214064 124234
rect 214012 124170 214064 124176
rect 214010 124128 214066 124137
rect 214010 124063 214066 124072
rect 213918 123448 213974 123457
rect 214024 123418 214052 124063
rect 213918 123383 213974 123392
rect 214012 123412 214064 123418
rect 213932 122874 213960 123383
rect 214012 123354 214064 123360
rect 213920 122868 213972 122874
rect 214668 122834 214696 139159
rect 213920 122810 213972 122816
rect 214576 122806 214696 122834
rect 214010 122768 214066 122777
rect 214010 122703 214066 122712
rect 213918 122088 213974 122097
rect 213918 122023 213974 122032
rect 213932 121514 213960 122023
rect 214024 121582 214052 122703
rect 214012 121576 214064 121582
rect 214012 121518 214064 121524
rect 213920 121508 213972 121514
rect 213920 121450 213972 121456
rect 214010 121408 214066 121417
rect 214010 121343 214066 121352
rect 213918 120728 213974 120737
rect 213918 120663 213974 120672
rect 213932 120154 213960 120663
rect 214024 120222 214052 121343
rect 214012 120216 214064 120222
rect 214012 120158 214064 120164
rect 213920 120148 213972 120154
rect 213920 120090 213972 120096
rect 214010 120048 214066 120057
rect 214010 119983 214066 119992
rect 213918 118824 213974 118833
rect 214024 118794 214052 119983
rect 214102 119504 214158 119513
rect 214102 119439 214158 119448
rect 214116 118862 214144 119439
rect 214104 118856 214156 118862
rect 214104 118798 214156 118804
rect 213918 118759 213974 118768
rect 214012 118788 214064 118794
rect 213932 118726 213960 118759
rect 214012 118730 214064 118736
rect 213920 118720 213972 118726
rect 213920 118662 213972 118668
rect 213918 118144 213974 118153
rect 213918 118079 213974 118088
rect 213276 117972 213328 117978
rect 213276 117914 213328 117920
rect 213182 117464 213238 117473
rect 213182 117399 213238 117408
rect 211988 114640 212040 114646
rect 211988 114582 212040 114588
rect 211894 91624 211950 91633
rect 211894 91559 211950 91568
rect 212000 84114 212028 114582
rect 212080 104984 212132 104990
rect 212080 104926 212132 104932
rect 212092 89690 212120 104926
rect 212080 89684 212132 89690
rect 212080 89626 212132 89632
rect 211988 84108 212040 84114
rect 211988 84050 212040 84056
rect 213196 82686 213224 117399
rect 213932 117366 213960 118079
rect 213920 117360 213972 117366
rect 213920 117302 213972 117308
rect 214010 116784 214066 116793
rect 214010 116719 214066 116728
rect 213918 116104 213974 116113
rect 213918 116039 213920 116048
rect 213972 116039 213974 116048
rect 213920 116010 213972 116016
rect 214024 116006 214052 116719
rect 214012 116000 214064 116006
rect 214012 115942 214064 115948
rect 214010 115424 214066 115433
rect 214010 115359 214066 115368
rect 213918 114880 213974 114889
rect 213918 114815 213974 114824
rect 213932 114578 213960 114815
rect 214024 114646 214052 115359
rect 214012 114640 214064 114646
rect 214012 114582 214064 114588
rect 213920 114572 213972 114578
rect 213920 114514 213972 114520
rect 214010 114200 214066 114209
rect 214010 114135 214066 114144
rect 213918 113520 213974 113529
rect 213918 113455 213974 113464
rect 213932 113218 213960 113455
rect 214024 113286 214052 114135
rect 214012 113280 214064 113286
rect 214012 113222 214064 113228
rect 213920 113212 213972 113218
rect 213920 113154 213972 113160
rect 214010 112840 214066 112849
rect 214010 112775 214066 112784
rect 213918 112160 213974 112169
rect 213918 112095 213974 112104
rect 213932 111858 213960 112095
rect 214024 111926 214052 112775
rect 214012 111920 214064 111926
rect 214012 111862 214064 111868
rect 213920 111852 213972 111858
rect 213920 111794 213972 111800
rect 214010 111480 214066 111489
rect 214010 111415 214066 111424
rect 213918 110800 213974 110809
rect 213918 110735 213974 110744
rect 213932 110566 213960 110735
rect 213920 110560 213972 110566
rect 213920 110502 213972 110508
rect 214024 110498 214052 111415
rect 214012 110492 214064 110498
rect 214012 110434 214064 110440
rect 213918 110256 213974 110265
rect 213918 110191 213974 110200
rect 213932 109070 213960 110191
rect 213920 109064 213972 109070
rect 213920 109006 213972 109012
rect 214010 108896 214066 108905
rect 214010 108831 214066 108840
rect 213918 108216 213974 108225
rect 213918 108151 213974 108160
rect 213932 107710 213960 108151
rect 214024 107778 214052 108831
rect 214012 107772 214064 107778
rect 214012 107714 214064 107720
rect 213920 107704 213972 107710
rect 213920 107646 213972 107652
rect 213918 107536 213974 107545
rect 213918 107471 213974 107480
rect 213932 106350 213960 107471
rect 213920 106344 213972 106350
rect 213920 106286 213972 106292
rect 214010 106176 214066 106185
rect 214010 106111 214066 106120
rect 213918 105632 213974 105641
rect 213918 105567 213974 105576
rect 213932 104922 213960 105567
rect 214024 104990 214052 106111
rect 214012 104984 214064 104990
rect 214012 104926 214064 104932
rect 213920 104916 213972 104922
rect 213920 104858 213972 104864
rect 213918 104272 213974 104281
rect 213918 104207 213974 104216
rect 213932 103562 213960 104207
rect 213920 103556 213972 103562
rect 213920 103498 213972 103504
rect 213918 102232 213974 102241
rect 213918 102167 213920 102176
rect 213972 102167 213974 102176
rect 213920 102138 213972 102144
rect 214010 101552 214066 101561
rect 214010 101487 214066 101496
rect 213918 101008 213974 101017
rect 213918 100943 213974 100952
rect 213932 100774 213960 100943
rect 214024 100842 214052 101487
rect 214012 100836 214064 100842
rect 214012 100778 214064 100784
rect 213920 100768 213972 100774
rect 213920 100710 213972 100716
rect 214010 100328 214066 100337
rect 214010 100263 214066 100272
rect 213918 99648 213974 99657
rect 213918 99583 213974 99592
rect 213932 99482 213960 99583
rect 213920 99476 213972 99482
rect 213920 99418 213972 99424
rect 214024 99414 214052 100263
rect 214012 99408 214064 99414
rect 214012 99350 214064 99356
rect 213918 98968 213974 98977
rect 213918 98903 213974 98912
rect 213932 98054 213960 98903
rect 213920 98048 213972 98054
rect 213920 97990 213972 97996
rect 213918 97608 213974 97617
rect 213918 97543 213974 97552
rect 213932 96694 213960 97543
rect 214576 97306 214604 122806
rect 214654 106856 214710 106865
rect 214654 106791 214710 106800
rect 214564 97300 214616 97306
rect 214564 97242 214616 97248
rect 213920 96688 213972 96694
rect 213920 96630 213972 96636
rect 214562 96384 214618 96393
rect 214562 96319 214618 96328
rect 214576 86970 214604 96319
rect 214564 86964 214616 86970
rect 214564 86906 214616 86912
rect 213184 82680 213236 82686
rect 213184 82622 213236 82628
rect 214668 81394 214696 106791
rect 214838 98288 214894 98297
rect 214838 98223 214894 98232
rect 214746 96928 214802 96937
rect 214746 96863 214802 96872
rect 214760 88330 214788 96863
rect 214852 93158 214880 98223
rect 214840 93152 214892 93158
rect 214840 93094 214892 93100
rect 215956 90914 215984 153711
rect 249996 150793 250024 199514
rect 250076 191208 250128 191214
rect 250076 191150 250128 191156
rect 250088 190454 250116 191150
rect 250088 190426 250208 190454
rect 250180 166705 250208 190426
rect 250166 166696 250222 166705
rect 250166 166631 250222 166640
rect 251192 159633 251220 214610
rect 251272 211880 251324 211886
rect 251272 211822 251324 211828
rect 251178 159624 251234 159633
rect 251178 159559 251234 159568
rect 251284 158817 251312 211822
rect 251456 181484 251508 181490
rect 251456 181426 251508 181432
rect 251364 165028 251416 165034
rect 251364 164970 251416 164976
rect 251376 164393 251404 164970
rect 251362 164384 251418 164393
rect 251362 164319 251418 164328
rect 251364 163124 251416 163130
rect 251364 163066 251416 163072
rect 251376 163033 251404 163066
rect 251362 163024 251418 163033
rect 251362 162959 251418 162968
rect 251468 161474 251496 181426
rect 251822 173360 251878 173369
rect 251822 173295 251878 173304
rect 251836 172718 251864 173295
rect 251824 172712 251876 172718
rect 251824 172654 251876 172660
rect 252008 172508 252060 172514
rect 252008 172450 252060 172456
rect 252020 171465 252048 172450
rect 252468 172440 252520 172446
rect 252466 172408 252468 172417
rect 252520 172408 252522 172417
rect 252466 172343 252522 172352
rect 252006 171456 252062 171465
rect 252006 171391 252062 171400
rect 252100 171080 252152 171086
rect 252100 171022 252152 171028
rect 251822 170504 251878 170513
rect 251822 170439 251878 170448
rect 251836 169998 251864 170439
rect 252112 170105 252140 171022
rect 252468 170944 252520 170950
rect 252466 170912 252468 170921
rect 252520 170912 252522 170921
rect 252466 170847 252522 170856
rect 252098 170096 252154 170105
rect 252098 170031 252154 170040
rect 251824 169992 251876 169998
rect 251824 169934 251876 169940
rect 252008 169244 252060 169250
rect 252008 169186 252060 169192
rect 252020 168609 252048 169186
rect 252466 169144 252522 169153
rect 252466 169079 252522 169088
rect 252006 168600 252062 168609
rect 252006 168535 252062 168544
rect 252480 168502 252508 169079
rect 252468 168496 252520 168502
rect 252468 168438 252520 168444
rect 252100 168360 252152 168366
rect 252100 168302 252152 168308
rect 251916 168224 251968 168230
rect 251914 168192 251916 168201
rect 251968 168192 251970 168201
rect 251914 168127 251970 168136
rect 252112 167249 252140 168302
rect 252468 168088 252520 168094
rect 252468 168030 252520 168036
rect 252480 167657 252508 168030
rect 252466 167648 252522 167657
rect 252466 167583 252522 167592
rect 252098 167240 252154 167249
rect 252098 167175 252154 167184
rect 251824 166932 251876 166938
rect 251824 166874 251876 166880
rect 251836 166297 251864 166874
rect 251822 166288 251878 166297
rect 251822 166223 251878 166232
rect 252468 165504 252520 165510
rect 252468 165446 252520 165452
rect 252376 165436 252428 165442
rect 252376 165378 252428 165384
rect 252388 164801 252416 165378
rect 252480 165345 252508 165446
rect 252466 165336 252522 165345
rect 252466 165271 252522 165280
rect 252374 164792 252430 164801
rect 252374 164727 252430 164736
rect 252468 164212 252520 164218
rect 252468 164154 252520 164160
rect 252480 163985 252508 164154
rect 252466 163976 252522 163985
rect 252466 163911 252522 163920
rect 252468 162852 252520 162858
rect 252468 162794 252520 162800
rect 252100 162784 252152 162790
rect 252100 162726 252152 162732
rect 252112 161537 252140 162726
rect 252480 162489 252508 162794
rect 252466 162480 252522 162489
rect 252466 162415 252522 162424
rect 251376 161446 251496 161474
rect 252098 161528 252154 161537
rect 252098 161463 252154 161472
rect 251270 158808 251326 158817
rect 251270 158743 251326 158752
rect 251180 154148 251232 154154
rect 251180 154090 251232 154096
rect 250442 152960 250498 152969
rect 250442 152895 250498 152904
rect 249982 150784 250038 150793
rect 249982 150719 250038 150728
rect 249890 138952 249946 138961
rect 249890 138887 249946 138896
rect 249904 138145 249932 138887
rect 249890 138136 249946 138145
rect 249890 138071 249946 138080
rect 250456 136649 250484 152895
rect 251192 152153 251220 154090
rect 251178 152144 251234 152153
rect 251178 152079 251234 152088
rect 251272 151496 251324 151502
rect 251272 151438 251324 151444
rect 251284 151201 251312 151438
rect 251270 151192 251326 151201
rect 251270 151127 251326 151136
rect 251272 148912 251324 148918
rect 251270 148880 251272 148889
rect 251324 148880 251326 148889
rect 251270 148815 251326 148824
rect 251376 142154 251404 161446
rect 252468 161424 252520 161430
rect 252468 161366 252520 161372
rect 252098 161120 252154 161129
rect 252098 161055 252154 161064
rect 252008 160880 252060 160886
rect 252008 160822 252060 160828
rect 252020 160177 252048 160822
rect 252112 160342 252140 161055
rect 252480 160585 252508 161366
rect 252466 160576 252522 160585
rect 252466 160511 252522 160520
rect 252100 160336 252152 160342
rect 252100 160278 252152 160284
rect 252006 160168 252062 160177
rect 252006 160103 252062 160112
rect 252468 160064 252520 160070
rect 252468 160006 252520 160012
rect 252480 159225 252508 160006
rect 252466 159216 252522 159225
rect 252466 159151 252522 159160
rect 252376 158704 252428 158710
rect 252376 158646 252428 158652
rect 252388 157865 252416 158646
rect 252468 158636 252520 158642
rect 252468 158578 252520 158584
rect 252480 158273 252508 158578
rect 252466 158264 252522 158273
rect 252466 158199 252522 158208
rect 252374 157856 252430 157865
rect 252374 157791 252430 157800
rect 252376 157344 252428 157350
rect 252376 157286 252428 157292
rect 252466 157312 252522 157321
rect 252388 156913 252416 157286
rect 252466 157247 252468 157256
rect 252520 157247 252522 157256
rect 252468 157218 252520 157224
rect 252374 156904 252430 156913
rect 252374 156839 252430 156848
rect 252466 155952 252522 155961
rect 252376 155916 252428 155922
rect 252466 155887 252522 155896
rect 252376 155858 252428 155864
rect 252388 155009 252416 155858
rect 252480 155854 252508 155887
rect 252468 155848 252520 155854
rect 252468 155790 252520 155796
rect 252374 155000 252430 155009
rect 252374 154935 252430 154944
rect 252376 154488 252428 154494
rect 252572 154465 252600 229774
rect 252652 221468 252704 221474
rect 252652 221410 252704 221416
rect 252664 169561 252692 221410
rect 252744 205012 252796 205018
rect 252744 204954 252796 204960
rect 252650 169552 252706 169561
rect 252650 169487 252706 169496
rect 252756 165753 252784 204954
rect 252836 192568 252888 192574
rect 252836 192510 252888 192516
rect 252742 165744 252798 165753
rect 252742 165679 252798 165688
rect 252848 165034 252876 192510
rect 252836 165028 252888 165034
rect 252836 164970 252888 164976
rect 253204 157412 253256 157418
rect 253204 157354 253256 157360
rect 252376 154430 252428 154436
rect 252558 154456 252614 154465
rect 252388 153513 252416 154430
rect 252468 154420 252520 154426
rect 252558 154391 252614 154400
rect 252468 154362 252520 154368
rect 252480 154057 252508 154362
rect 252466 154048 252522 154057
rect 252466 153983 252522 153992
rect 252374 153504 252430 153513
rect 252374 153439 252430 153448
rect 252468 153196 252520 153202
rect 252468 153138 252520 153144
rect 252480 153105 252508 153138
rect 252466 153096 252522 153105
rect 252466 153031 252522 153040
rect 252468 151768 252520 151774
rect 252466 151736 252468 151745
rect 252520 151736 252522 151745
rect 252466 151671 252522 151680
rect 252284 150408 252336 150414
rect 252284 150350 252336 150356
rect 252296 149841 252324 150350
rect 252282 149832 252338 149841
rect 252282 149767 252338 149776
rect 251732 149320 251784 149326
rect 251730 149288 251732 149297
rect 251784 149288 251786 149297
rect 251730 149223 251786 149232
rect 252468 149048 252520 149054
rect 252468 148990 252520 148996
rect 251916 148776 251968 148782
rect 251916 148718 251968 148724
rect 251928 148345 251956 148718
rect 251914 148336 251970 148345
rect 251914 148271 251970 148280
rect 252480 147937 252508 148990
rect 252466 147928 252522 147937
rect 252466 147863 252522 147872
rect 252468 147620 252520 147626
rect 252468 147562 252520 147568
rect 251732 147552 251784 147558
rect 252480 147529 252508 147562
rect 251732 147494 251784 147500
rect 252466 147520 252522 147529
rect 251744 146985 251772 147494
rect 252466 147455 252522 147464
rect 251730 146976 251786 146985
rect 251730 146911 251786 146920
rect 251732 146872 251784 146878
rect 251732 146814 251784 146820
rect 251744 146577 251772 146814
rect 251730 146568 251786 146577
rect 251730 146503 251786 146512
rect 251916 146260 251968 146266
rect 251916 146202 251968 146208
rect 251732 146192 251784 146198
rect 251732 146134 251784 146140
rect 251744 145625 251772 146134
rect 251928 146033 251956 146202
rect 252100 146124 252152 146130
rect 252100 146066 252152 146072
rect 251914 146024 251970 146033
rect 251914 145959 251970 145968
rect 251730 145616 251786 145625
rect 251730 145551 251786 145560
rect 252112 145081 252140 146066
rect 252098 145072 252154 145081
rect 252098 145007 252154 145016
rect 252376 144900 252428 144906
rect 252376 144842 252428 144848
rect 252100 144220 252152 144226
rect 252100 144162 252152 144168
rect 251916 142860 251968 142866
rect 251916 142802 251968 142808
rect 251284 142126 251404 142154
rect 251284 140865 251312 142126
rect 251824 141432 251876 141438
rect 251824 141374 251876 141380
rect 251270 140856 251326 140865
rect 251270 140791 251326 140800
rect 251364 139936 251416 139942
rect 251362 139904 251364 139913
rect 251416 139904 251418 139913
rect 251362 139839 251418 139848
rect 251548 138712 251600 138718
rect 251548 138654 251600 138660
rect 251362 138000 251418 138009
rect 251362 137935 251418 137944
rect 251376 137902 251404 137935
rect 251364 137896 251416 137902
rect 251364 137838 251416 137844
rect 250442 136640 250498 136649
rect 250442 136575 250498 136584
rect 251560 136241 251588 138654
rect 251546 136232 251602 136241
rect 251546 136167 251602 136176
rect 251640 135244 251692 135250
rect 251640 135186 251692 135192
rect 251652 134745 251680 135186
rect 251638 134736 251694 134745
rect 251638 134671 251694 134680
rect 251548 134564 251600 134570
rect 251548 134506 251600 134512
rect 251456 133884 251508 133890
rect 251456 133826 251508 133832
rect 251468 133385 251496 133826
rect 251454 133376 251510 133385
rect 251454 133311 251510 133320
rect 251362 132424 251418 132433
rect 251362 132359 251418 132368
rect 251376 132326 251404 132359
rect 251364 132320 251416 132326
rect 251364 132262 251416 132268
rect 251560 127673 251588 134506
rect 251732 131096 251784 131102
rect 251732 131038 251784 131044
rect 251744 130529 251772 131038
rect 251730 130520 251786 130529
rect 251730 130455 251786 130464
rect 251732 129736 251784 129742
rect 251732 129678 251784 129684
rect 251744 129169 251772 129678
rect 251730 129160 251786 129169
rect 251730 129095 251786 129104
rect 251546 127664 251602 127673
rect 251546 127599 251602 127608
rect 251272 126268 251324 126274
rect 251272 126210 251324 126216
rect 251284 124409 251312 126210
rect 251270 124400 251326 124409
rect 251270 124335 251326 124344
rect 251364 120012 251416 120018
rect 251364 119954 251416 119960
rect 251376 119649 251404 119954
rect 251362 119640 251418 119649
rect 251362 119575 251418 119584
rect 251836 119241 251864 141374
rect 251928 126313 251956 142802
rect 252008 132388 252060 132394
rect 252008 132330 252060 132336
rect 252020 131481 252048 132330
rect 252006 131472 252062 131481
rect 252006 131407 252062 131416
rect 252008 131028 252060 131034
rect 252008 130970 252060 130976
rect 252020 130121 252048 130970
rect 252006 130112 252062 130121
rect 252006 130047 252062 130056
rect 252112 129826 252140 144162
rect 252388 144129 252416 144842
rect 252468 144832 252520 144838
rect 252468 144774 252520 144780
rect 252480 144673 252508 144774
rect 252466 144664 252522 144673
rect 252466 144599 252522 144608
rect 252374 144120 252430 144129
rect 252374 144055 252430 144064
rect 252468 144084 252520 144090
rect 252468 144026 252520 144032
rect 252480 143721 252508 144026
rect 252466 143712 252522 143721
rect 252466 143647 252522 143656
rect 252468 143540 252520 143546
rect 252468 143482 252520 143488
rect 252480 143177 252508 143482
rect 252466 143168 252522 143177
rect 252466 143103 252522 143112
rect 252468 142112 252520 142118
rect 252468 142054 252520 142060
rect 252480 141409 252508 142054
rect 252466 141400 252522 141409
rect 252466 141335 252522 141344
rect 252468 139392 252520 139398
rect 252468 139334 252520 139340
rect 252480 138553 252508 139334
rect 252466 138544 252522 138553
rect 252466 138479 252522 138488
rect 252468 137964 252520 137970
rect 252468 137906 252520 137912
rect 252480 137057 252508 137906
rect 252466 137048 252522 137057
rect 252466 136983 252522 136992
rect 252468 136604 252520 136610
rect 252468 136546 252520 136552
rect 252376 136536 252428 136542
rect 252376 136478 252428 136484
rect 252388 135289 252416 136478
rect 252480 135697 252508 136546
rect 252466 135688 252522 135697
rect 252466 135623 252522 135632
rect 252374 135280 252430 135289
rect 252374 135215 252430 135224
rect 252468 134632 252520 134638
rect 252468 134574 252520 134580
rect 252480 134337 252508 134574
rect 252466 134328 252522 134337
rect 252466 134263 252522 134272
rect 252468 133816 252520 133822
rect 252468 133758 252520 133764
rect 252480 132841 252508 133758
rect 252466 132832 252522 132841
rect 252466 132767 252522 132776
rect 252284 132456 252336 132462
rect 252284 132398 252336 132404
rect 252296 131889 252324 132398
rect 252282 131880 252338 131889
rect 252282 131815 252338 131824
rect 252466 130928 252522 130937
rect 252466 130863 252522 130872
rect 252480 129946 252508 130863
rect 252468 129940 252520 129946
rect 252468 129882 252520 129888
rect 252020 129798 252140 129826
rect 252020 129577 252048 129798
rect 252100 129668 252152 129674
rect 252100 129610 252152 129616
rect 252006 129568 252062 129577
rect 252006 129503 252062 129512
rect 252112 128625 252140 129610
rect 252098 128616 252154 128625
rect 252098 128551 252154 128560
rect 252008 128308 252060 128314
rect 252008 128250 252060 128256
rect 252020 127265 252048 128250
rect 252468 128240 252520 128246
rect 252466 128208 252468 128217
rect 252520 128208 252522 128217
rect 252466 128143 252522 128152
rect 252006 127256 252062 127265
rect 252006 127191 252062 127200
rect 252100 126948 252152 126954
rect 252100 126890 252152 126896
rect 251914 126304 251970 126313
rect 251914 126239 251970 126248
rect 252112 125769 252140 126890
rect 252468 126880 252520 126886
rect 252468 126822 252520 126828
rect 252480 126721 252508 126822
rect 252466 126712 252522 126721
rect 252466 126647 252522 126656
rect 252098 125760 252154 125769
rect 252098 125695 252154 125704
rect 252468 125588 252520 125594
rect 252468 125530 252520 125536
rect 252376 125520 252428 125526
rect 252376 125462 252428 125468
rect 252284 124908 252336 124914
rect 252284 124850 252336 124856
rect 252008 124092 252060 124098
rect 252008 124034 252060 124040
rect 252020 123049 252048 124034
rect 252296 124001 252324 124850
rect 252388 124817 252416 125462
rect 252480 125361 252508 125530
rect 252466 125352 252522 125361
rect 252466 125287 252522 125296
rect 252374 124808 252430 124817
rect 252374 124743 252430 124752
rect 252468 124160 252520 124166
rect 252468 124102 252520 124108
rect 252282 123992 252338 124001
rect 252282 123927 252338 123936
rect 252100 123480 252152 123486
rect 252480 123457 252508 124102
rect 252100 123422 252152 123428
rect 252466 123448 252522 123457
rect 252006 123040 252062 123049
rect 252006 122975 252062 122984
rect 252112 122834 252140 123422
rect 252466 123383 252522 123392
rect 252020 122806 252140 122834
rect 251916 121440 251968 121446
rect 251916 121382 251968 121388
rect 251928 120193 251956 121382
rect 251914 120184 251970 120193
rect 251914 120119 251970 120128
rect 251822 119232 251878 119241
rect 251822 119167 251878 119176
rect 251180 118788 251232 118794
rect 251180 118730 251232 118736
rect 251192 117337 251220 118730
rect 251824 118652 251876 118658
rect 251824 118594 251876 118600
rect 251640 117972 251692 117978
rect 251640 117914 251692 117920
rect 251178 117328 251234 117337
rect 251178 117263 251234 117272
rect 251652 114481 251680 117914
rect 251836 117881 251864 118594
rect 251822 117872 251878 117881
rect 251822 117807 251878 117816
rect 251916 117292 251968 117298
rect 251916 117234 251968 117240
rect 251928 116385 251956 117234
rect 251914 116376 251970 116385
rect 251914 116311 251970 116320
rect 251638 114472 251694 114481
rect 251638 114407 251694 114416
rect 252020 112713 252048 122806
rect 252468 122800 252520 122806
rect 252468 122742 252520 122748
rect 252376 122732 252428 122738
rect 252376 122674 252428 122680
rect 252388 122097 252416 122674
rect 252480 122505 252508 122742
rect 252466 122496 252522 122505
rect 252466 122431 252522 122440
rect 252374 122088 252430 122097
rect 252374 122023 252430 122032
rect 252468 122052 252520 122058
rect 252468 121994 252520 122000
rect 252480 121553 252508 121994
rect 252466 121544 252522 121553
rect 252466 121479 252522 121488
rect 252468 121372 252520 121378
rect 252468 121314 252520 121320
rect 252376 121304 252428 121310
rect 252376 121246 252428 121252
rect 252388 120601 252416 121246
rect 252480 121145 252508 121314
rect 252466 121136 252522 121145
rect 252466 121071 252522 121080
rect 252374 120592 252430 120601
rect 252374 120527 252430 120536
rect 252468 120080 252520 120086
rect 252468 120022 252520 120028
rect 252480 118833 252508 120022
rect 252466 118824 252522 118833
rect 253216 118794 253244 157354
rect 253952 154154 253980 274654
rect 254032 262880 254084 262886
rect 254032 262822 254084 262828
rect 254044 163130 254072 262822
rect 254124 220244 254176 220250
rect 254124 220186 254176 220192
rect 254032 163124 254084 163130
rect 254032 163066 254084 163072
rect 253940 154148 253992 154154
rect 253940 154090 253992 154096
rect 254136 148918 254164 220186
rect 254216 200932 254268 200938
rect 254216 200874 254268 200880
rect 254228 151502 254256 200874
rect 255332 168230 255360 294170
rect 263600 292800 263652 292806
rect 263600 292742 263652 292748
rect 255412 267028 255464 267034
rect 255412 266970 255464 266976
rect 255320 168224 255372 168230
rect 255320 168166 255372 168172
rect 255424 160886 255452 266970
rect 262220 217456 262272 217462
rect 262220 217398 262272 217404
rect 260840 200864 260892 200870
rect 260840 200806 260892 200812
rect 258172 199436 258224 199442
rect 258172 199378 258224 199384
rect 256700 191276 256752 191282
rect 256700 191218 256752 191224
rect 255504 185768 255556 185774
rect 255504 185710 255556 185716
rect 255412 160880 255464 160886
rect 255412 160822 255464 160828
rect 254676 153264 254728 153270
rect 254676 153206 254728 153212
rect 254216 151496 254268 151502
rect 254216 151438 254268 151444
rect 254124 148912 254176 148918
rect 254124 148854 254176 148860
rect 253480 144968 253532 144974
rect 253480 144910 253532 144916
rect 253386 142760 253442 142769
rect 253386 142695 253442 142704
rect 253400 142361 253428 142695
rect 253386 142352 253442 142361
rect 253386 142287 253442 142296
rect 253388 140072 253440 140078
rect 253388 140014 253440 140020
rect 253296 137284 253348 137290
rect 253296 137226 253348 137232
rect 252466 118759 252522 118768
rect 253204 118788 253256 118794
rect 253204 118730 253256 118736
rect 252468 118584 252520 118590
rect 252468 118526 252520 118532
rect 252480 118289 252508 118526
rect 252466 118280 252522 118289
rect 252466 118215 252522 118224
rect 252376 117224 252428 117230
rect 252376 117166 252428 117172
rect 252388 115977 252416 117166
rect 252468 117156 252520 117162
rect 252468 117098 252520 117104
rect 252480 116929 252508 117098
rect 252466 116920 252522 116929
rect 252466 116855 252522 116864
rect 252374 115968 252430 115977
rect 252374 115903 252430 115912
rect 252468 115932 252520 115938
rect 252468 115874 252520 115880
rect 252376 115864 252428 115870
rect 252376 115806 252428 115812
rect 252388 115025 252416 115806
rect 252480 115433 252508 115874
rect 252466 115424 252522 115433
rect 252466 115359 252522 115368
rect 252374 115016 252430 115025
rect 252374 114951 252430 114960
rect 252468 114504 252520 114510
rect 252468 114446 252520 114452
rect 252376 114436 252428 114442
rect 252376 114378 252428 114384
rect 252100 113756 252152 113762
rect 252100 113698 252152 113704
rect 252112 113121 252140 113698
rect 252388 113529 252416 114378
rect 252480 114073 252508 114446
rect 252466 114064 252522 114073
rect 252466 113999 252522 114008
rect 252374 113520 252430 113529
rect 252374 113455 252430 113464
rect 252468 113144 252520 113150
rect 252098 113112 252154 113121
rect 252468 113086 252520 113092
rect 252098 113047 252154 113056
rect 252006 112704 252062 112713
rect 252006 112639 252062 112648
rect 252376 112464 252428 112470
rect 252376 112406 252428 112412
rect 251548 111852 251600 111858
rect 251548 111794 251600 111800
rect 251560 110809 251588 111794
rect 252282 111752 252338 111761
rect 252282 111687 252284 111696
rect 252336 111687 252338 111696
rect 252284 111658 252336 111664
rect 251732 111104 251784 111110
rect 251732 111046 251784 111052
rect 251546 110800 251602 110809
rect 251546 110735 251602 110744
rect 251272 110356 251324 110362
rect 251272 110298 251324 110304
rect 251180 107908 251232 107914
rect 251180 107850 251232 107856
rect 251192 103737 251220 107850
rect 251284 107545 251312 110298
rect 251364 108996 251416 109002
rect 251364 108938 251416 108944
rect 251376 107953 251404 108938
rect 251744 108361 251772 111046
rect 252388 109857 252416 112406
rect 252480 112169 252508 113086
rect 252466 112160 252522 112169
rect 252466 112095 252522 112104
rect 252468 111784 252520 111790
rect 252468 111726 252520 111732
rect 252480 111217 252508 111726
rect 252466 111208 252522 111217
rect 252466 111143 252522 111152
rect 252468 110424 252520 110430
rect 252468 110366 252520 110372
rect 252480 110265 252508 110366
rect 252466 110256 252522 110265
rect 252466 110191 252522 110200
rect 252374 109848 252430 109857
rect 252374 109783 252430 109792
rect 251916 109336 251968 109342
rect 251914 109304 251916 109313
rect 251968 109304 251970 109313
rect 251914 109239 251970 109248
rect 252468 108928 252520 108934
rect 252466 108896 252468 108905
rect 252520 108896 252522 108905
rect 252466 108831 252522 108840
rect 251730 108352 251786 108361
rect 251730 108287 251786 108296
rect 251362 107944 251418 107953
rect 251362 107879 251418 107888
rect 251364 107636 251416 107642
rect 251364 107578 251416 107584
rect 251270 107536 251326 107545
rect 251270 107471 251326 107480
rect 251376 106593 251404 107578
rect 252468 107568 252520 107574
rect 252468 107510 252520 107516
rect 252480 107001 252508 107510
rect 252466 106992 252522 107001
rect 252466 106927 252522 106936
rect 251362 106584 251418 106593
rect 251362 106519 251418 106528
rect 252008 106276 252060 106282
rect 252008 106218 252060 106224
rect 252020 106049 252048 106218
rect 252284 106208 252336 106214
rect 252284 106150 252336 106156
rect 252006 106040 252062 106049
rect 252006 105975 252062 105984
rect 252296 105641 252324 106150
rect 252282 105632 252338 105641
rect 252008 105596 252060 105602
rect 252282 105567 252338 105576
rect 252008 105538 252060 105544
rect 252020 104689 252048 105538
rect 252468 104848 252520 104854
rect 252468 104790 252520 104796
rect 252006 104680 252062 104689
rect 252006 104615 252062 104624
rect 251548 104168 251600 104174
rect 252480 104145 252508 104790
rect 251548 104110 251600 104116
rect 252466 104136 252522 104145
rect 251178 103728 251234 103737
rect 251178 103663 251234 103672
rect 216034 102912 216090 102921
rect 216034 102847 216090 102856
rect 215944 90908 215996 90914
rect 215944 90850 215996 90856
rect 214748 88324 214800 88330
rect 214748 88266 214800 88272
rect 216048 84182 216076 102847
rect 251180 102808 251232 102814
rect 251178 102776 251180 102785
rect 251232 102776 251234 102785
rect 251178 102711 251234 102720
rect 251560 102241 251588 104110
rect 252466 104071 252522 104080
rect 253204 103692 253256 103698
rect 253204 103634 253256 103640
rect 252468 103488 252520 103494
rect 252468 103430 252520 103436
rect 252480 103193 252508 103430
rect 252466 103184 252522 103193
rect 252466 103119 252522 103128
rect 252100 102264 252152 102270
rect 251546 102232 251602 102241
rect 252100 102206 252152 102212
rect 251546 102167 251602 102176
rect 252112 100881 252140 102206
rect 252468 102128 252520 102134
rect 252468 102070 252520 102076
rect 252376 102060 252428 102066
rect 252376 102002 252428 102008
rect 252388 101425 252416 102002
rect 252480 101833 252508 102070
rect 252466 101824 252522 101833
rect 252466 101759 252522 101768
rect 252374 101416 252430 101425
rect 252374 101351 252430 101360
rect 252098 100872 252154 100881
rect 252098 100807 252154 100816
rect 252100 100700 252152 100706
rect 252100 100642 252152 100648
rect 251180 100156 251232 100162
rect 251180 100098 251232 100104
rect 251192 99929 251220 100098
rect 251178 99920 251234 99929
rect 251178 99855 251234 99864
rect 252112 99521 252140 100642
rect 252468 100632 252520 100638
rect 252468 100574 252520 100580
rect 252480 100473 252508 100574
rect 252466 100464 252522 100473
rect 252466 100399 252522 100408
rect 252098 99512 252154 99521
rect 252098 99447 252154 99456
rect 252192 99340 252244 99346
rect 252192 99282 252244 99288
rect 251180 98660 251232 98666
rect 251180 98602 251232 98608
rect 251192 98569 251220 98602
rect 251178 98560 251234 98569
rect 251178 98495 251234 98504
rect 252204 98025 252232 99282
rect 252284 99204 252336 99210
rect 252284 99146 252336 99152
rect 252296 98977 252324 99146
rect 252282 98968 252338 98977
rect 252282 98903 252338 98912
rect 252190 98016 252246 98025
rect 252190 97951 252246 97960
rect 252468 97912 252520 97918
rect 252468 97854 252520 97860
rect 252480 97617 252508 97854
rect 252466 97608 252522 97617
rect 249524 97572 249576 97578
rect 252466 97543 252522 97552
rect 249524 97514 249576 97520
rect 249536 96665 249564 97514
rect 251178 97064 251234 97073
rect 251178 96999 251234 97008
rect 249154 96656 249210 96665
rect 249154 96591 249210 96600
rect 249522 96656 249578 96665
rect 249522 96591 249578 96600
rect 248418 95704 248474 95713
rect 248418 95639 248474 95648
rect 248432 94518 248460 95639
rect 239404 94512 239456 94518
rect 239404 94454 239456 94460
rect 248420 94512 248472 94518
rect 248420 94454 248472 94460
rect 216036 84176 216088 84182
rect 216036 84118 216088 84124
rect 214656 81388 214708 81394
rect 214656 81330 214708 81336
rect 211804 78600 211856 78606
rect 211804 78542 211856 78548
rect 239416 4010 239444 94454
rect 249168 84194 249196 96591
rect 250444 95260 250496 95266
rect 250444 95202 250496 95208
rect 248432 84166 249196 84194
rect 248432 8294 248460 84166
rect 248420 8288 248472 8294
rect 248420 8230 248472 8236
rect 235816 4004 235868 4010
rect 235816 3946 235868 3952
rect 239404 4004 239456 4010
rect 239404 3946 239456 3952
rect 207664 3596 207716 3602
rect 207664 3538 207716 3544
rect 125874 3360 125930 3369
rect 125874 3295 125930 3304
rect 125888 480 125916 3295
rect 235828 480 235856 3946
rect 250456 2106 250484 95202
rect 251192 9654 251220 96999
rect 251180 9648 251232 9654
rect 251180 9590 251232 9596
rect 253216 3466 253244 103634
rect 253308 100162 253336 137226
rect 253400 102814 253428 140014
rect 253492 107914 253520 144910
rect 254584 140820 254636 140826
rect 254584 140762 254636 140768
rect 253480 107908 253532 107914
rect 253480 107850 253532 107856
rect 253388 102808 253440 102814
rect 253388 102750 253440 102756
rect 253296 100156 253348 100162
rect 253296 100098 253348 100104
rect 254596 98666 254624 140762
rect 254688 113762 254716 153206
rect 254768 151836 254820 151842
rect 254768 151778 254820 151784
rect 254676 113756 254728 113762
rect 254676 113698 254728 113704
rect 254780 111858 254808 151778
rect 255516 148782 255544 185710
rect 255596 176044 255648 176050
rect 255596 175986 255648 175992
rect 255504 148776 255556 148782
rect 255504 148718 255556 148724
rect 255608 146878 255636 175986
rect 256148 150476 256200 150482
rect 256148 150418 256200 150424
rect 256056 149728 256108 149734
rect 256056 149670 256108 149676
rect 255596 146872 255648 146878
rect 255596 146814 255648 146820
rect 255962 144120 256018 144129
rect 255962 144055 256018 144064
rect 254768 111852 254820 111858
rect 254768 111794 254820 111800
rect 254584 98660 254636 98666
rect 254584 98602 254636 98608
rect 255976 97578 256004 144055
rect 256068 99210 256096 149670
rect 256160 109342 256188 150418
rect 256240 146328 256292 146334
rect 256240 146270 256292 146276
rect 256148 109336 256200 109342
rect 256148 109278 256200 109284
rect 256252 106214 256280 146270
rect 256712 139942 256740 191218
rect 256792 187060 256844 187066
rect 256792 187002 256844 187008
rect 256804 149326 256832 187002
rect 258080 178900 258132 178906
rect 258080 178842 258132 178848
rect 256974 175944 257030 175953
rect 256974 175879 257030 175888
rect 256988 170950 257016 175879
rect 258092 172514 258120 178842
rect 258080 172508 258132 172514
rect 258080 172450 258132 172456
rect 258080 172372 258132 172378
rect 258080 172314 258132 172320
rect 256976 170944 257028 170950
rect 256976 170886 257028 170892
rect 258092 169250 258120 172314
rect 258184 169998 258212 199378
rect 259552 198076 259604 198082
rect 259552 198018 259604 198024
rect 259460 181620 259512 181626
rect 259460 181562 259512 181568
rect 258448 180328 258500 180334
rect 258448 180270 258500 180276
rect 258356 179104 258408 179110
rect 258356 179046 258408 179052
rect 258264 178968 258316 178974
rect 258264 178910 258316 178916
rect 258276 172378 258304 178910
rect 258264 172372 258316 172378
rect 258264 172314 258316 172320
rect 258264 172236 258316 172242
rect 258264 172178 258316 172184
rect 258172 169992 258224 169998
rect 258172 169934 258224 169940
rect 258080 169244 258132 169250
rect 258080 169186 258132 169192
rect 258276 160342 258304 172178
rect 258264 160336 258316 160342
rect 258264 160278 258316 160284
rect 257344 151904 257396 151910
rect 257344 151846 257396 151852
rect 256792 149320 256844 149326
rect 256792 149262 256844 149268
rect 256700 139936 256752 139942
rect 256700 139878 256752 139884
rect 257356 111722 257384 151846
rect 257528 147688 257580 147694
rect 257528 147630 257580 147636
rect 257436 142180 257488 142186
rect 257436 142122 257488 142128
rect 257344 111716 257396 111722
rect 257344 111658 257396 111664
rect 256240 106208 256292 106214
rect 256240 106150 256292 106156
rect 257448 102270 257476 142122
rect 257540 110362 257568 147630
rect 258368 142118 258396 179046
rect 258460 172242 258488 180270
rect 259472 172718 259500 181562
rect 259460 172712 259512 172718
rect 259460 172654 259512 172660
rect 258448 172236 258500 172242
rect 258448 172178 258500 172184
rect 258816 169788 258868 169794
rect 258816 169730 258868 169736
rect 258724 160132 258776 160138
rect 258724 160074 258776 160080
rect 258356 142112 258408 142118
rect 258356 142054 258408 142060
rect 258736 121310 258764 160074
rect 258828 129946 258856 169730
rect 259564 168502 259592 198018
rect 259644 181688 259696 181694
rect 259644 181630 259696 181636
rect 259552 168496 259604 168502
rect 259552 168438 259604 168444
rect 259656 168094 259684 181630
rect 259736 177608 259788 177614
rect 259736 177550 259788 177556
rect 259644 168088 259696 168094
rect 259644 168030 259696 168036
rect 258908 153876 258960 153882
rect 258908 153818 258960 153824
rect 258816 129940 258868 129946
rect 258816 129882 258868 129888
rect 258724 121304 258776 121310
rect 258724 121246 258776 121252
rect 258920 117162 258948 153818
rect 259748 144090 259776 177550
rect 260288 172576 260340 172582
rect 260288 172518 260340 172524
rect 260196 161492 260248 161498
rect 260196 161434 260248 161440
rect 260104 157480 260156 157486
rect 260104 157422 260156 157428
rect 259736 144084 259788 144090
rect 259736 144026 259788 144032
rect 260116 118590 260144 157422
rect 260208 122058 260236 161434
rect 260300 134638 260328 172518
rect 260852 166938 260880 200806
rect 260932 183184 260984 183190
rect 260932 183126 260984 183132
rect 260944 168366 260972 183126
rect 261116 183116 261168 183122
rect 261116 183058 261168 183064
rect 261024 177676 261076 177682
rect 261024 177618 261076 177624
rect 260932 168360 260984 168366
rect 260932 168302 260984 168308
rect 260840 166932 260892 166938
rect 260840 166874 260892 166880
rect 261036 165510 261064 177618
rect 261128 172446 261156 183058
rect 261116 172440 261168 172446
rect 261116 172382 261168 172388
rect 261760 171148 261812 171154
rect 261760 171090 261812 171096
rect 261668 165640 261720 165646
rect 261668 165582 261720 165588
rect 261024 165504 261076 165510
rect 261024 165446 261076 165452
rect 261576 162920 261628 162926
rect 261576 162862 261628 162868
rect 261484 155984 261536 155990
rect 261484 155926 261536 155932
rect 260288 134632 260340 134638
rect 260288 134574 260340 134580
rect 260196 122052 260248 122058
rect 260196 121994 260248 122000
rect 260104 118584 260156 118590
rect 260104 118526 260156 118532
rect 261496 117230 261524 155926
rect 261588 124098 261616 162862
rect 261680 126886 261708 165582
rect 261772 132326 261800 171090
rect 262232 171086 262260 217398
rect 262312 196716 262364 196722
rect 262312 196658 262364 196664
rect 262220 171080 262272 171086
rect 262220 171022 262272 171028
rect 262324 151774 262352 196658
rect 262496 175976 262548 175982
rect 262496 175918 262548 175924
rect 262508 160070 262536 175918
rect 262496 160064 262548 160070
rect 262496 160006 262548 160012
rect 262956 158772 263008 158778
rect 262956 158714 263008 158720
rect 262864 154624 262916 154630
rect 262864 154566 262916 154572
rect 262312 151768 262364 151774
rect 262312 151710 262364 151716
rect 261760 132320 261812 132326
rect 261760 132262 261812 132268
rect 261668 126880 261720 126886
rect 261668 126822 261720 126828
rect 261576 124092 261628 124098
rect 261576 124034 261628 124040
rect 261484 117224 261536 117230
rect 261484 117166 261536 117172
rect 258908 117156 258960 117162
rect 258908 117098 258960 117104
rect 262876 115870 262904 154566
rect 262968 120018 262996 158714
rect 263612 157282 263640 292742
rect 264256 235958 264284 699654
rect 269776 323610 269804 700334
rect 269764 323604 269816 323610
rect 269764 323546 269816 323552
rect 282932 313954 282960 702406
rect 300136 696250 300164 703520
rect 332520 700398 332548 703520
rect 348804 703050 348832 703520
rect 348792 703044 348844 703050
rect 348792 702986 348844 702992
rect 332508 700392 332560 700398
rect 332508 700334 332560 700340
rect 364996 700330 365024 703520
rect 397472 702846 397500 703520
rect 413664 702982 413692 703520
rect 413652 702976 413704 702982
rect 413652 702918 413704 702924
rect 397460 702840 397512 702846
rect 397460 702782 397512 702788
rect 429856 702778 429884 703520
rect 462332 702914 462360 703520
rect 462320 702908 462372 702914
rect 462320 702850 462372 702856
rect 429844 702772 429896 702778
rect 429844 702714 429896 702720
rect 478524 702710 478552 703520
rect 478512 702704 478564 702710
rect 478512 702646 478564 702652
rect 364984 700324 365036 700330
rect 364984 700266 365036 700272
rect 300124 696244 300176 696250
rect 300124 696186 300176 696192
rect 282920 313948 282972 313954
rect 282920 313890 282972 313896
rect 283564 307828 283616 307834
rect 283564 307770 283616 307776
rect 281540 305040 281592 305046
rect 281540 304982 281592 304988
rect 278780 303680 278832 303686
rect 278780 303622 278832 303628
rect 273260 302252 273312 302258
rect 273260 302194 273312 302200
rect 269120 289876 269172 289882
rect 269120 289818 269172 289824
rect 267740 259480 267792 259486
rect 267740 259422 267792 259428
rect 264244 235952 264296 235958
rect 264244 235894 264296 235900
rect 263692 220176 263744 220182
rect 263692 220118 263744 220124
rect 263600 157276 263652 157282
rect 263600 157218 263652 157224
rect 263704 146130 263732 220118
rect 266452 206304 266504 206310
rect 266452 206246 266504 206252
rect 266360 202292 266412 202298
rect 266360 202234 266412 202240
rect 264980 196648 265032 196654
rect 264980 196590 265032 196596
rect 264336 171216 264388 171222
rect 264336 171158 264388 171164
rect 264244 168428 264296 168434
rect 264244 168370 264296 168376
rect 263692 146124 263744 146130
rect 263692 146066 263744 146072
rect 264256 144226 264284 168370
rect 264244 144220 264296 144226
rect 264244 144162 264296 144168
rect 264244 136672 264296 136678
rect 264244 136614 264296 136620
rect 262956 120012 263008 120018
rect 262956 119954 263008 119960
rect 263048 119400 263100 119406
rect 263048 119342 263100 119348
rect 262864 115864 262916 115870
rect 262864 115806 262916 115812
rect 257528 110356 257580 110362
rect 257528 110298 257580 110304
rect 261484 109064 261536 109070
rect 261484 109006 261536 109012
rect 257436 102264 257488 102270
rect 257436 102206 257488 102212
rect 257344 102196 257396 102202
rect 257344 102138 257396 102144
rect 256056 99204 256108 99210
rect 256056 99146 256108 99152
rect 255964 97572 256016 97578
rect 255964 97514 256016 97520
rect 256056 96688 256108 96694
rect 256056 96630 256108 96636
rect 256068 17270 256096 96630
rect 257356 55962 257384 102138
rect 260104 98048 260156 98054
rect 260104 97990 260156 97996
rect 257344 55956 257396 55962
rect 257344 55898 257396 55904
rect 256056 17264 256108 17270
rect 256056 17206 256108 17212
rect 260116 15910 260144 97990
rect 260104 15904 260156 15910
rect 260104 15846 260156 15852
rect 261496 4894 261524 109006
rect 263060 97918 263088 119342
rect 263048 97912 263100 97918
rect 263048 97854 263100 97860
rect 264256 10402 264284 136614
rect 264348 133822 264376 171158
rect 264992 162790 265020 196590
rect 265072 181552 265124 181558
rect 265072 181494 265124 181500
rect 264980 162784 265032 162790
rect 264980 162726 265032 162732
rect 265084 158642 265112 181494
rect 265900 167068 265952 167074
rect 265900 167010 265952 167016
rect 265808 164484 265860 164490
rect 265808 164426 265860 164432
rect 265716 160200 265768 160206
rect 265716 160142 265768 160148
rect 265072 158636 265124 158642
rect 265072 158578 265124 158584
rect 264428 150544 264480 150550
rect 264428 150486 264480 150492
rect 264336 133816 264388 133822
rect 264336 133758 264388 133764
rect 264336 114572 264388 114578
rect 264336 114514 264388 114520
rect 264348 29646 264376 114514
rect 264440 112470 264468 150486
rect 265624 128376 265676 128382
rect 265624 128318 265676 128324
rect 264428 112464 264480 112470
rect 264428 112406 264480 112412
rect 265636 37942 265664 128318
rect 265728 121378 265756 160142
rect 265820 125526 265848 164426
rect 265912 128246 265940 167010
rect 266372 161430 266400 202234
rect 266464 165442 266492 206246
rect 266544 177472 266596 177478
rect 266544 177414 266596 177420
rect 266452 165436 266504 165442
rect 266452 165378 266504 165384
rect 266360 161424 266412 161430
rect 266360 161366 266412 161372
rect 266556 146198 266584 177414
rect 267004 173936 267056 173942
rect 267004 173878 267056 173884
rect 266544 146192 266596 146198
rect 266544 146134 266596 146140
rect 267016 136542 267044 173878
rect 267752 157350 267780 259422
rect 267924 188420 267976 188426
rect 267924 188362 267976 188368
rect 267832 177540 267884 177546
rect 267832 177482 267884 177488
rect 267740 157344 267792 157350
rect 267740 157286 267792 157292
rect 267096 145036 267148 145042
rect 267096 144978 267148 144984
rect 267004 136536 267056 136542
rect 267004 136478 267056 136484
rect 265900 128240 265952 128246
rect 265900 128182 265952 128188
rect 265808 125520 265860 125526
rect 265808 125462 265860 125468
rect 265716 121372 265768 121378
rect 265716 121314 265768 121320
rect 267004 120148 267056 120154
rect 267004 120090 267056 120096
rect 265716 116000 265768 116006
rect 265716 115942 265768 115948
rect 265624 37936 265676 37942
rect 265624 37878 265676 37884
rect 264336 29640 264388 29646
rect 264336 29582 264388 29588
rect 265728 28286 265756 115942
rect 267016 62898 267044 120090
rect 267108 103494 267136 144978
rect 267844 144838 267872 177482
rect 267936 164218 267964 188362
rect 267924 164212 267976 164218
rect 267924 164154 267976 164160
rect 268384 162988 268436 162994
rect 268384 162930 268436 162936
rect 267832 144832 267884 144838
rect 267832 144774 267884 144780
rect 268396 124166 268424 162930
rect 269132 143546 269160 289818
rect 270500 245676 270552 245682
rect 270500 245618 270552 245624
rect 269212 193860 269264 193866
rect 269212 193802 269264 193808
rect 269224 154494 269252 193802
rect 269304 188488 269356 188494
rect 269304 188430 269356 188436
rect 269316 162858 269344 188430
rect 269856 164348 269908 164354
rect 269856 164290 269908 164296
rect 269304 162852 269356 162858
rect 269304 162794 269356 162800
rect 269764 161560 269816 161566
rect 269764 161502 269816 161508
rect 269212 154488 269264 154494
rect 269212 154430 269264 154436
rect 269120 143540 269172 143546
rect 269120 143482 269172 143488
rect 268384 124160 268436 124166
rect 268384 124102 268436 124108
rect 269776 122738 269804 161502
rect 269868 126954 269896 164290
rect 270512 144906 270540 245618
rect 271880 211812 271932 211818
rect 271880 211754 271932 211760
rect 270592 203720 270644 203726
rect 270592 203662 270644 203668
rect 270604 155854 270632 203662
rect 271328 169856 271380 169862
rect 271328 169798 271380 169804
rect 271144 165708 271196 165714
rect 271144 165650 271196 165656
rect 270592 155848 270644 155854
rect 270592 155790 270644 155796
rect 270500 144900 270552 144906
rect 270500 144842 270552 144848
rect 269946 133104 270002 133113
rect 269946 133039 270002 133048
rect 269856 126948 269908 126954
rect 269856 126890 269908 126896
rect 269764 122732 269816 122738
rect 269764 122674 269816 122680
rect 268384 121508 268436 121514
rect 268384 121450 268436 121456
rect 267096 103488 267148 103494
rect 267096 103430 267148 103436
rect 267004 62892 267056 62898
rect 267004 62834 267056 62840
rect 268396 61402 268424 121450
rect 269396 112464 269448 112470
rect 269396 112406 269448 112412
rect 269408 107574 269436 112406
rect 269396 107568 269448 107574
rect 269396 107510 269448 107516
rect 269856 106344 269908 106350
rect 269856 106286 269908 106292
rect 269764 102264 269816 102270
rect 269764 102206 269816 102212
rect 268384 61396 268436 61402
rect 268384 61338 268436 61344
rect 265716 28280 265768 28286
rect 265716 28222 265768 28228
rect 269776 13122 269804 102206
rect 269868 66978 269896 106286
rect 269960 99346 269988 133039
rect 271156 128314 271184 165650
rect 271236 135312 271288 135318
rect 271236 135254 271288 135260
rect 271144 128308 271196 128314
rect 271144 128250 271196 128256
rect 271144 125656 271196 125662
rect 271144 125598 271196 125604
rect 269948 99340 270000 99346
rect 269948 99282 270000 99288
rect 269856 66972 269908 66978
rect 269856 66914 269908 66920
rect 271156 24138 271184 125598
rect 271248 54602 271276 135254
rect 271340 132394 271368 169798
rect 271892 149054 271920 211754
rect 271972 202224 272024 202230
rect 271972 202166 272024 202172
rect 271984 154426 272012 202166
rect 272524 167136 272576 167142
rect 272524 167078 272576 167084
rect 271972 154420 272024 154426
rect 271972 154362 272024 154368
rect 271880 149048 271932 149054
rect 271880 148990 271932 148996
rect 271328 132388 271380 132394
rect 271328 132330 271380 132336
rect 272536 129674 272564 167078
rect 273272 153202 273300 302194
rect 274640 298308 274692 298314
rect 274640 298250 274692 298256
rect 273352 198008 273404 198014
rect 273352 197950 273404 197956
rect 273260 153196 273312 153202
rect 273260 153138 273312 153144
rect 273364 146266 273392 197950
rect 273996 172644 274048 172650
rect 273996 172586 274048 172592
rect 273352 146260 273404 146266
rect 273352 146202 273404 146208
rect 273904 138032 273956 138038
rect 273904 137974 273956 137980
rect 272524 129668 272576 129674
rect 272524 129610 272576 129616
rect 272524 127016 272576 127022
rect 272524 126958 272576 126964
rect 271236 54596 271288 54602
rect 271236 54538 271288 54544
rect 272536 50386 272564 126958
rect 272524 50380 272576 50386
rect 272524 50322 272576 50328
rect 271144 24132 271196 24138
rect 271144 24074 271196 24080
rect 269764 13116 269816 13122
rect 269764 13058 269816 13064
rect 264244 10396 264296 10402
rect 264244 10338 264296 10344
rect 261484 4888 261536 4894
rect 261484 4830 261536 4836
rect 273916 3534 273944 137974
rect 274008 135250 274036 172586
rect 274088 146396 274140 146402
rect 274088 146338 274140 146344
rect 274100 138689 274128 146338
rect 274086 138680 274142 138689
rect 274086 138615 274142 138624
rect 274652 137902 274680 298250
rect 278044 295452 278096 295458
rect 278044 295394 278096 295400
rect 276020 227112 276072 227118
rect 276020 227054 276072 227060
rect 274732 203652 274784 203658
rect 274732 203594 274784 203600
rect 274744 147558 274772 203594
rect 275284 158840 275336 158846
rect 275284 158782 275336 158788
rect 274732 147552 274784 147558
rect 274732 147494 274784 147500
rect 275296 141438 275324 158782
rect 276032 158710 276060 227054
rect 277400 217388 277452 217394
rect 277400 217330 277452 217336
rect 276020 158704 276072 158710
rect 276020 158646 276072 158652
rect 275376 156052 275428 156058
rect 275376 155994 275428 156000
rect 275284 141432 275336 141438
rect 275284 141374 275336 141380
rect 274640 137896 274692 137902
rect 274640 137838 274692 137844
rect 273996 135244 274048 135250
rect 273996 135186 274048 135192
rect 275284 133952 275336 133958
rect 275284 133894 275336 133900
rect 273996 128444 274048 128450
rect 273996 128386 274048 128392
rect 274008 21418 274036 128386
rect 275296 42158 275324 133894
rect 275388 115938 275416 155994
rect 276756 141432 276808 141438
rect 276756 141374 276808 141380
rect 276664 129804 276716 129810
rect 276664 129746 276716 129752
rect 275376 115932 275428 115938
rect 275376 115874 275428 115880
rect 275284 42152 275336 42158
rect 275284 42094 275336 42100
rect 276676 36582 276704 129746
rect 276768 114442 276796 141374
rect 277412 137970 277440 217330
rect 277400 137964 277452 137970
rect 277400 137906 277452 137912
rect 276756 114436 276808 114442
rect 276756 114378 276808 114384
rect 278056 96626 278084 295394
rect 278228 174004 278280 174010
rect 278228 173946 278280 173952
rect 278240 138718 278268 173946
rect 278792 155922 278820 303622
rect 280160 235408 280212 235414
rect 280160 235350 280212 235356
rect 278872 213308 278924 213314
rect 278872 213250 278924 213256
rect 278780 155916 278832 155922
rect 278780 155858 278832 155864
rect 278884 150414 278912 213250
rect 279608 168496 279660 168502
rect 279608 168438 279660 168444
rect 278872 150408 278924 150414
rect 278872 150350 278924 150356
rect 278228 138712 278280 138718
rect 278228 138654 278280 138660
rect 278136 138100 278188 138106
rect 278136 138042 278188 138048
rect 278044 96620 278096 96626
rect 278044 96562 278096 96568
rect 276664 36576 276716 36582
rect 276664 36518 276716 36524
rect 273996 21412 274048 21418
rect 273996 21354 274048 21360
rect 278148 11830 278176 138042
rect 279516 131164 279568 131170
rect 279516 131106 279568 131112
rect 279424 129872 279476 129878
rect 279424 129814 279476 129820
rect 278228 109132 278280 109138
rect 278228 109074 278280 109080
rect 278240 25634 278268 109074
rect 278228 25628 278280 25634
rect 278228 25570 278280 25576
rect 279436 18630 279464 129814
rect 279528 44878 279556 131106
rect 279620 131034 279648 168438
rect 279700 144220 279752 144226
rect 279700 144162 279752 144168
rect 279608 131028 279660 131034
rect 279608 130970 279660 130976
rect 279608 113212 279660 113218
rect 279608 113154 279660 113160
rect 279620 51746 279648 113154
rect 279712 106282 279740 144162
rect 280172 139398 280200 235350
rect 280896 147756 280948 147762
rect 280896 147698 280948 147704
rect 280804 139460 280856 139466
rect 280804 139402 280856 139408
rect 280160 139392 280212 139398
rect 280160 139334 280212 139340
rect 279700 106276 279752 106282
rect 279700 106218 279752 106224
rect 279608 51740 279660 51746
rect 279608 51682 279660 51688
rect 279516 44872 279568 44878
rect 279516 44814 279568 44820
rect 279424 18624 279476 18630
rect 279424 18566 279476 18572
rect 280816 13190 280844 139402
rect 280908 107642 280936 147698
rect 281552 147626 281580 304982
rect 283576 181490 283604 307770
rect 342260 306400 342312 306406
rect 342260 306342 342312 306348
rect 319444 300892 319496 300898
rect 319444 300834 319496 300840
rect 308404 299600 308456 299606
rect 308404 299542 308456 299548
rect 307024 282940 307076 282946
rect 307024 282882 307076 282888
rect 305644 249076 305696 249082
rect 305644 249018 305696 249024
rect 287704 223032 287756 223038
rect 287704 222974 287756 222980
rect 283564 181484 283616 181490
rect 283564 181426 283616 181432
rect 287716 180334 287744 222974
rect 291844 215960 291896 215966
rect 291844 215902 291896 215908
rect 291856 181558 291884 215902
rect 300124 209160 300176 209166
rect 300124 209102 300176 209108
rect 291844 181552 291896 181558
rect 291844 181494 291896 181500
rect 300136 181393 300164 209102
rect 300122 181384 300178 181393
rect 300122 181319 300178 181328
rect 287704 180328 287756 180334
rect 287704 180270 287756 180276
rect 305656 178809 305684 249018
rect 305642 178800 305698 178809
rect 305642 178735 305698 178744
rect 307036 177410 307064 282882
rect 307116 210520 307168 210526
rect 307116 210462 307168 210468
rect 307128 178673 307156 210462
rect 307114 178664 307170 178673
rect 307114 178599 307170 178608
rect 307024 177404 307076 177410
rect 307024 177346 307076 177352
rect 307022 175264 307078 175273
rect 307022 175199 307078 175208
rect 306746 174856 306802 174865
rect 306746 174791 306802 174800
rect 291844 174072 291896 174078
rect 291844 174014 291896 174020
rect 282184 172712 282236 172718
rect 282184 172654 282236 172660
rect 282196 155281 282224 172654
rect 289268 171284 289320 171290
rect 289268 171226 289320 171232
rect 287888 169924 287940 169930
rect 287888 169866 287940 169872
rect 283564 168564 283616 168570
rect 283564 168506 283616 168512
rect 282182 155272 282238 155281
rect 282182 155207 282238 155216
rect 282368 154692 282420 154698
rect 282368 154634 282420 154640
rect 281540 147620 281592 147626
rect 281540 147562 281592 147568
rect 282276 136740 282328 136746
rect 282276 136682 282328 136688
rect 282184 114640 282236 114646
rect 282184 114582 282236 114588
rect 280896 107636 280948 107642
rect 280896 107578 280948 107584
rect 280896 105052 280948 105058
rect 280896 104994 280948 105000
rect 280908 15978 280936 104994
rect 280896 15972 280948 15978
rect 280896 15914 280948 15920
rect 280804 13184 280856 13190
rect 280804 13126 280856 13132
rect 278136 11824 278188 11830
rect 278136 11766 278188 11772
rect 282196 6186 282224 114582
rect 282288 46238 282316 136682
rect 282380 114510 282408 154634
rect 282460 149116 282512 149122
rect 282460 149058 282512 149064
rect 282368 114504 282420 114510
rect 282368 114446 282420 114452
rect 282472 108934 282500 149058
rect 283576 129742 283604 168506
rect 283656 167204 283708 167210
rect 283656 167146 283708 167152
rect 283668 134570 283696 167146
rect 285036 160744 285088 160750
rect 285036 160686 285088 160692
rect 284944 135380 284996 135386
rect 284944 135322 284996 135328
rect 283656 134564 283708 134570
rect 283656 134506 283708 134512
rect 283748 134020 283800 134026
rect 283748 133962 283800 133968
rect 283564 129736 283616 129742
rect 283564 129678 283616 129684
rect 283564 122868 283616 122874
rect 283564 122810 283616 122816
rect 282460 108928 282512 108934
rect 282460 108870 282512 108876
rect 282368 107908 282420 107914
rect 282368 107850 282420 107856
rect 282380 65550 282408 107850
rect 282368 65544 282420 65550
rect 282368 65486 282420 65492
rect 282276 46232 282328 46238
rect 282276 46174 282328 46180
rect 283576 14482 283604 122810
rect 283656 106412 283708 106418
rect 283656 106354 283708 106360
rect 283668 22778 283696 106354
rect 283760 57254 283788 133962
rect 283748 57248 283800 57254
rect 283748 57190 283800 57196
rect 284956 53174 284984 135322
rect 285048 131102 285076 160686
rect 286416 143608 286468 143614
rect 286416 143550 286468 143556
rect 286324 142248 286376 142254
rect 286324 142190 286376 142196
rect 285036 131096 285088 131102
rect 285036 131038 285088 131044
rect 285036 127084 285088 127090
rect 285036 127026 285088 127032
rect 284944 53168 284996 53174
rect 284944 53110 284996 53116
rect 285048 49026 285076 127026
rect 286336 102066 286364 142190
rect 286428 104174 286456 143550
rect 287704 132524 287756 132530
rect 287704 132466 287756 132472
rect 286416 104168 286468 104174
rect 286416 104110 286468 104116
rect 286324 102060 286376 102066
rect 286324 102002 286376 102008
rect 286416 100768 286468 100774
rect 286416 100710 286468 100716
rect 286324 98116 286376 98122
rect 286324 98058 286376 98064
rect 285036 49020 285088 49026
rect 285036 48962 285088 48968
rect 283656 22772 283708 22778
rect 283656 22714 283708 22720
rect 283564 14476 283616 14482
rect 283564 14418 283616 14424
rect 286336 11762 286364 98058
rect 286428 64190 286456 100710
rect 286416 64184 286468 64190
rect 286416 64126 286468 64132
rect 286324 11756 286376 11762
rect 286324 11698 286376 11704
rect 287716 7614 287744 132466
rect 287900 132462 287928 169866
rect 289176 150612 289228 150618
rect 289176 150554 289228 150560
rect 287980 146940 288032 146946
rect 287980 146882 288032 146888
rect 287888 132456 287940 132462
rect 287888 132398 287940 132404
rect 287796 131232 287848 131238
rect 287796 131174 287848 131180
rect 287808 25566 287836 131174
rect 287992 121446 288020 146882
rect 289084 139528 289136 139534
rect 289084 139470 289136 139476
rect 287980 121440 288032 121446
rect 287980 121382 288032 121388
rect 287888 120216 287940 120222
rect 287888 120158 287940 120164
rect 287900 50454 287928 120158
rect 287980 103624 288032 103630
rect 287980 103566 288032 103572
rect 287992 68406 288020 103566
rect 287980 68400 288032 68406
rect 287980 68342 288032 68348
rect 287888 50448 287940 50454
rect 287888 50390 287940 50396
rect 287796 25560 287848 25566
rect 287796 25502 287848 25508
rect 289096 10334 289124 139470
rect 289188 110430 289216 150554
rect 289280 133890 289308 171226
rect 291856 136610 291884 174014
rect 306760 174010 306788 174791
rect 306748 174004 306800 174010
rect 306748 173946 306800 173952
rect 306930 173224 306986 173233
rect 306930 173159 306986 173168
rect 306944 172582 306972 173159
rect 306932 172576 306984 172582
rect 306932 172518 306984 172524
rect 306930 171048 306986 171057
rect 306930 170983 306986 170992
rect 306944 169930 306972 170983
rect 306932 169924 306984 169930
rect 306932 169866 306984 169872
rect 293224 165776 293276 165782
rect 293224 165718 293276 165724
rect 291936 156120 291988 156126
rect 291936 156062 291988 156068
rect 291844 136604 291896 136610
rect 291844 136546 291896 136552
rect 290648 134088 290700 134094
rect 290648 134030 290700 134036
rect 289268 133884 289320 133890
rect 289268 133826 289320 133832
rect 290556 129940 290608 129946
rect 290556 129882 290608 129888
rect 289360 125724 289412 125730
rect 289360 125666 289412 125672
rect 289176 110424 289228 110430
rect 289176 110366 289228 110372
rect 289176 104984 289228 104990
rect 289176 104926 289228 104932
rect 289188 18698 289216 104926
rect 289268 99408 289320 99414
rect 289268 99350 289320 99356
rect 289280 35222 289308 99350
rect 289372 72554 289400 125666
rect 290464 124228 290516 124234
rect 290464 124170 290516 124176
rect 289360 72548 289412 72554
rect 289360 72490 289412 72496
rect 289268 35216 289320 35222
rect 289268 35158 289320 35164
rect 289176 18692 289228 18698
rect 289176 18634 289228 18640
rect 289084 10328 289136 10334
rect 289084 10270 289136 10276
rect 287704 7608 287756 7614
rect 287704 7550 287756 7556
rect 282184 6180 282236 6186
rect 282184 6122 282236 6128
rect 273904 3528 273956 3534
rect 273904 3470 273956 3476
rect 253204 3460 253256 3466
rect 253204 3402 253256 3408
rect 290476 2174 290504 124170
rect 290568 26926 290596 129882
rect 290660 76634 290688 134030
rect 291844 131300 291896 131306
rect 291844 131242 291896 131248
rect 290648 76628 290700 76634
rect 290648 76570 290700 76576
rect 291856 43450 291884 131242
rect 291948 117298 291976 156062
rect 293236 142866 293264 165718
rect 306562 165064 306618 165073
rect 306562 164999 306618 165008
rect 294788 164416 294840 164422
rect 294788 164358 294840 164364
rect 293592 157548 293644 157554
rect 293592 157490 293644 157496
rect 293224 142860 293276 142866
rect 293224 142802 293276 142808
rect 293498 142760 293554 142769
rect 293498 142695 293554 142704
rect 292118 141400 292174 141409
rect 292118 141335 292174 141344
rect 291936 117292 291988 117298
rect 291936 117234 291988 117240
rect 292028 116068 292080 116074
rect 292028 116010 292080 116016
rect 291936 113280 291988 113286
rect 291936 113222 291988 113228
rect 291948 47598 291976 113222
rect 292040 58682 292068 116010
rect 292132 100638 292160 141335
rect 293224 132592 293276 132598
rect 293224 132534 293276 132540
rect 292120 100632 292172 100638
rect 292120 100574 292172 100580
rect 292120 96756 292172 96762
rect 292120 96698 292172 96704
rect 292028 58676 292080 58682
rect 292028 58618 292080 58624
rect 292132 54534 292160 96698
rect 292120 54528 292172 54534
rect 292120 54470 292172 54476
rect 291936 47592 291988 47598
rect 291936 47534 291988 47540
rect 291844 43444 291896 43450
rect 291844 43386 291896 43392
rect 290556 26920 290608 26926
rect 290556 26862 290608 26868
rect 293236 8974 293264 132534
rect 293316 121576 293368 121582
rect 293316 121518 293368 121524
rect 293328 40798 293356 121518
rect 293408 117360 293460 117366
rect 293408 117302 293460 117308
rect 293420 71126 293448 117302
rect 293512 102134 293540 142695
rect 293604 118658 293632 157490
rect 294604 128512 294656 128518
rect 294604 128454 294656 128460
rect 293592 118652 293644 118658
rect 293592 118594 293644 118600
rect 293500 102128 293552 102134
rect 293500 102070 293552 102076
rect 293592 100836 293644 100842
rect 293592 100778 293644 100784
rect 293408 71120 293460 71126
rect 293408 71062 293460 71068
rect 293604 66910 293632 100778
rect 293592 66904 293644 66910
rect 293592 66846 293644 66852
rect 293316 40792 293368 40798
rect 293316 40734 293368 40740
rect 294616 39370 294644 128454
rect 294800 126274 294828 164358
rect 306576 164286 306604 164999
rect 304356 164280 304408 164286
rect 304356 164222 304408 164228
rect 306564 164280 306616 164286
rect 306564 164222 306616 164228
rect 300124 163056 300176 163062
rect 300124 162998 300176 163004
rect 296076 161628 296128 161634
rect 296076 161570 296128 161576
rect 295984 127152 296036 127158
rect 295984 127094 296036 127100
rect 294788 126268 294840 126274
rect 294788 126210 294840 126216
rect 294696 125792 294748 125798
rect 294696 125734 294748 125740
rect 294708 73846 294736 125734
rect 294788 98184 294840 98190
rect 294788 98126 294840 98132
rect 294696 73840 294748 73846
rect 294696 73782 294748 73788
rect 294800 53106 294828 98126
rect 294788 53100 294840 53106
rect 294788 53042 294840 53048
rect 295996 40730 296024 127094
rect 296088 122806 296116 161570
rect 296260 158908 296312 158914
rect 296260 158850 296312 158856
rect 296076 122800 296128 122806
rect 296076 122742 296128 122748
rect 296272 120086 296300 158850
rect 298836 154760 298888 154766
rect 298836 154702 298888 154708
rect 297640 149184 297692 149190
rect 297640 149126 297692 149132
rect 297364 135448 297416 135454
rect 297364 135390 297416 135396
rect 296260 120080 296312 120086
rect 296260 120022 296312 120028
rect 296168 118856 296220 118862
rect 296168 118798 296220 118804
rect 296076 117428 296128 117434
rect 296076 117370 296128 117376
rect 295984 40724 296036 40730
rect 295984 40666 296036 40672
rect 294604 39364 294656 39370
rect 294604 39306 294656 39312
rect 296088 33794 296116 117370
rect 296180 36650 296208 118798
rect 296260 110492 296312 110498
rect 296260 110434 296312 110440
rect 296168 36644 296220 36650
rect 296168 36586 296220 36592
rect 296076 33788 296128 33794
rect 296076 33730 296128 33736
rect 296272 28354 296300 110434
rect 297376 39438 297404 135390
rect 297548 121644 297600 121650
rect 297548 121586 297600 121592
rect 297456 111852 297508 111858
rect 297456 111794 297508 111800
rect 297364 39432 297416 39438
rect 297364 39374 297416 39380
rect 297468 29714 297496 111794
rect 297560 49094 297588 121586
rect 297652 111110 297680 149126
rect 298744 138168 298796 138174
rect 298744 138110 298796 138116
rect 297640 111104 297692 111110
rect 297640 111046 297692 111052
rect 297548 49088 297600 49094
rect 297548 49030 297600 49036
rect 298756 33862 298784 138110
rect 298848 117978 298876 154702
rect 300136 124914 300164 162998
rect 301596 153332 301648 153338
rect 301596 153274 301648 153280
rect 301504 151972 301556 151978
rect 301504 151914 301556 151920
rect 300492 146124 300544 146130
rect 300492 146066 300544 146072
rect 300124 124908 300176 124914
rect 300124 124850 300176 124856
rect 300308 124364 300360 124370
rect 300308 124306 300360 124312
rect 300216 123004 300268 123010
rect 300216 122946 300268 122952
rect 299020 118788 299072 118794
rect 299020 118730 299072 118736
rect 298836 117972 298888 117978
rect 298836 117914 298888 117920
rect 298836 113348 298888 113354
rect 298836 113290 298888 113296
rect 298744 33856 298796 33862
rect 298744 33798 298796 33804
rect 298848 32434 298876 113290
rect 298928 102332 298980 102338
rect 298928 102274 298980 102280
rect 298836 32428 298888 32434
rect 298836 32370 298888 32376
rect 298940 31074 298968 102274
rect 299032 69698 299060 118730
rect 300124 111920 300176 111926
rect 300124 111862 300176 111868
rect 299020 69692 299072 69698
rect 299020 69634 299072 69640
rect 298928 31068 298980 31074
rect 298928 31010 298980 31016
rect 297456 29708 297508 29714
rect 297456 29650 297508 29656
rect 296260 28348 296312 28354
rect 296260 28290 296312 28296
rect 300136 26994 300164 111862
rect 300228 42090 300256 122946
rect 300320 60042 300348 124306
rect 300400 117496 300452 117502
rect 300400 117438 300452 117444
rect 300308 60036 300360 60042
rect 300308 59978 300360 59984
rect 300412 55894 300440 117438
rect 300504 113150 300532 146066
rect 300492 113144 300544 113150
rect 300492 113086 300544 113092
rect 301516 111790 301544 151914
rect 301608 123486 301636 153274
rect 303068 147824 303120 147830
rect 303068 147766 303120 147772
rect 302884 135516 302936 135522
rect 302884 135458 302936 135464
rect 301596 123480 301648 123486
rect 301596 123422 301648 123428
rect 301688 120284 301740 120290
rect 301688 120226 301740 120232
rect 301504 111784 301556 111790
rect 301504 111726 301556 111732
rect 301596 107772 301648 107778
rect 301596 107714 301648 107720
rect 301504 106480 301556 106486
rect 301504 106422 301556 106428
rect 300400 55888 300452 55894
rect 300400 55830 300452 55836
rect 300216 42084 300268 42090
rect 300216 42026 300268 42032
rect 300124 26988 300176 26994
rect 300124 26930 300176 26936
rect 301516 21486 301544 106422
rect 301608 24206 301636 107714
rect 301700 38010 301728 120226
rect 301780 110628 301832 110634
rect 301780 110570 301832 110576
rect 301792 58750 301820 110570
rect 301780 58744 301832 58750
rect 301780 58686 301832 58692
rect 302896 47666 302924 135458
rect 302976 122936 303028 122942
rect 302976 122878 303028 122884
rect 302884 47660 302936 47666
rect 302884 47602 302936 47608
rect 302988 44946 303016 122878
rect 303080 109002 303108 147766
rect 304368 125594 304396 164222
rect 306562 160848 306618 160857
rect 306562 160783 306618 160792
rect 306576 160138 306604 160783
rect 306564 160132 306616 160138
rect 306564 160074 306616 160080
rect 306930 160032 306986 160041
rect 306930 159967 306986 159976
rect 306944 158778 306972 159967
rect 306932 158772 306984 158778
rect 306932 158714 306984 158720
rect 306930 158672 306986 158681
rect 306930 158607 306986 158616
rect 306944 157486 306972 158607
rect 306932 157480 306984 157486
rect 306932 157422 306984 157428
rect 306746 157040 306802 157049
rect 306746 156975 306802 156984
rect 306760 156126 306788 156975
rect 306748 156120 306800 156126
rect 306748 156062 306800 156068
rect 306654 153232 306710 153241
rect 306654 153167 306710 153176
rect 305826 146432 305882 146441
rect 305826 146367 305882 146376
rect 304448 139596 304500 139602
rect 304448 139538 304500 139544
rect 304356 125588 304408 125594
rect 304356 125530 304408 125536
rect 304264 124296 304316 124302
rect 304264 124238 304316 124244
rect 303160 110560 303212 110566
rect 303160 110502 303212 110508
rect 303068 108996 303120 109002
rect 303068 108938 303120 108944
rect 303068 100904 303120 100910
rect 303068 100846 303120 100852
rect 303080 62830 303108 100846
rect 303172 75206 303200 110502
rect 303160 75200 303212 75206
rect 303160 75142 303212 75148
rect 303068 62824 303120 62830
rect 303068 62766 303120 62772
rect 302976 44940 303028 44946
rect 302976 44882 303028 44888
rect 301688 38004 301740 38010
rect 301688 37946 301740 37952
rect 301596 24200 301648 24206
rect 301596 24142 301648 24148
rect 301504 21480 301556 21486
rect 301504 21422 301556 21428
rect 304276 19990 304304 124238
rect 304356 107704 304408 107710
rect 304356 107646 304408 107652
rect 304368 31142 304396 107646
rect 304460 100706 304488 139538
rect 305734 118960 305790 118969
rect 305734 118895 305790 118904
rect 304540 109200 304592 109206
rect 304540 109142 304592 109148
rect 304448 100700 304500 100706
rect 304448 100642 304500 100648
rect 304552 73914 304580 109142
rect 305642 105496 305698 105505
rect 305642 105431 305698 105440
rect 304632 99476 304684 99482
rect 304632 99418 304684 99424
rect 304540 73908 304592 73914
rect 304540 73850 304592 73856
rect 304644 68338 304672 99418
rect 304632 68332 304684 68338
rect 304632 68274 304684 68280
rect 304356 31136 304408 31142
rect 304356 31078 304408 31084
rect 304264 19984 304316 19990
rect 304264 19926 304316 19932
rect 305656 17338 305684 105431
rect 305748 35290 305776 118895
rect 305840 105602 305868 146367
rect 306668 146130 306696 153167
rect 306930 150648 306986 150657
rect 306930 150583 306986 150592
rect 306944 150482 306972 150583
rect 306932 150476 306984 150482
rect 306932 150418 306984 150424
rect 306930 150240 306986 150249
rect 306930 150175 306986 150184
rect 306944 149122 306972 150175
rect 307036 149734 307064 175199
rect 307666 174448 307722 174457
rect 307666 174383 307722 174392
rect 307680 174078 307708 174383
rect 307668 174072 307720 174078
rect 307574 174040 307630 174049
rect 307668 174014 307720 174020
rect 307574 173975 307630 173984
rect 307588 173942 307616 173975
rect 307576 173936 307628 173942
rect 307576 173878 307628 173884
rect 307666 173632 307722 173641
rect 307666 173567 307722 173576
rect 307300 172712 307352 172718
rect 307298 172680 307300 172689
rect 307352 172680 307354 172689
rect 307680 172650 307708 173567
rect 307298 172615 307354 172624
rect 307668 172644 307720 172650
rect 307668 172586 307720 172592
rect 307482 172272 307538 172281
rect 307482 172207 307538 172216
rect 307496 171290 307524 172207
rect 307574 171864 307630 171873
rect 307574 171799 307630 171808
rect 307484 171284 307536 171290
rect 307484 171226 307536 171232
rect 307588 171222 307616 171799
rect 307666 171456 307722 171465
rect 307666 171391 307722 171400
rect 307576 171216 307628 171222
rect 307576 171158 307628 171164
rect 307680 171154 307708 171391
rect 307668 171148 307720 171154
rect 307668 171090 307720 171096
rect 307482 170640 307538 170649
rect 307482 170575 307538 170584
rect 307496 169862 307524 170575
rect 307666 170232 307722 170241
rect 307666 170167 307722 170176
rect 307484 169856 307536 169862
rect 307206 169824 307262 169833
rect 307484 169798 307536 169804
rect 307680 169794 307708 170167
rect 307206 169759 307262 169768
rect 307668 169788 307720 169794
rect 307220 160750 307248 169759
rect 307668 169730 307720 169736
rect 307482 169280 307538 169289
rect 307482 169215 307538 169224
rect 307300 168564 307352 168570
rect 307300 168506 307352 168512
rect 307312 168473 307340 168506
rect 307496 168502 307524 169215
rect 307666 168872 307722 168881
rect 307666 168807 307722 168816
rect 307484 168496 307536 168502
rect 307298 168464 307354 168473
rect 307484 168438 307536 168444
rect 307680 168434 307708 168807
rect 307298 168399 307354 168408
rect 307668 168428 307720 168434
rect 307668 168370 307720 168376
rect 307482 168056 307538 168065
rect 307482 167991 307538 168000
rect 307496 167142 307524 167991
rect 307574 167648 307630 167657
rect 307574 167583 307630 167592
rect 307484 167136 307536 167142
rect 307484 167078 307536 167084
rect 307588 167074 307616 167583
rect 307666 167240 307722 167249
rect 307666 167175 307668 167184
rect 307720 167175 307722 167184
rect 307668 167146 307720 167152
rect 307576 167068 307628 167074
rect 307576 167010 307628 167016
rect 307666 166832 307722 166841
rect 307666 166767 307722 166776
rect 307482 166424 307538 166433
rect 307482 166359 307538 166368
rect 307298 165880 307354 165889
rect 307298 165815 307354 165824
rect 307312 165782 307340 165815
rect 307300 165776 307352 165782
rect 307300 165718 307352 165724
rect 307496 165646 307524 166359
rect 307680 165714 307708 166767
rect 307668 165708 307720 165714
rect 307668 165650 307720 165656
rect 307484 165640 307536 165646
rect 307484 165582 307536 165588
rect 307482 165472 307538 165481
rect 307482 165407 307538 165416
rect 307496 164354 307524 165407
rect 307666 164656 307722 164665
rect 307666 164591 307722 164600
rect 307680 164490 307708 164591
rect 307668 164484 307720 164490
rect 307668 164426 307720 164432
rect 307576 164416 307628 164422
rect 307576 164358 307628 164364
rect 307484 164348 307536 164354
rect 307484 164290 307536 164296
rect 307588 164257 307616 164358
rect 307574 164248 307630 164257
rect 307574 164183 307630 164192
rect 307482 163840 307538 163849
rect 307482 163775 307538 163784
rect 307496 163062 307524 163775
rect 307666 163432 307722 163441
rect 307666 163367 307722 163376
rect 307484 163056 307536 163062
rect 307298 163024 307354 163033
rect 307484 162998 307536 163004
rect 307680 162994 307708 163367
rect 307298 162959 307354 162968
rect 307668 162988 307720 162994
rect 307312 162926 307340 162959
rect 307668 162930 307720 162936
rect 307300 162920 307352 162926
rect 307300 162862 307352 162868
rect 307482 162480 307538 162489
rect 307482 162415 307538 162424
rect 307298 162072 307354 162081
rect 307298 162007 307354 162016
rect 307312 161566 307340 162007
rect 307496 161634 307524 162415
rect 307666 161664 307722 161673
rect 307484 161628 307536 161634
rect 307666 161599 307722 161608
rect 307484 161570 307536 161576
rect 307300 161560 307352 161566
rect 307300 161502 307352 161508
rect 307680 161498 307708 161599
rect 307668 161492 307720 161498
rect 307668 161434 307720 161440
rect 307666 161256 307722 161265
rect 307666 161191 307722 161200
rect 307208 160744 307260 160750
rect 307208 160686 307260 160692
rect 307114 160440 307170 160449
rect 307114 160375 307170 160384
rect 307024 149728 307076 149734
rect 307024 149670 307076 149676
rect 306932 149116 306984 149122
rect 306932 149058 306984 149064
rect 306930 148880 306986 148889
rect 306930 148815 306986 148824
rect 306944 147694 306972 148815
rect 307022 148472 307078 148481
rect 307022 148407 307078 148416
rect 306932 147688 306984 147694
rect 306932 147630 306984 147636
rect 306746 147248 306802 147257
rect 306746 147183 306802 147192
rect 306760 146334 306788 147183
rect 306748 146328 306800 146334
rect 306748 146270 306800 146276
rect 306656 146124 306708 146130
rect 306656 146066 306708 146072
rect 306562 144664 306618 144673
rect 306562 144599 306618 144608
rect 305920 140888 305972 140894
rect 305920 140830 305972 140836
rect 305828 105596 305880 105602
rect 305828 105538 305880 105544
rect 305932 104854 305960 140830
rect 306576 140078 306604 144599
rect 306746 143032 306802 143041
rect 306746 142967 306802 142976
rect 306760 142186 306788 142967
rect 306748 142180 306800 142186
rect 306748 142122 306800 142128
rect 306564 140072 306616 140078
rect 306564 140014 306616 140020
rect 306930 137864 306986 137873
rect 306930 137799 306986 137808
rect 306944 136678 306972 137799
rect 306932 136672 306984 136678
rect 306932 136614 306984 136620
rect 306746 134872 306802 134881
rect 306746 134807 306802 134816
rect 306760 133958 306788 134807
rect 306748 133952 306800 133958
rect 306748 133894 306800 133900
rect 306746 131472 306802 131481
rect 306746 131407 306802 131416
rect 306760 131306 306788 131407
rect 306748 131300 306800 131306
rect 306748 131242 306800 131248
rect 306746 131064 306802 131073
rect 306746 130999 306802 131008
rect 306760 129946 306788 130999
rect 306930 130248 306986 130257
rect 306930 130183 306986 130192
rect 306748 129940 306800 129946
rect 306748 129882 306800 129888
rect 306944 129878 306972 130183
rect 306932 129872 306984 129878
rect 306932 129814 306984 129820
rect 306746 125896 306802 125905
rect 306746 125831 306802 125840
rect 306760 125730 306788 125831
rect 306748 125724 306800 125730
rect 306748 125666 306800 125672
rect 306746 125488 306802 125497
rect 306746 125423 306802 125432
rect 306760 124370 306788 125423
rect 306748 124364 306800 124370
rect 306748 124306 306800 124312
rect 306562 123856 306618 123865
rect 306562 123791 306618 123800
rect 306576 122874 306604 123791
rect 306564 122868 306616 122874
rect 306564 122810 306616 122816
rect 306746 120048 306802 120057
rect 306746 119983 306802 119992
rect 306760 118862 306788 119983
rect 306748 118856 306800 118862
rect 306748 118798 306800 118804
rect 306746 116648 306802 116657
rect 306746 116583 306802 116592
rect 306760 116006 306788 116583
rect 306748 116000 306800 116006
rect 306748 115942 306800 115948
rect 306746 115696 306802 115705
rect 306746 115631 306802 115640
rect 306760 114578 306788 115631
rect 306748 114572 306800 114578
rect 306748 114514 306800 114520
rect 306746 114472 306802 114481
rect 306746 114407 306802 114416
rect 306760 113354 306788 114407
rect 306748 113348 306800 113354
rect 306748 113290 306800 113296
rect 307036 112470 307064 148407
rect 307128 146946 307156 160375
rect 307680 160206 307708 161191
rect 307668 160200 307720 160206
rect 307668 160142 307720 160148
rect 307482 159624 307538 159633
rect 307482 159559 307538 159568
rect 307496 158846 307524 159559
rect 307666 159080 307722 159089
rect 307666 159015 307722 159024
rect 307680 158914 307708 159015
rect 307668 158908 307720 158914
rect 307668 158850 307720 158856
rect 307484 158840 307536 158846
rect 307484 158782 307536 158788
rect 307482 158264 307538 158273
rect 307482 158199 307538 158208
rect 307298 157856 307354 157865
rect 307298 157791 307354 157800
rect 307312 157418 307340 157791
rect 307496 157554 307524 158199
rect 307484 157548 307536 157554
rect 307484 157490 307536 157496
rect 307390 157448 307446 157457
rect 307300 157412 307352 157418
rect 307390 157383 307446 157392
rect 307300 157354 307352 157360
rect 307206 154456 307262 154465
rect 307206 154391 307262 154400
rect 307116 146940 307168 146946
rect 307116 146882 307168 146888
rect 307220 141438 307248 154391
rect 307404 153882 307432 157383
rect 307574 156632 307630 156641
rect 307574 156567 307630 156576
rect 307588 155990 307616 156567
rect 307666 156224 307722 156233
rect 307666 156159 307722 156168
rect 307680 156058 307708 156159
rect 307668 156052 307720 156058
rect 307668 155994 307720 156000
rect 307576 155984 307628 155990
rect 307576 155926 307628 155932
rect 307482 155680 307538 155689
rect 307482 155615 307538 155624
rect 307496 154630 307524 155615
rect 307574 155272 307630 155281
rect 307574 155207 307630 155216
rect 307588 154766 307616 155207
rect 307666 154864 307722 154873
rect 307666 154799 307722 154808
rect 307576 154760 307628 154766
rect 307576 154702 307628 154708
rect 307680 154698 307708 154799
rect 307668 154692 307720 154698
rect 307668 154634 307720 154640
rect 307484 154624 307536 154630
rect 307484 154566 307536 154572
rect 307482 154048 307538 154057
rect 307482 153983 307538 153992
rect 307392 153876 307444 153882
rect 307392 153818 307444 153824
rect 307496 153270 307524 153983
rect 307666 153640 307722 153649
rect 307666 153575 307722 153584
rect 307680 153338 307708 153575
rect 307668 153332 307720 153338
rect 307668 153274 307720 153280
rect 307484 153264 307536 153270
rect 307484 153206 307536 153212
rect 307482 152688 307538 152697
rect 307482 152623 307538 152632
rect 307496 151910 307524 152623
rect 307666 152280 307722 152289
rect 307666 152215 307722 152224
rect 307680 151978 307708 152215
rect 307668 151972 307720 151978
rect 307668 151914 307720 151920
rect 307484 151904 307536 151910
rect 307484 151846 307536 151852
rect 307666 151872 307722 151881
rect 307666 151807 307668 151816
rect 307720 151807 307722 151816
rect 307668 151778 307720 151784
rect 307482 151464 307538 151473
rect 307482 151399 307538 151408
rect 307496 150618 307524 151399
rect 307666 151056 307722 151065
rect 307666 150991 307722 151000
rect 307484 150612 307536 150618
rect 307484 150554 307536 150560
rect 307680 150550 307708 150991
rect 307668 150544 307720 150550
rect 307668 150486 307720 150492
rect 307666 149832 307722 149841
rect 307666 149767 307722 149776
rect 307574 149288 307630 149297
rect 307574 149223 307630 149232
rect 307588 147830 307616 149223
rect 307680 149190 307708 149767
rect 307668 149184 307720 149190
rect 307668 149126 307720 149132
rect 307666 148064 307722 148073
rect 307666 147999 307722 148008
rect 307576 147824 307628 147830
rect 307576 147766 307628 147772
rect 307680 147762 307708 147999
rect 307668 147756 307720 147762
rect 307668 147698 307720 147704
rect 307390 147656 307446 147665
rect 307390 147591 307446 147600
rect 307404 144226 307432 147591
rect 307666 146840 307722 146849
rect 307666 146775 307722 146784
rect 307680 146402 307708 146775
rect 307668 146396 307720 146402
rect 307668 146338 307720 146344
rect 307482 145888 307538 145897
rect 307482 145823 307538 145832
rect 307392 144220 307444 144226
rect 307392 144162 307444 144168
rect 307298 142080 307354 142089
rect 307298 142015 307354 142024
rect 307208 141432 307260 141438
rect 307208 141374 307260 141380
rect 307206 140448 307262 140457
rect 307206 140383 307262 140392
rect 307114 137048 307170 137057
rect 307114 136983 307170 136992
rect 307024 112464 307076 112470
rect 307024 112406 307076 112412
rect 306746 108896 306802 108905
rect 306746 108831 306802 108840
rect 306010 108488 306066 108497
rect 306010 108423 306066 108432
rect 305920 104848 305972 104854
rect 305920 104790 305972 104796
rect 305826 104272 305882 104281
rect 305826 104207 305882 104216
rect 305840 72486 305868 104207
rect 306024 76566 306052 108423
rect 306760 107778 306788 108831
rect 306748 107772 306800 107778
rect 306748 107714 306800 107720
rect 306562 105904 306618 105913
rect 306562 105839 306618 105848
rect 306576 104990 306604 105839
rect 306564 104984 306616 104990
rect 306564 104926 306616 104932
rect 306746 103456 306802 103465
rect 306746 103391 306802 103400
rect 306760 102270 306788 103391
rect 306930 102504 306986 102513
rect 306930 102439 306986 102448
rect 306748 102264 306800 102270
rect 306748 102206 306800 102212
rect 306944 102202 306972 102439
rect 306932 102196 306984 102202
rect 306932 102138 306984 102144
rect 306746 97880 306802 97889
rect 306746 97815 306802 97824
rect 306760 96762 306788 97815
rect 307022 97064 307078 97073
rect 307022 96999 307078 97008
rect 306748 96756 306800 96762
rect 306748 96698 306800 96704
rect 306012 76560 306064 76566
rect 306012 76502 306064 76508
rect 305828 72480 305880 72486
rect 305828 72422 305880 72428
rect 305736 35284 305788 35290
rect 305736 35226 305788 35232
rect 305644 17332 305696 17338
rect 305644 17274 305696 17280
rect 293224 8968 293276 8974
rect 293224 8910 293276 8916
rect 307036 4826 307064 96999
rect 307128 90370 307156 136983
rect 307220 119406 307248 140383
rect 307312 137290 307340 142015
rect 307390 141672 307446 141681
rect 307390 141607 307446 141616
rect 307404 139602 307432 141607
rect 307496 140894 307524 145823
rect 307574 145480 307630 145489
rect 307574 145415 307630 145424
rect 307588 144974 307616 145415
rect 307666 145072 307722 145081
rect 307666 145007 307668 145016
rect 307720 145007 307722 145016
rect 307668 144978 307720 144984
rect 307576 144968 307628 144974
rect 307576 144910 307628 144916
rect 307666 144256 307722 144265
rect 307666 144191 307722 144200
rect 307680 143614 307708 144191
rect 307668 143608 307720 143614
rect 307668 143550 307720 143556
rect 307666 143440 307722 143449
rect 307666 143375 307722 143384
rect 307680 142254 307708 143375
rect 307668 142248 307720 142254
rect 307668 142190 307720 142196
rect 307666 141264 307722 141273
rect 307666 141199 307722 141208
rect 307484 140888 307536 140894
rect 307484 140830 307536 140836
rect 307680 140826 307708 141199
rect 307668 140820 307720 140826
rect 307668 140762 307720 140768
rect 307574 140040 307630 140049
rect 307574 139975 307630 139984
rect 307392 139596 307444 139602
rect 307392 139538 307444 139544
rect 307588 139534 307616 139975
rect 307666 139632 307722 139641
rect 307666 139567 307722 139576
rect 307576 139528 307628 139534
rect 307576 139470 307628 139476
rect 307680 139466 307708 139567
rect 307668 139460 307720 139466
rect 307668 139402 307720 139408
rect 307482 139088 307538 139097
rect 307482 139023 307538 139032
rect 307496 138038 307524 139023
rect 307574 138680 307630 138689
rect 307574 138615 307630 138624
rect 307588 138106 307616 138615
rect 307666 138272 307722 138281
rect 307666 138207 307722 138216
rect 307680 138174 307708 138207
rect 307668 138168 307720 138174
rect 307668 138110 307720 138116
rect 307576 138100 307628 138106
rect 307576 138042 307628 138048
rect 307484 138032 307536 138038
rect 307484 137974 307536 137980
rect 307482 137456 307538 137465
rect 307482 137391 307538 137400
rect 307300 137284 307352 137290
rect 307300 137226 307352 137232
rect 307496 136746 307524 137391
rect 307484 136740 307536 136746
rect 307484 136682 307536 136688
rect 307390 136640 307446 136649
rect 307390 136575 307446 136584
rect 307404 135386 307432 136575
rect 307666 136232 307722 136241
rect 307666 136167 307722 136176
rect 307482 135688 307538 135697
rect 307482 135623 307538 135632
rect 307392 135380 307444 135386
rect 307392 135322 307444 135328
rect 307496 135318 307524 135623
rect 307576 135516 307628 135522
rect 307576 135458 307628 135464
rect 307484 135312 307536 135318
rect 307588 135289 307616 135458
rect 307680 135454 307708 136167
rect 307668 135448 307720 135454
rect 307668 135390 307720 135396
rect 307484 135254 307536 135260
rect 307574 135280 307630 135289
rect 307574 135215 307630 135224
rect 307574 134464 307630 134473
rect 307574 134399 307630 134408
rect 307588 134026 307616 134399
rect 307668 134088 307720 134094
rect 307666 134056 307668 134065
rect 307720 134056 307722 134065
rect 307576 134020 307628 134026
rect 307666 133991 307722 134000
rect 307576 133962 307628 133968
rect 307666 133648 307722 133657
rect 307666 133583 307722 133592
rect 307482 133240 307538 133249
rect 307482 133175 307538 133184
rect 307496 132530 307524 133175
rect 307680 132598 307708 133583
rect 307668 132592 307720 132598
rect 307668 132534 307720 132540
rect 307484 132524 307536 132530
rect 307484 132466 307536 132472
rect 307482 132288 307538 132297
rect 307482 132223 307538 132232
rect 307496 131170 307524 132223
rect 307666 131880 307722 131889
rect 307666 131815 307722 131824
rect 307680 131238 307708 131815
rect 307668 131232 307720 131238
rect 307668 131174 307720 131180
rect 307484 131164 307536 131170
rect 307484 131106 307536 131112
rect 307666 129840 307722 129849
rect 307666 129775 307668 129784
rect 307720 129775 307722 129784
rect 307668 129746 307720 129752
rect 307482 129296 307538 129305
rect 307482 129231 307538 129240
rect 307496 128382 307524 129231
rect 307574 128888 307630 128897
rect 307574 128823 307630 128832
rect 307588 128450 307616 128823
rect 307668 128512 307720 128518
rect 307666 128480 307668 128489
rect 307720 128480 307722 128489
rect 307576 128444 307628 128450
rect 307666 128415 307722 128424
rect 307576 128386 307628 128392
rect 307484 128376 307536 128382
rect 307484 128318 307536 128324
rect 307482 128072 307538 128081
rect 307482 128007 307538 128016
rect 307496 127022 307524 128007
rect 307574 127664 307630 127673
rect 307574 127599 307630 127608
rect 307588 127090 307616 127599
rect 307666 127256 307722 127265
rect 307666 127191 307722 127200
rect 307680 127158 307708 127191
rect 307668 127152 307720 127158
rect 307668 127094 307720 127100
rect 307576 127084 307628 127090
rect 307576 127026 307628 127032
rect 307484 127016 307536 127022
rect 307484 126958 307536 126964
rect 307482 126848 307538 126857
rect 307482 126783 307538 126792
rect 307496 125662 307524 126783
rect 307666 126440 307722 126449
rect 307666 126375 307722 126384
rect 307680 125798 307708 126375
rect 307668 125792 307720 125798
rect 307668 125734 307720 125740
rect 307484 125656 307536 125662
rect 307484 125598 307536 125604
rect 307482 125080 307538 125089
rect 307482 125015 307538 125024
rect 307298 124672 307354 124681
rect 307298 124607 307354 124616
rect 307208 119400 307260 119406
rect 307208 119342 307260 119348
rect 307206 116240 307262 116249
rect 307206 116175 307262 116184
rect 307116 90364 307168 90370
rect 307116 90306 307168 90312
rect 307220 71058 307248 116175
rect 307312 91798 307340 124607
rect 307496 124302 307524 125015
rect 307484 124296 307536 124302
rect 307484 124238 307536 124244
rect 307666 124264 307722 124273
rect 307666 124199 307668 124208
rect 307720 124199 307722 124208
rect 307668 124170 307720 124176
rect 307574 123448 307630 123457
rect 307574 123383 307630 123392
rect 307588 122942 307616 123383
rect 307666 123040 307722 123049
rect 307666 122975 307668 122984
rect 307720 122975 307722 122984
rect 307668 122946 307720 122952
rect 307576 122936 307628 122942
rect 307576 122878 307628 122884
rect 307482 122496 307538 122505
rect 307482 122431 307538 122440
rect 307496 121514 307524 122431
rect 307574 122088 307630 122097
rect 307574 122023 307630 122032
rect 307588 121582 307616 122023
rect 307666 121680 307722 121689
rect 307666 121615 307668 121624
rect 307720 121615 307722 121624
rect 307668 121586 307720 121592
rect 307576 121576 307628 121582
rect 307576 121518 307628 121524
rect 307484 121508 307536 121514
rect 307484 121450 307536 121456
rect 307482 121272 307538 121281
rect 307482 121207 307538 121216
rect 307496 120222 307524 121207
rect 307574 120864 307630 120873
rect 307574 120799 307630 120808
rect 307484 120216 307536 120222
rect 307484 120158 307536 120164
rect 307588 120154 307616 120799
rect 307666 120456 307722 120465
rect 307666 120391 307722 120400
rect 307680 120290 307708 120391
rect 307668 120284 307720 120290
rect 307668 120226 307720 120232
rect 307576 120148 307628 120154
rect 307576 120090 307628 120096
rect 307574 119640 307630 119649
rect 307574 119575 307630 119584
rect 307588 118969 307616 119575
rect 307666 119096 307722 119105
rect 307666 119031 307722 119040
rect 307574 118960 307630 118969
rect 307574 118895 307630 118904
rect 307680 118794 307708 119031
rect 307668 118788 307720 118794
rect 307668 118730 307720 118736
rect 307482 118688 307538 118697
rect 307482 118623 307538 118632
rect 307496 117366 307524 118623
rect 307574 117872 307630 117881
rect 307574 117807 307630 117816
rect 307588 117502 307616 117807
rect 307576 117496 307628 117502
rect 307576 117438 307628 117444
rect 307666 117464 307722 117473
rect 307666 117399 307668 117408
rect 307720 117399 307722 117408
rect 307668 117370 307720 117376
rect 307484 117360 307536 117366
rect 307484 117302 307536 117308
rect 307666 117056 307722 117065
rect 307666 116991 307722 117000
rect 307680 116074 307708 116991
rect 307668 116068 307720 116074
rect 307668 116010 307720 116016
rect 307666 114880 307722 114889
rect 307666 114815 307722 114824
rect 307680 114646 307708 114815
rect 307668 114640 307720 114646
rect 307668 114582 307720 114588
rect 307574 113656 307630 113665
rect 307574 113591 307630 113600
rect 307588 113286 307616 113591
rect 307576 113280 307628 113286
rect 307576 113222 307628 113228
rect 307666 113248 307722 113257
rect 307666 113183 307668 113192
rect 307720 113183 307722 113192
rect 307668 113154 307720 113160
rect 307574 112296 307630 112305
rect 307574 112231 307630 112240
rect 307588 111926 307616 112231
rect 307576 111920 307628 111926
rect 307576 111862 307628 111868
rect 307666 111888 307722 111897
rect 307666 111823 307668 111832
rect 307720 111823 307722 111832
rect 307668 111794 307720 111800
rect 307482 111480 307538 111489
rect 307482 111415 307538 111424
rect 307496 110498 307524 111415
rect 307574 111072 307630 111081
rect 307574 111007 307630 111016
rect 307588 110634 307616 111007
rect 307666 110664 307722 110673
rect 307576 110628 307628 110634
rect 307666 110599 307722 110608
rect 307576 110570 307628 110576
rect 307680 110566 307708 110599
rect 307668 110560 307720 110566
rect 307668 110502 307720 110508
rect 307484 110492 307536 110498
rect 307484 110434 307536 110440
rect 307482 110256 307538 110265
rect 307482 110191 307538 110200
rect 307496 109206 307524 110191
rect 307574 109848 307630 109857
rect 307574 109783 307630 109792
rect 307484 109200 307536 109206
rect 307484 109142 307536 109148
rect 307588 109138 307616 109783
rect 307666 109304 307722 109313
rect 307666 109239 307722 109248
rect 307576 109132 307628 109138
rect 307576 109074 307628 109080
rect 307680 109070 307708 109239
rect 307668 109064 307720 109070
rect 307668 109006 307720 109012
rect 307574 108080 307630 108089
rect 307574 108015 307630 108024
rect 307588 107710 307616 108015
rect 307668 107908 307720 107914
rect 307668 107850 307720 107856
rect 307576 107704 307628 107710
rect 307680 107681 307708 107850
rect 307576 107646 307628 107652
rect 307666 107672 307722 107681
rect 307666 107607 307722 107616
rect 307482 107264 307538 107273
rect 307482 107199 307538 107208
rect 307496 106486 307524 107199
rect 307574 106856 307630 106865
rect 307574 106791 307630 106800
rect 307484 106480 307536 106486
rect 307484 106422 307536 106428
rect 307588 106418 307616 106791
rect 307666 106448 307722 106457
rect 307576 106412 307628 106418
rect 307666 106383 307722 106392
rect 307576 106354 307628 106360
rect 307680 106350 307708 106383
rect 307668 106344 307720 106350
rect 307668 106286 307720 106292
rect 307666 105088 307722 105097
rect 307666 105023 307668 105032
rect 307720 105023 307722 105032
rect 307668 104994 307720 105000
rect 307574 104680 307630 104689
rect 307574 104615 307630 104624
rect 307588 103630 307616 104615
rect 307666 103864 307722 103873
rect 307666 103799 307722 103808
rect 307680 103698 307708 103799
rect 307668 103692 307720 103698
rect 307668 103634 307720 103640
rect 307576 103624 307628 103630
rect 307576 103566 307628 103572
rect 307482 103048 307538 103057
rect 307482 102983 307538 102992
rect 307496 102338 307524 102983
rect 307484 102332 307536 102338
rect 307484 102274 307536 102280
rect 307574 102096 307630 102105
rect 307574 102031 307630 102040
rect 307482 101688 307538 101697
rect 307482 101623 307538 101632
rect 307496 100774 307524 101623
rect 307588 100910 307616 102031
rect 307576 100904 307628 100910
rect 307576 100846 307628 100852
rect 307666 100872 307722 100881
rect 307666 100807 307668 100816
rect 307720 100807 307722 100816
rect 307668 100778 307720 100784
rect 307484 100768 307536 100774
rect 307484 100710 307536 100716
rect 307482 100464 307538 100473
rect 307482 100399 307538 100408
rect 307496 99482 307524 100399
rect 307666 100056 307722 100065
rect 307666 99991 307722 100000
rect 307484 99476 307536 99482
rect 307484 99418 307536 99424
rect 307680 99414 307708 99991
rect 307668 99408 307720 99414
rect 307668 99350 307720 99356
rect 307482 99104 307538 99113
rect 307482 99039 307538 99048
rect 307496 98122 307524 99039
rect 307666 98696 307722 98705
rect 307666 98631 307722 98640
rect 307574 98288 307630 98297
rect 307574 98223 307630 98232
rect 307484 98116 307536 98122
rect 307484 98058 307536 98064
rect 307588 98054 307616 98223
rect 307680 98190 307708 98631
rect 307668 98184 307720 98190
rect 307668 98126 307720 98132
rect 307576 98048 307628 98054
rect 307576 97990 307628 97996
rect 307482 97472 307538 97481
rect 307482 97407 307538 97416
rect 307496 96694 307524 97407
rect 307484 96688 307536 96694
rect 307484 96630 307536 96636
rect 307666 96248 307722 96257
rect 307666 96183 307722 96192
rect 307680 95266 307708 96183
rect 307668 95260 307720 95266
rect 307668 95202 307720 95208
rect 308416 94994 308444 299542
rect 308496 294160 308548 294166
rect 308496 294102 308548 294108
rect 308508 95985 308536 294102
rect 318064 292732 318116 292738
rect 318064 292674 318116 292680
rect 313924 288448 313976 288454
rect 313924 288390 313976 288396
rect 311164 267776 311216 267782
rect 311164 267718 311216 267724
rect 308588 265056 308640 265062
rect 308588 264998 308640 265004
rect 308494 95976 308550 95985
rect 308494 95911 308550 95920
rect 308600 95130 308628 264998
rect 309784 248464 309836 248470
rect 309784 248406 309836 248412
rect 308588 95124 308640 95130
rect 308588 95066 308640 95072
rect 309796 95062 309824 248406
rect 309876 225616 309928 225622
rect 309876 225558 309928 225564
rect 309888 176662 309916 225558
rect 311176 178770 311204 267718
rect 311256 242956 311308 242962
rect 311256 242898 311308 242904
rect 311164 178764 311216 178770
rect 311164 178706 311216 178712
rect 311268 177478 311296 242898
rect 312544 222896 312596 222902
rect 312544 222838 312596 222844
rect 311256 177472 311308 177478
rect 311256 177414 311308 177420
rect 309876 176656 309928 176662
rect 309876 176598 309928 176604
rect 312556 175953 312584 222838
rect 313936 177313 313964 288390
rect 315304 225684 315356 225690
rect 315304 225626 315356 225632
rect 314016 216028 314068 216034
rect 314016 215970 314068 215976
rect 314028 177614 314056 215970
rect 314016 177608 314068 177614
rect 314016 177550 314068 177556
rect 313922 177304 313978 177313
rect 313922 177239 313978 177248
rect 315316 176050 315344 225626
rect 318076 177546 318104 292674
rect 318156 278792 318208 278798
rect 318156 278734 318208 278740
rect 318064 177540 318116 177546
rect 318064 177482 318116 177488
rect 316038 176760 316094 176769
rect 316038 176695 316094 176704
rect 315304 176044 315356 176050
rect 315304 175986 315356 175992
rect 312542 175944 312598 175953
rect 316052 175930 316080 176695
rect 316020 175902 316080 175930
rect 312542 175879 312598 175888
rect 318168 175642 318196 278734
rect 318248 217320 318300 217326
rect 318248 217262 318300 217268
rect 318260 175982 318288 217262
rect 319456 176633 319484 300834
rect 333980 298240 334032 298246
rect 333980 298182 334032 298188
rect 325792 296744 325844 296750
rect 325792 296686 325844 296692
rect 320180 292664 320232 292670
rect 320180 292606 320232 292612
rect 320192 176769 320220 292606
rect 325698 290592 325754 290601
rect 325698 290527 325754 290536
rect 323676 253972 323728 253978
rect 323676 253914 323728 253920
rect 323584 244316 323636 244322
rect 323584 244258 323636 244264
rect 321652 228404 321704 228410
rect 321652 228346 321704 228352
rect 321560 200796 321612 200802
rect 321560 200738 321612 200744
rect 321284 184204 321336 184210
rect 321284 184146 321336 184152
rect 320178 176760 320234 176769
rect 320178 176695 320234 176704
rect 319442 176624 319498 176633
rect 319442 176559 319498 176568
rect 318248 175976 318300 175982
rect 318248 175918 318300 175924
rect 318156 175636 318208 175642
rect 318156 175578 318208 175584
rect 321296 165073 321324 184146
rect 321376 177336 321428 177342
rect 321376 177278 321428 177284
rect 321388 173777 321416 177278
rect 321468 176656 321520 176662
rect 321468 176598 321520 176604
rect 321480 176089 321508 176598
rect 321466 176080 321522 176089
rect 321466 176015 321522 176024
rect 321468 175636 321520 175642
rect 321468 175578 321520 175584
rect 321480 175273 321508 175578
rect 321466 175264 321522 175273
rect 321466 175199 321522 175208
rect 321374 173768 321430 173777
rect 321374 173703 321430 173712
rect 321282 165064 321338 165073
rect 321282 164999 321338 165008
rect 321572 106049 321600 200738
rect 321664 165753 321692 228346
rect 321836 185700 321888 185706
rect 321836 185642 321888 185648
rect 321848 172689 321876 185642
rect 322940 185632 322992 185638
rect 322940 185574 322992 185580
rect 321928 182980 321980 182986
rect 321928 182922 321980 182928
rect 321834 172680 321890 172689
rect 321834 172615 321890 172624
rect 321650 165744 321706 165753
rect 321650 165679 321706 165688
rect 321940 161474 321968 182922
rect 321756 161446 321968 161474
rect 321756 151337 321784 161446
rect 322952 153241 322980 185574
rect 322938 153232 322994 153241
rect 322938 153167 322994 153176
rect 321742 151328 321798 151337
rect 321742 151263 321798 151272
rect 323596 124098 323624 244258
rect 323688 141710 323716 253914
rect 324412 232552 324464 232558
rect 324412 232494 324464 232500
rect 324320 169720 324372 169726
rect 324320 169662 324372 169668
rect 324332 169425 324360 169662
rect 324318 169416 324374 169425
rect 324318 169351 324374 169360
rect 324424 168609 324452 232494
rect 324596 209092 324648 209098
rect 324596 209034 324648 209040
rect 324504 195356 324556 195362
rect 324504 195298 324556 195304
rect 324410 168600 324466 168609
rect 324410 168535 324466 168544
rect 324412 168360 324464 168366
rect 324412 168302 324464 168308
rect 324320 168292 324372 168298
rect 324320 168234 324372 168240
rect 324332 167793 324360 168234
rect 324318 167784 324374 167793
rect 324318 167719 324374 167728
rect 324424 167113 324452 168302
rect 324410 167104 324466 167113
rect 324410 167039 324466 167048
rect 324320 167000 324372 167006
rect 324320 166942 324372 166948
rect 324332 166297 324360 166942
rect 324318 166288 324374 166297
rect 324318 166223 324374 166232
rect 324412 164212 324464 164218
rect 324412 164154 324464 164160
rect 324320 164144 324372 164150
rect 324320 164086 324372 164092
rect 324332 163985 324360 164086
rect 324318 163976 324374 163985
rect 324318 163911 324374 163920
rect 324424 163169 324452 164154
rect 324410 163160 324466 163169
rect 324410 163095 324466 163104
rect 324320 162852 324372 162858
rect 324320 162794 324372 162800
rect 324332 162489 324360 162794
rect 324412 162784 324464 162790
rect 324412 162726 324464 162732
rect 324318 162480 324374 162489
rect 324318 162415 324374 162424
rect 324424 161673 324452 162726
rect 324410 161664 324466 161673
rect 324410 161599 324466 161608
rect 324320 161356 324372 161362
rect 324320 161298 324372 161304
rect 324332 160177 324360 161298
rect 324318 160168 324374 160177
rect 324318 160103 324374 160112
rect 324320 160064 324372 160070
rect 324320 160006 324372 160012
rect 324332 159361 324360 160006
rect 324318 159352 324374 159361
rect 324318 159287 324374 159296
rect 324412 158704 324464 158710
rect 324412 158646 324464 158652
rect 324320 158636 324372 158642
rect 324320 158578 324372 158584
rect 324332 158545 324360 158578
rect 324318 158536 324374 158545
rect 324318 158471 324374 158480
rect 324424 157865 324452 158646
rect 324410 157856 324466 157865
rect 324410 157791 324466 157800
rect 324320 157344 324372 157350
rect 324320 157286 324372 157292
rect 324332 157049 324360 157286
rect 324412 157276 324464 157282
rect 324412 157218 324464 157224
rect 324318 157040 324374 157049
rect 324318 156975 324374 156984
rect 324424 156369 324452 157218
rect 324410 156360 324466 156369
rect 324410 156295 324466 156304
rect 324320 155916 324372 155922
rect 324320 155858 324372 155864
rect 324332 155553 324360 155858
rect 324318 155544 324374 155553
rect 324318 155479 324374 155488
rect 324516 154737 324544 195298
rect 324502 154728 324558 154737
rect 324502 154663 324558 154672
rect 324320 154556 324372 154562
rect 324320 154498 324372 154504
rect 324332 154057 324360 154498
rect 324318 154048 324374 154057
rect 324318 153983 324374 153992
rect 324320 153196 324372 153202
rect 324320 153138 324372 153144
rect 324332 152425 324360 153138
rect 324318 152416 324374 152425
rect 324318 152351 324374 152360
rect 324320 151768 324372 151774
rect 324318 151736 324320 151745
rect 324372 151736 324374 151745
rect 324318 151671 324374 151680
rect 324320 150408 324372 150414
rect 324320 150350 324372 150356
rect 324332 150113 324360 150350
rect 324412 150340 324464 150346
rect 324412 150282 324464 150288
rect 324318 150104 324374 150113
rect 324318 150039 324374 150048
rect 324424 149433 324452 150282
rect 324410 149424 324466 149433
rect 324410 149359 324466 149368
rect 324320 149048 324372 149054
rect 324320 148990 324372 148996
rect 324332 148617 324360 148990
rect 324412 148980 324464 148986
rect 324412 148922 324464 148928
rect 324318 148608 324374 148617
rect 324318 148543 324374 148552
rect 324424 147801 324452 148922
rect 324410 147792 324466 147801
rect 324410 147727 324466 147736
rect 324320 147620 324372 147626
rect 324320 147562 324372 147568
rect 324332 147121 324360 147562
rect 324318 147112 324374 147121
rect 324318 147047 324374 147056
rect 324318 146296 324374 146305
rect 324318 146231 324374 146240
rect 324412 146260 324464 146266
rect 324332 146198 324360 146231
rect 324412 146202 324464 146208
rect 324320 146192 324372 146198
rect 324320 146134 324372 146140
rect 324424 145489 324452 146202
rect 324410 145480 324466 145489
rect 324410 145415 324466 145424
rect 324320 144900 324372 144906
rect 324320 144842 324372 144848
rect 324332 144809 324360 144842
rect 324412 144832 324464 144838
rect 324318 144800 324374 144809
rect 324412 144774 324464 144780
rect 324318 144735 324374 144744
rect 324424 143993 324452 144774
rect 324410 143984 324466 143993
rect 324410 143919 324466 143928
rect 324320 142724 324372 142730
rect 324320 142666 324372 142672
rect 324332 142497 324360 142666
rect 324318 142488 324374 142497
rect 324318 142423 324374 142432
rect 324320 142112 324372 142118
rect 324320 142054 324372 142060
rect 323676 141704 323728 141710
rect 324332 141681 324360 142054
rect 324504 142044 324556 142050
rect 324504 141986 324556 141992
rect 324412 141704 324464 141710
rect 323676 141646 323728 141652
rect 324318 141672 324374 141681
rect 324412 141646 324464 141652
rect 324318 141607 324374 141616
rect 324320 139392 324372 139398
rect 324318 139360 324320 139369
rect 324372 139360 324374 139369
rect 324318 139295 324374 139304
rect 324320 137964 324372 137970
rect 324320 137906 324372 137912
rect 324332 137873 324360 137906
rect 324318 137864 324374 137873
rect 324318 137799 324374 137808
rect 324320 136536 324372 136542
rect 324320 136478 324372 136484
rect 324332 136377 324360 136478
rect 324318 136368 324374 136377
rect 324318 136303 324374 136312
rect 324320 133884 324372 133890
rect 324320 133826 324372 133832
rect 324332 133249 324360 133826
rect 324318 133240 324374 133249
rect 324318 133175 324374 133184
rect 324318 132424 324374 132433
rect 324318 132359 324320 132368
rect 324372 132359 324374 132368
rect 324320 132330 324372 132336
rect 324424 131186 324452 141646
rect 324516 140865 324544 141986
rect 324502 140856 324558 140865
rect 324502 140791 324558 140800
rect 324504 139324 324556 139330
rect 324504 139266 324556 139272
rect 324516 138553 324544 139266
rect 324502 138544 324558 138553
rect 324502 138479 324558 138488
rect 324504 137896 324556 137902
rect 324504 137838 324556 137844
rect 324516 137057 324544 137838
rect 324502 137048 324558 137057
rect 324502 136983 324558 136992
rect 324504 136604 324556 136610
rect 324504 136546 324556 136552
rect 324516 135561 324544 136546
rect 324502 135552 324558 135561
rect 324502 135487 324558 135496
rect 324504 132456 324556 132462
rect 324504 132398 324556 132404
rect 324516 131753 324544 132398
rect 324502 131744 324558 131753
rect 324502 131679 324558 131688
rect 324424 131158 324544 131186
rect 324320 131096 324372 131102
rect 324320 131038 324372 131044
rect 324332 130937 324360 131038
rect 324412 131028 324464 131034
rect 324412 130970 324464 130976
rect 324318 130928 324374 130937
rect 324318 130863 324374 130872
rect 324424 130121 324452 130970
rect 324410 130112 324466 130121
rect 324410 130047 324466 130056
rect 324320 129736 324372 129742
rect 324320 129678 324372 129684
rect 324332 128625 324360 129678
rect 324318 128616 324374 128625
rect 324318 128551 324374 128560
rect 324320 128308 324372 128314
rect 324320 128250 324372 128256
rect 324332 127809 324360 128250
rect 324318 127800 324374 127809
rect 324318 127735 324374 127744
rect 324320 126948 324372 126954
rect 324320 126890 324372 126896
rect 324332 126313 324360 126890
rect 324318 126304 324374 126313
rect 324318 126239 324374 126248
rect 324516 125497 324544 131158
rect 324502 125488 324558 125497
rect 324502 125423 324558 125432
rect 324320 124160 324372 124166
rect 324320 124102 324372 124108
rect 323584 124092 323636 124098
rect 323584 124034 323636 124040
rect 324332 124001 324360 124102
rect 324504 124092 324556 124098
rect 324504 124034 324556 124040
rect 324318 123992 324374 124001
rect 324318 123927 324374 123936
rect 324320 122732 324372 122738
rect 324320 122674 324372 122680
rect 324332 121689 324360 122674
rect 324318 121680 324374 121689
rect 324318 121615 324374 121624
rect 324412 121440 324464 121446
rect 324412 121382 324464 121388
rect 324320 121372 324372 121378
rect 324320 121314 324372 121320
rect 324332 120873 324360 121314
rect 324318 120864 324374 120873
rect 324318 120799 324374 120808
rect 324424 120193 324452 121382
rect 324410 120184 324466 120193
rect 324410 120119 324466 120128
rect 324516 119377 324544 124034
rect 324502 119368 324558 119377
rect 324502 119303 324558 119312
rect 324412 118652 324464 118658
rect 324412 118594 324464 118600
rect 324320 118584 324372 118590
rect 324318 118552 324320 118561
rect 324372 118552 324374 118561
rect 324318 118487 324374 118496
rect 324424 117881 324452 118594
rect 324410 117872 324466 117881
rect 324410 117807 324466 117816
rect 324412 117292 324464 117298
rect 324412 117234 324464 117240
rect 324320 117224 324372 117230
rect 324320 117166 324372 117172
rect 324332 117065 324360 117166
rect 324318 117056 324374 117065
rect 324318 116991 324374 117000
rect 324424 116385 324452 117234
rect 324410 116376 324466 116385
rect 324410 116311 324466 116320
rect 324320 115932 324372 115938
rect 324320 115874 324372 115880
rect 324332 115569 324360 115874
rect 324318 115560 324374 115569
rect 324318 115495 324374 115504
rect 324320 114504 324372 114510
rect 324320 114446 324372 114452
rect 324332 114073 324360 114446
rect 324412 114436 324464 114442
rect 324412 114378 324464 114384
rect 324318 114064 324374 114073
rect 324318 113999 324374 114008
rect 324424 113257 324452 114378
rect 324410 113248 324466 113257
rect 324410 113183 324466 113192
rect 324320 113144 324372 113150
rect 324320 113086 324372 113092
rect 324332 112441 324360 113086
rect 324318 112432 324374 112441
rect 324318 112367 324374 112376
rect 324320 111784 324372 111790
rect 324318 111752 324320 111761
rect 324372 111752 324374 111761
rect 324318 111687 324374 111696
rect 324410 108624 324466 108633
rect 324410 108559 324466 108568
rect 324320 108044 324372 108050
rect 324320 107986 324372 107992
rect 324332 107817 324360 107986
rect 324318 107808 324374 107817
rect 324318 107743 324374 107752
rect 323490 106584 323546 106593
rect 323490 106519 323546 106528
rect 323504 106321 323532 106519
rect 323490 106312 323546 106321
rect 323490 106247 323546 106256
rect 321558 106040 321614 106049
rect 321558 105975 321614 105984
rect 324318 103184 324374 103193
rect 324318 103119 324374 103128
rect 321742 98152 321798 98161
rect 321742 98087 321798 98096
rect 321558 97336 321614 97345
rect 321558 97271 321614 97280
rect 321466 96656 321522 96665
rect 321466 96591 321468 96600
rect 321520 96591 321522 96600
rect 321468 96562 321520 96568
rect 321572 95130 321600 97271
rect 321650 96656 321706 96665
rect 321650 96591 321706 96600
rect 321664 95169 321692 96591
rect 321650 95160 321706 95169
rect 321560 95124 321612 95130
rect 321650 95095 321706 95104
rect 321560 95066 321612 95072
rect 309784 95056 309836 95062
rect 309784 94998 309836 95004
rect 321756 94994 321784 98087
rect 324332 95198 324360 103119
rect 324320 95192 324372 95198
rect 324320 95134 324372 95140
rect 324424 95062 324452 108559
rect 324608 100881 324636 209034
rect 324688 161424 324740 161430
rect 324688 161366 324740 161372
rect 324700 160857 324728 161366
rect 324686 160848 324742 160857
rect 324686 160783 324742 160792
rect 324686 142760 324742 142769
rect 324686 142695 324742 142704
rect 324700 140185 324728 142695
rect 324686 140176 324742 140185
rect 324686 140111 324742 140120
rect 324964 139256 325016 139262
rect 324964 139198 325016 139204
rect 324976 123185 325004 139198
rect 325606 124808 325662 124817
rect 325712 124794 325740 290527
rect 325804 134065 325832 296686
rect 327080 286340 327132 286346
rect 327080 286282 327132 286288
rect 325882 176624 325938 176633
rect 325882 176559 325938 176568
rect 325896 171737 325924 176559
rect 325882 171728 325938 171737
rect 325882 171663 325938 171672
rect 327092 142730 327120 286282
rect 328460 277500 328512 277506
rect 328460 277442 328512 277448
rect 327172 262268 327224 262274
rect 327172 262210 327224 262216
rect 327080 142724 327132 142730
rect 327080 142666 327132 142672
rect 327184 139262 327212 262210
rect 327356 235340 327408 235346
rect 327356 235282 327408 235288
rect 327264 203584 327316 203590
rect 327264 203526 327316 203532
rect 327172 139256 327224 139262
rect 327172 139198 327224 139204
rect 325790 134056 325846 134065
rect 325790 133991 325846 134000
rect 325662 124766 325740 124794
rect 325606 124743 325662 124752
rect 324962 123176 325018 123185
rect 324962 123111 325018 123120
rect 324688 122800 324740 122806
rect 324688 122742 324740 122748
rect 324700 122505 324728 122742
rect 324686 122496 324742 122505
rect 324686 122431 324742 122440
rect 327276 108050 327304 203526
rect 327368 151774 327396 235282
rect 327356 151768 327408 151774
rect 327356 151710 327408 151716
rect 328472 126954 328500 277442
rect 331220 276072 331272 276078
rect 331220 276014 331272 276020
rect 328552 240236 328604 240242
rect 328552 240178 328604 240184
rect 328564 133890 328592 240178
rect 330116 240168 330168 240174
rect 330116 240110 330168 240116
rect 329932 222964 329984 222970
rect 329932 222906 329984 222912
rect 328644 188352 328696 188358
rect 328644 188294 328696 188300
rect 328656 154562 328684 188294
rect 328736 178696 328788 178702
rect 328736 178638 328788 178644
rect 328748 160070 328776 178638
rect 328736 160064 328788 160070
rect 328736 160006 328788 160012
rect 328644 154556 328696 154562
rect 328644 154498 328696 154504
rect 328552 133884 328604 133890
rect 328552 133826 328604 133832
rect 329944 128314 329972 222906
rect 330024 214600 330076 214606
rect 330024 214542 330076 214548
rect 330036 137902 330064 214542
rect 330024 137896 330076 137902
rect 330024 137838 330076 137844
rect 330128 129742 330156 240110
rect 331232 144838 331260 276014
rect 332876 257372 332928 257378
rect 332876 257314 332928 257320
rect 331312 250504 331364 250510
rect 331312 250446 331364 250452
rect 331220 144832 331272 144838
rect 331220 144774 331272 144780
rect 331324 131102 331352 250446
rect 331404 231124 331456 231130
rect 331404 231066 331456 231072
rect 331312 131096 331364 131102
rect 331312 131038 331364 131044
rect 331416 131034 331444 231066
rect 332784 183048 332836 183054
rect 332784 182990 332836 182996
rect 332692 181552 332744 181558
rect 332692 181494 332744 181500
rect 331496 177472 331548 177478
rect 331496 177414 331548 177420
rect 331508 162790 331536 177414
rect 332600 176044 332652 176050
rect 332600 175986 332652 175992
rect 332612 169726 332640 175986
rect 332600 169720 332652 169726
rect 332600 169662 332652 169668
rect 331496 162784 331548 162790
rect 331496 162726 331548 162732
rect 331404 131028 331456 131034
rect 331404 130970 331456 130976
rect 330116 129736 330168 129742
rect 330116 129678 330168 129684
rect 329932 128308 329984 128314
rect 329932 128250 329984 128256
rect 328460 126948 328512 126954
rect 328460 126890 328512 126896
rect 332704 117230 332732 181494
rect 332796 139330 332824 182990
rect 332888 158642 332916 257314
rect 332876 158636 332928 158642
rect 332876 158578 332928 158584
rect 333992 142050 334020 298182
rect 339500 296880 339552 296886
rect 339500 296822 339552 296828
rect 336740 292596 336792 292602
rect 336740 292538 336792 292544
rect 335360 284368 335412 284374
rect 335360 284310 335412 284316
rect 334256 220108 334308 220114
rect 334256 220050 334308 220056
rect 334164 199504 334216 199510
rect 334164 199446 334216 199452
rect 334072 177608 334124 177614
rect 334072 177550 334124 177556
rect 333980 142044 334032 142050
rect 333980 141986 334032 141992
rect 332784 139324 332836 139330
rect 332784 139266 332836 139272
rect 332692 117224 332744 117230
rect 332692 117166 332744 117172
rect 334084 114442 334112 177550
rect 334176 146198 334204 199446
rect 334268 168298 334296 220050
rect 334256 168292 334308 168298
rect 334256 168234 334308 168240
rect 335372 161362 335400 284310
rect 335544 180328 335596 180334
rect 335544 180270 335596 180276
rect 335452 178764 335504 178770
rect 335452 178706 335504 178712
rect 335360 161356 335412 161362
rect 335360 161298 335412 161304
rect 334164 146192 334216 146198
rect 334164 146134 334216 146140
rect 334072 114436 334124 114442
rect 334072 114378 334124 114384
rect 335464 113150 335492 178706
rect 335556 121378 335584 180270
rect 335636 175976 335688 175982
rect 335636 175918 335688 175924
rect 335648 164150 335676 175918
rect 335636 164144 335688 164150
rect 335636 164086 335688 164092
rect 336752 162858 336780 292538
rect 338120 238060 338172 238066
rect 338120 238002 338172 238008
rect 336832 195288 336884 195294
rect 336832 195230 336884 195236
rect 336740 162852 336792 162858
rect 336740 162794 336792 162800
rect 335544 121372 335596 121378
rect 335544 121314 335596 121320
rect 336844 115938 336872 195230
rect 337016 192500 337068 192506
rect 337016 192442 337068 192448
rect 336924 180260 336976 180266
rect 336924 180202 336976 180208
rect 336936 117298 336964 180202
rect 337028 148986 337056 192442
rect 337016 148980 337068 148986
rect 337016 148922 337068 148928
rect 338132 122738 338160 238002
rect 338212 186992 338264 186998
rect 338212 186934 338264 186940
rect 338224 146266 338252 186934
rect 338396 182912 338448 182918
rect 338396 182854 338448 182860
rect 338304 177540 338356 177546
rect 338304 177482 338356 177488
rect 338316 158710 338344 177482
rect 338408 168366 338436 182854
rect 338396 168360 338448 168366
rect 338396 168302 338448 168308
rect 338304 158704 338356 158710
rect 338304 158646 338356 158652
rect 338212 146260 338264 146266
rect 338212 146202 338264 146208
rect 338120 122732 338172 122738
rect 338120 122674 338172 122680
rect 339512 121446 339540 296822
rect 340880 296812 340932 296818
rect 340880 296754 340932 296760
rect 339592 202156 339644 202162
rect 339592 202098 339644 202104
rect 339500 121440 339552 121446
rect 339500 121382 339552 121388
rect 339604 118590 339632 202098
rect 339776 189780 339828 189786
rect 339776 189722 339828 189728
rect 339684 180192 339736 180198
rect 339684 180134 339736 180140
rect 339696 136542 339724 180134
rect 339788 161430 339816 189722
rect 339776 161424 339828 161430
rect 339776 161366 339828 161372
rect 340892 147626 340920 296754
rect 340972 243568 341024 243574
rect 340972 243510 341024 243516
rect 340984 242894 341012 243510
rect 340972 242888 341024 242894
rect 340972 242830 341024 242836
rect 340972 236700 341024 236706
rect 340972 236642 341024 236648
rect 340880 147620 340932 147626
rect 340880 147562 340932 147568
rect 339684 136536 339736 136542
rect 339684 136478 339736 136484
rect 339592 118584 339644 118590
rect 339592 118526 339644 118532
rect 336924 117292 336976 117298
rect 336924 117234 336976 117240
rect 336832 115932 336884 115938
rect 336832 115874 336884 115880
rect 340984 114510 341012 236642
rect 341064 213240 341116 213246
rect 341064 213182 341116 213188
rect 341076 118658 341104 213182
rect 341156 177404 341208 177410
rect 341156 177346 341208 177352
rect 341168 132394 341196 177346
rect 341156 132388 341208 132394
rect 341156 132330 341208 132336
rect 341064 118652 341116 118658
rect 341064 118594 341116 118600
rect 340972 114504 341024 114510
rect 340972 114446 341024 114452
rect 335452 113144 335504 113150
rect 335452 113086 335504 113092
rect 342272 111790 342300 306342
rect 343640 299532 343692 299538
rect 343640 299474 343692 299480
rect 342352 280220 342404 280226
rect 342352 280162 342404 280168
rect 342364 124166 342392 280162
rect 342444 260908 342496 260914
rect 342444 260850 342496 260856
rect 342456 137970 342484 260850
rect 342536 180124 342588 180130
rect 342536 180066 342588 180072
rect 342548 144906 342576 180066
rect 342536 144900 342588 144906
rect 342536 144842 342588 144848
rect 342444 137964 342496 137970
rect 342444 137906 342496 137912
rect 343652 136610 343680 299474
rect 347044 295384 347096 295390
rect 347044 295326 347096 295332
rect 345020 294092 345072 294098
rect 345020 294034 345072 294040
rect 343732 227044 343784 227050
rect 343732 226986 343784 226992
rect 343744 157282 343772 226986
rect 343824 181484 343876 181490
rect 343824 181426 343876 181432
rect 343732 157276 343784 157282
rect 343732 157218 343784 157224
rect 343640 136604 343692 136610
rect 343640 136546 343692 136552
rect 342352 124160 342404 124166
rect 342352 124102 342404 124108
rect 343836 122806 343864 181426
rect 345032 132462 345060 294034
rect 346398 292632 346454 292641
rect 346398 292567 346454 292576
rect 345112 291304 345164 291310
rect 345110 291272 345112 291281
rect 345164 291272 345166 291281
rect 345110 291207 345166 291216
rect 345112 266416 345164 266422
rect 345112 266358 345164 266364
rect 345124 149054 345152 266358
rect 345294 182880 345350 182889
rect 345204 182844 345256 182850
rect 345294 182815 345350 182824
rect 345204 182786 345256 182792
rect 345216 164218 345244 182786
rect 345308 167006 345336 182815
rect 345296 167000 345348 167006
rect 345296 166942 345348 166948
rect 345204 164212 345256 164218
rect 345204 164154 345256 164160
rect 346412 157350 346440 292567
rect 346492 251252 346544 251258
rect 346492 251194 346544 251200
rect 346400 157344 346452 157350
rect 346400 157286 346452 157292
rect 346504 150346 346532 251194
rect 346584 218748 346636 218754
rect 346584 218690 346636 218696
rect 346596 150414 346624 218690
rect 347056 179382 347084 295326
rect 350540 294024 350592 294030
rect 350540 293966 350592 293972
rect 347780 277432 347832 277438
rect 347780 277374 347832 277380
rect 347044 179376 347096 179382
rect 347044 179318 347096 179324
rect 347792 155922 347820 277374
rect 349160 264988 349212 264994
rect 349160 264930 349212 264936
rect 347872 252612 347924 252618
rect 347872 252554 347924 252560
rect 347780 155916 347832 155922
rect 347780 155858 347832 155864
rect 347884 153202 347912 252554
rect 347872 153196 347924 153202
rect 347872 153138 347924 153144
rect 346584 150408 346636 150414
rect 346584 150350 346636 150356
rect 346492 150340 346544 150346
rect 346492 150282 346544 150288
rect 345112 149048 345164 149054
rect 345112 148990 345164 148996
rect 349172 142118 349200 264930
rect 349160 142112 349212 142118
rect 349160 142054 349212 142060
rect 350552 139398 350580 293966
rect 392584 275324 392636 275330
rect 392584 275266 392636 275272
rect 350540 139392 350592 139398
rect 350540 139334 350592 139340
rect 345020 132456 345072 132462
rect 345020 132398 345072 132404
rect 392596 126954 392624 275266
rect 395344 272536 395396 272542
rect 395344 272478 395396 272484
rect 392584 126948 392636 126954
rect 392584 126890 392636 126896
rect 343824 122800 343876 122806
rect 343824 122742 343876 122748
rect 342260 111784 342312 111790
rect 342260 111726 342312 111732
rect 327264 108044 327316 108050
rect 327264 107986 327316 107992
rect 324594 100872 324650 100881
rect 324594 100807 324650 100816
rect 395356 100706 395384 272478
rect 494072 238746 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 527192 702642 527220 703520
rect 527180 702636 527232 702642
rect 527180 702578 527232 702584
rect 543476 702434 543504 703520
rect 559668 702574 559696 703520
rect 559656 702568 559708 702574
rect 559656 702510 559708 702516
rect 580908 702500 580960 702506
rect 580908 702442 580960 702448
rect 542372 702406 543504 702434
rect 494060 238740 494112 238746
rect 494060 238682 494112 238688
rect 542372 229090 542400 702406
rect 580920 697241 580948 702442
rect 580906 697232 580962 697241
rect 580906 697167 580962 697176
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 582378 591016 582434 591025
rect 582378 590951 582434 590960
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580262 511320 580318 511329
rect 580262 511255 580318 511264
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 580184 470626 580212 471407
rect 580172 470620 580224 470626
rect 580172 470562 580224 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 579894 431624 579950 431633
rect 579894 431559 579950 431568
rect 579908 430642 579936 431559
rect 579896 430636 579948 430642
rect 579896 430578 579948 430584
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 579618 365120 579674 365129
rect 579618 365055 579674 365064
rect 579632 364410 579660 365055
rect 579620 364404 579672 364410
rect 579620 364346 579672 364352
rect 580172 351960 580224 351966
rect 580170 351928 580172 351937
rect 580224 351928 580226 351937
rect 580170 351863 580226 351872
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 324358 580212 325207
rect 580172 324352 580224 324358
rect 580172 324294 580224 324300
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580184 311914 580212 312015
rect 580172 311908 580224 311914
rect 580172 311850 580224 311856
rect 580276 307086 580304 511255
rect 580264 307080 580316 307086
rect 580264 307022 580316 307028
rect 580264 282192 580316 282198
rect 580264 282134 580316 282140
rect 579620 259412 579672 259418
rect 579620 259354 579672 259360
rect 579632 258913 579660 259354
rect 579618 258904 579674 258913
rect 579618 258839 579674 258848
rect 579894 245576 579950 245585
rect 579894 245511 579950 245520
rect 579908 243574 579936 245511
rect 579896 243568 579948 243574
rect 579896 243510 579948 243516
rect 542360 229084 542412 229090
rect 542360 229026 542412 229032
rect 580172 206984 580224 206990
rect 580172 206926 580224 206932
rect 580184 205737 580212 206926
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 579988 179376 580040 179382
rect 579988 179318 580040 179324
rect 580000 179217 580028 179318
rect 579986 179208 580042 179217
rect 579986 179143 580042 179152
rect 580276 152697 580304 282134
rect 580354 279712 580410 279721
rect 580354 279647 580410 279656
rect 580368 219065 580396 279647
rect 580446 272232 580502 272241
rect 580446 272167 580502 272176
rect 580460 264217 580488 272167
rect 580446 264208 580502 264217
rect 580446 264143 580502 264152
rect 580448 247716 580500 247722
rect 580448 247658 580500 247664
rect 580460 232393 580488 247658
rect 582392 233238 582420 590951
rect 582470 537840 582526 537849
rect 582470 537775 582526 537784
rect 582484 238814 582512 537775
rect 582746 298752 582802 298761
rect 582746 298687 582802 298696
rect 582564 298172 582616 298178
rect 582564 298114 582616 298120
rect 582472 238808 582524 238814
rect 582472 238750 582524 238756
rect 582472 233912 582524 233918
rect 582472 233854 582524 233860
rect 582380 233232 582432 233238
rect 582380 233174 582432 233180
rect 580446 232384 580502 232393
rect 580446 232319 580502 232328
rect 582380 229764 582432 229770
rect 582380 229706 582432 229712
rect 580354 219056 580410 219065
rect 580354 218991 580410 219000
rect 580262 152688 580318 152697
rect 580262 152623 580318 152632
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 395344 100700 395396 100706
rect 395344 100642 395396 100648
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 324502 100192 324558 100201
rect 324502 100127 324558 100136
rect 324412 95056 324464 95062
rect 324412 94998 324464 95004
rect 308404 94988 308456 94994
rect 308404 94930 308456 94936
rect 321744 94988 321796 94994
rect 321744 94930 321796 94936
rect 324516 93770 324544 100127
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 324504 93764 324556 93770
rect 324504 93706 324556 93712
rect 307300 91792 307352 91798
rect 307300 91734 307352 91740
rect 307208 71052 307260 71058
rect 307208 70994 307260 71000
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 582392 6633 582420 229706
rect 582484 46345 582512 233854
rect 582470 46336 582526 46345
rect 582470 46271 582526 46280
rect 582576 19825 582604 298114
rect 582656 291236 582708 291242
rect 582656 291178 582708 291184
rect 582668 112849 582696 291178
rect 582760 237386 582788 298687
rect 582748 237380 582800 237386
rect 582748 237322 582800 237328
rect 582838 231160 582894 231169
rect 582838 231095 582894 231104
rect 582748 191140 582800 191146
rect 582748 191082 582800 191088
rect 582654 112840 582710 112849
rect 582654 112775 582710 112784
rect 582760 33153 582788 191082
rect 582852 86193 582880 231095
rect 582838 86184 582894 86193
rect 582838 86119 582894 86128
rect 582746 33144 582802 33153
rect 582746 33079 582802 33088
rect 582562 19816 582618 19825
rect 582562 19751 582618 19760
rect 582378 6624 582434 6633
rect 582378 6559 582434 6568
rect 307024 4820 307076 4826
rect 307024 4762 307076 4768
rect 290464 2168 290516 2174
rect 290464 2110 290516 2116
rect 250444 2100 250496 2106
rect 250444 2042 250496 2048
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 2778 606056 2834 606112
rect 3330 579944 3386 580000
rect 3238 566888 3294 566944
rect 3330 553832 3386 553888
rect 2962 527856 3018 527912
rect 3330 501744 3386 501800
rect 3054 475632 3110 475688
rect 3330 462576 3386 462632
rect 3330 449520 3386 449576
rect 3330 423544 3386 423600
rect 3330 410488 3386 410544
rect 3330 397468 3332 397488
rect 3332 397468 3384 397488
rect 3384 397468 3386 397488
rect 3330 397432 3386 397468
rect 3330 371320 3386 371376
rect 3330 358400 3386 358456
rect 3330 345344 3386 345400
rect 3514 671200 3570 671256
rect 3514 658144 3570 658200
rect 3514 632068 3516 632088
rect 3516 632068 3568 632088
rect 3568 632068 3570 632088
rect 3514 632032 3570 632068
rect 3514 619112 3570 619168
rect 3514 514800 3570 514856
rect 3330 319232 3386 319288
rect 3422 306176 3478 306232
rect 2778 293120 2834 293176
rect 3146 254088 3202 254144
rect 3054 241032 3110 241088
rect 3054 201864 3110 201920
rect 3514 267144 3570 267200
rect 3514 214956 3516 214976
rect 3516 214956 3568 214976
rect 3568 214956 3570 214976
rect 3514 214920 3570 214956
rect 3422 188808 3478 188864
rect 3238 162832 3294 162888
rect 3422 149776 3478 149832
rect 3238 136720 3294 136776
rect 3422 110608 3478 110664
rect 2778 97552 2834 97608
rect 3146 84632 3202 84688
rect 2778 61376 2834 61432
rect 3054 58520 3110 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3238 32408 3294 32464
rect 3514 19352 3570 19408
rect 3422 6432 3478 6488
rect 8298 57160 8354 57216
rect 11058 22616 11114 22672
rect 22098 46144 22154 46200
rect 28998 65456 29054 65512
rect 34518 69536 34574 69592
rect 46846 206216 46902 206272
rect 52366 197920 52422 197976
rect 54942 232464 54998 232520
rect 55034 208936 55090 208992
rect 49698 75112 49754 75168
rect 57794 207576 57850 207632
rect 61842 193840 61898 193896
rect 60646 184184 60702 184240
rect 64694 125568 64750 125624
rect 64694 94832 64750 94888
rect 59358 64096 59414 64152
rect 67454 285640 67510 285696
rect 67638 291080 67694 291136
rect 68834 296792 68890 296848
rect 68834 290400 68890 290456
rect 68742 289720 68798 289776
rect 68190 289040 68246 289096
rect 67638 287680 67694 287736
rect 67730 287000 67786 287056
rect 67638 286320 67694 286376
rect 67638 284316 67640 284336
rect 67640 284316 67692 284336
rect 67692 284316 67694 284336
rect 67638 284280 67694 284316
rect 67546 282920 67602 282976
rect 68834 283600 68890 283656
rect 68558 281560 68614 281616
rect 67638 280880 67694 280936
rect 68374 280200 68430 280256
rect 67638 279520 67694 279576
rect 67730 278160 67786 278216
rect 67638 277500 67694 277536
rect 67638 277480 67640 277500
rect 67640 277480 67692 277500
rect 67692 277480 67694 277500
rect 67730 276800 67786 276856
rect 67638 276120 67694 276176
rect 67730 275440 67786 275496
rect 67638 274780 67694 274816
rect 67638 274760 67640 274780
rect 67640 274760 67692 274780
rect 67692 274760 67694 274780
rect 67638 274080 67694 274136
rect 68006 273400 68062 273456
rect 67822 272720 67878 272776
rect 67638 272040 67694 272096
rect 67638 271360 67694 271416
rect 67730 270680 67786 270736
rect 67638 270000 67694 270056
rect 68282 269320 68338 269376
rect 67546 268640 67602 268696
rect 67362 261160 67418 261216
rect 67454 251640 67510 251696
rect 67638 267960 67694 268016
rect 67638 267280 67694 267336
rect 67730 266600 67786 266656
rect 67822 265920 67878 265976
rect 67638 265240 67694 265296
rect 67730 264560 67786 264616
rect 67638 263880 67694 263936
rect 67638 263200 67694 263256
rect 67638 262520 67694 262576
rect 67730 261840 67786 261896
rect 67638 260480 67694 260536
rect 67638 259800 67694 259856
rect 67730 259120 67786 259176
rect 67638 258440 67694 258496
rect 67730 257760 67786 257816
rect 67638 257080 67694 257136
rect 67638 256400 67694 256456
rect 67730 255720 67786 255776
rect 67638 255040 67694 255096
rect 67638 253680 67694 253736
rect 68098 253000 68154 253056
rect 67638 250960 67694 251016
rect 67730 250280 67786 250336
rect 67638 249600 67694 249656
rect 67638 248920 67694 248976
rect 67638 248240 67694 248296
rect 67730 247560 67786 247616
rect 67638 246880 67694 246936
rect 75366 302232 75422 302288
rect 80518 299512 80574 299568
rect 80334 294072 80390 294128
rect 95790 294208 95846 294264
rect 99654 295432 99710 295488
rect 101586 292576 101642 292632
rect 104162 292576 104218 292632
rect 105450 292712 105506 292768
rect 108210 291896 108266 291952
rect 111798 295296 111854 295352
rect 113178 293936 113234 293992
rect 116582 293120 116638 293176
rect 69754 291236 69810 291272
rect 69754 291216 69756 291236
rect 69756 291216 69808 291236
rect 69808 291216 69810 291236
rect 69110 288360 69166 288416
rect 119894 290536 119950 290592
rect 119802 286728 119858 286784
rect 69018 278840 69074 278896
rect 69018 246200 69074 246256
rect 68282 245656 68338 245712
rect 67638 245556 67640 245576
rect 67640 245556 67692 245576
rect 67692 245556 67694 245576
rect 67638 245520 67694 245556
rect 67638 244840 67694 244896
rect 67822 244160 67878 244216
rect 67730 243480 67786 243536
rect 67638 242836 67640 242856
rect 67640 242836 67692 242856
rect 67692 242836 67694 242856
rect 67638 242800 67694 242836
rect 67730 242120 67786 242176
rect 67638 241460 67694 241496
rect 67638 241440 67640 241460
rect 67640 241440 67692 241460
rect 67692 241440 67694 241460
rect 120722 293936 120778 293992
rect 120170 261160 120226 261216
rect 120170 250960 120226 251016
rect 120078 247560 120134 247616
rect 70582 239808 70638 239864
rect 77114 224168 77170 224224
rect 77298 189624 77354 189680
rect 73250 186904 73306 186960
rect 84382 221448 84438 221504
rect 91282 238448 91338 238504
rect 97354 179424 97410 179480
rect 97354 176840 97410 176896
rect 103610 204856 103666 204912
rect 110418 214512 110474 214568
rect 100666 177520 100722 177576
rect 106186 177520 106242 177576
rect 107566 177520 107622 177576
rect 118330 238584 118386 238640
rect 121642 291760 121698 291816
rect 121734 291080 121790 291136
rect 121642 290400 121698 290456
rect 121642 289756 121644 289776
rect 121644 289756 121696 289776
rect 121696 289756 121698 289776
rect 121642 289720 121698 289756
rect 121642 289040 121698 289096
rect 121826 288360 121882 288416
rect 121642 287020 121698 287056
rect 121642 287000 121644 287020
rect 121644 287000 121696 287020
rect 121696 287000 121698 287020
rect 122194 287680 122250 287736
rect 121550 285676 121552 285696
rect 121552 285676 121604 285696
rect 121604 285676 121606 285696
rect 121550 285640 121606 285676
rect 121550 284960 121606 285016
rect 121642 284280 121698 284336
rect 121550 283600 121606 283656
rect 121550 282940 121606 282976
rect 121550 282920 121552 282940
rect 121552 282920 121604 282940
rect 121604 282920 121606 282940
rect 121550 282240 121606 282296
rect 121642 280880 121698 280936
rect 121550 280236 121552 280256
rect 121552 280236 121604 280256
rect 121604 280236 121606 280256
rect 121550 280200 121606 280236
rect 121642 279520 121698 279576
rect 121550 278860 121606 278896
rect 121550 278840 121552 278860
rect 121552 278840 121604 278860
rect 121604 278840 121606 278860
rect 121642 278160 121698 278216
rect 121550 277480 121606 277536
rect 122102 281560 122158 281616
rect 121642 276800 121698 276856
rect 121550 276120 121606 276176
rect 121734 275440 121790 275496
rect 121550 274760 121606 274816
rect 121642 274080 121698 274136
rect 121550 273400 121606 273456
rect 121642 272720 121698 272776
rect 121550 271360 121606 271416
rect 121642 270000 121698 270056
rect 121550 269320 121606 269376
rect 121826 268640 121882 268696
rect 121550 267960 121606 268016
rect 121458 267280 121514 267336
rect 121550 265920 121606 265976
rect 121458 265240 121514 265296
rect 121458 264560 121514 264616
rect 121458 263880 121514 263936
rect 122194 266600 122250 266656
rect 121642 263200 121698 263256
rect 121458 262520 121514 262576
rect 121458 261840 121514 261896
rect 121458 259800 121514 259856
rect 122102 259120 122158 259176
rect 121458 258440 121514 258496
rect 121642 257760 121698 257816
rect 121458 257116 121460 257136
rect 121460 257116 121512 257136
rect 121512 257116 121514 257136
rect 121458 257080 121514 257116
rect 121458 256436 121460 256456
rect 121460 256436 121512 256456
rect 121512 256436 121514 256456
rect 121458 256400 121514 256436
rect 121550 255720 121606 255776
rect 121550 255040 121606 255096
rect 121458 254360 121514 254416
rect 121550 253680 121606 253736
rect 121458 253000 121514 253056
rect 121642 252320 121698 252376
rect 121458 251640 121514 251696
rect 125046 292712 125102 292768
rect 121550 250280 121606 250336
rect 121458 249600 121514 249656
rect 121458 248920 121514 248976
rect 121458 248240 121514 248296
rect 121550 246880 121606 246936
rect 120722 246336 120778 246392
rect 121642 246200 121698 246256
rect 121550 245520 121606 245576
rect 121458 244840 121514 244896
rect 121550 244160 121606 244216
rect 121458 243480 121514 243536
rect 121642 243480 121698 243536
rect 121458 242836 121460 242856
rect 121460 242836 121512 242856
rect 121512 242836 121514 242856
rect 121458 242800 121514 242836
rect 121550 242120 121606 242176
rect 121458 241440 121514 241496
rect 122102 240760 122158 240816
rect 121550 240080 121606 240136
rect 126978 293120 127034 293176
rect 152462 196560 152518 196616
rect 166262 236544 166318 236600
rect 110694 177520 110750 177576
rect 112166 177520 112222 177576
rect 114374 177520 114430 177576
rect 117226 177520 117282 177576
rect 118606 177520 118662 177576
rect 124126 177520 124182 177576
rect 125046 177520 125102 177576
rect 126794 177520 126850 177576
rect 121182 177112 121238 177168
rect 133142 177112 133198 177168
rect 99102 176704 99158 176760
rect 102046 176704 102102 176760
rect 108118 176704 108174 176760
rect 110050 176704 110106 176760
rect 115846 176704 115902 176760
rect 127070 176724 127126 176760
rect 127070 176704 127072 176724
rect 127072 176704 127124 176724
rect 127124 176704 127126 176724
rect 128174 176704 128230 176760
rect 129462 176704 129518 176760
rect 132038 176704 132094 176760
rect 134706 176704 134762 176760
rect 135718 176740 135720 176760
rect 135720 176740 135772 176760
rect 135772 176740 135774 176760
rect 135718 176704 135774 176740
rect 148230 176704 148286 176760
rect 100758 175344 100814 175400
rect 130750 175480 130806 175536
rect 158902 175480 158958 175536
rect 121918 175344 121974 175400
rect 119434 174936 119490 174992
rect 67362 129240 67418 129296
rect 64970 126248 65026 126304
rect 64970 125568 65026 125624
rect 66166 125160 66222 125216
rect 66074 123528 66130 123584
rect 66074 102312 66130 102368
rect 67270 100680 67326 100736
rect 66166 91024 66222 91080
rect 67638 128016 67694 128072
rect 67454 122576 67510 122632
rect 67546 120808 67602 120864
rect 167642 171536 167698 171592
rect 105450 94696 105506 94752
rect 117962 94696 118018 94752
rect 119526 94696 119582 94752
rect 129370 94696 129426 94752
rect 134338 94696 134394 94752
rect 67638 93744 67694 93800
rect 130750 93608 130806 93664
rect 151726 93608 151782 93664
rect 110694 93472 110750 93528
rect 115846 93472 115902 93528
rect 110326 93200 110382 93256
rect 85670 92384 85726 92440
rect 91650 92384 91706 92440
rect 107750 92384 107806 92440
rect 89350 91704 89406 91760
rect 90546 91704 90602 91760
rect 75366 91160 75422 91216
rect 85486 91160 85542 91216
rect 86866 91160 86922 91216
rect 88062 91160 88118 91216
rect 99746 91704 99802 91760
rect 99286 91432 99342 91488
rect 95054 91296 95110 91352
rect 97814 91296 97870 91352
rect 99102 91296 99158 91352
rect 93766 91160 93822 91216
rect 95146 91160 95202 91216
rect 96526 91160 96582 91216
rect 96526 84088 96582 84144
rect 97906 91160 97962 91216
rect 99194 91160 99250 91216
rect 103150 91568 103206 91624
rect 102046 91432 102102 91488
rect 101862 91296 101918 91352
rect 100574 91160 100630 91216
rect 101954 91160 102010 91216
rect 101954 82728 102010 82784
rect 107566 91296 107622 91352
rect 103426 91160 103482 91216
rect 104346 91160 104402 91216
rect 104622 91160 104678 91216
rect 107474 91160 107530 91216
rect 104622 88168 104678 88224
rect 109222 91160 109278 91216
rect 109774 91160 109830 91216
rect 128174 93200 128230 93256
rect 114190 92384 114246 92440
rect 115478 92420 115480 92440
rect 115480 92420 115532 92440
rect 115532 92420 115534 92440
rect 115478 92384 115534 92420
rect 116766 92404 116822 92440
rect 116766 92384 116768 92404
rect 116768 92384 116820 92404
rect 116820 92384 116822 92404
rect 111614 91160 111670 91216
rect 111982 91160 112038 91216
rect 112350 91160 112406 91216
rect 119710 92384 119766 92440
rect 122470 92384 122526 92440
rect 117134 91704 117190 91760
rect 114466 91160 114522 91216
rect 115294 91160 115350 91216
rect 107566 80008 107622 80064
rect 121274 91296 121330 91352
rect 118606 91160 118662 91216
rect 121366 91160 121422 91216
rect 121274 83952 121330 84008
rect 125782 92384 125838 92440
rect 125506 92112 125562 92168
rect 122838 91432 122894 91488
rect 122746 91160 122802 91216
rect 123574 91160 123630 91216
rect 124126 91160 124182 91216
rect 125414 91160 125470 91216
rect 123574 86808 123630 86864
rect 126518 91160 126574 91216
rect 126886 91160 126942 91216
rect 151542 92384 151598 92440
rect 152094 92384 152150 92440
rect 151450 92112 151506 92168
rect 136454 91432 136510 91488
rect 132038 91160 132094 91216
rect 133142 91160 133198 91216
rect 128174 89664 128230 89720
rect 167918 111732 167920 111752
rect 167920 111732 167972 111752
rect 167972 111732 167974 111752
rect 167918 111696 167974 111732
rect 168194 110064 168250 110120
rect 167734 108704 167790 108760
rect 174542 89664 174598 89720
rect 112442 43424 112498 43480
rect 180062 294208 180118 294264
rect 178682 184320 178738 184376
rect 180062 95104 180118 95160
rect 180154 92248 180210 92304
rect 189722 179968 189778 180024
rect 210422 175888 210478 175944
rect 214562 188264 214618 188320
rect 213918 175616 213974 175672
rect 213918 174936 213974 174992
rect 214010 174256 214066 174312
rect 213918 173576 213974 173632
rect 214102 172896 214158 172952
rect 213918 172216 213974 172272
rect 214010 171536 214066 171592
rect 214010 171012 214066 171048
rect 214010 170992 214012 171012
rect 214012 170992 214064 171012
rect 214064 170992 214066 171012
rect 213918 170312 213974 170368
rect 214010 169652 214066 169688
rect 214010 169632 214012 169652
rect 214012 169632 214064 169652
rect 214064 169632 214066 169652
rect 213918 168952 213974 169008
rect 213918 168292 213974 168328
rect 213918 168272 213920 168292
rect 213920 168272 213972 168292
rect 213972 168272 213974 168292
rect 214010 167592 214066 167648
rect 213918 166948 213920 166968
rect 213920 166948 213972 166968
rect 213972 166948 213974 166968
rect 213918 166912 213974 166948
rect 214010 166368 214066 166424
rect 213918 165008 213974 165064
rect 214010 164328 214066 164384
rect 213918 162968 213974 163024
rect 213918 162288 213974 162344
rect 213918 161064 213974 161120
rect 214010 160384 214066 160440
rect 214470 159704 214526 159760
rect 213918 157664 213974 157720
rect 214010 157120 214066 157176
rect 213918 156440 213974 156496
rect 213918 155760 213974 155816
rect 213918 154400 213974 154456
rect 214010 153040 214066 153096
rect 213918 152496 213974 152552
rect 213274 151816 213330 151872
rect 209134 94832 209190 94888
rect 214010 151136 214066 151192
rect 213918 149776 213974 149832
rect 214010 149096 214066 149152
rect 224314 180104 224370 180160
rect 214654 165688 214710 165744
rect 240782 176024 240838 176080
rect 248418 177520 248474 177576
rect 248050 175752 248106 175808
rect 249246 175208 249302 175264
rect 249154 174664 249210 174720
rect 249154 172760 249210 172816
rect 249798 171808 249854 171864
rect 214746 161744 214802 161800
rect 249798 155352 249854 155408
rect 215942 153720 215998 153776
rect 214654 150456 214710 150512
rect 214562 148416 214618 148472
rect 213918 147872 213974 147928
rect 214010 147192 214066 147248
rect 213918 146512 213974 146568
rect 214010 145832 214066 145888
rect 213918 145152 213974 145208
rect 214010 144472 214066 144528
rect 213918 143792 213974 143848
rect 214010 143248 214066 143304
rect 213918 142568 213974 142624
rect 213918 141888 213974 141944
rect 213918 140528 213974 140584
rect 213918 138624 213974 138680
rect 214102 137944 214158 138000
rect 213918 137264 213974 137320
rect 214010 136584 214066 136640
rect 213918 135260 213920 135280
rect 213920 135260 213972 135280
rect 213972 135260 213974 135280
rect 213918 135224 213974 135260
rect 214010 134544 214066 134600
rect 213918 133864 213974 133920
rect 213918 133320 213974 133376
rect 214654 139168 214710 139224
rect 213918 131960 213974 132016
rect 213918 130600 213974 130656
rect 214010 129240 214066 129296
rect 213918 128696 213974 128752
rect 214010 128016 214066 128072
rect 213918 127336 213974 127392
rect 214010 126656 214066 126712
rect 213918 125976 213974 126032
rect 214010 125296 214066 125352
rect 213918 124616 213974 124672
rect 214010 124072 214066 124128
rect 213918 123392 213974 123448
rect 214010 122712 214066 122768
rect 213918 122032 213974 122088
rect 214010 121352 214066 121408
rect 213918 120672 213974 120728
rect 214010 119992 214066 120048
rect 213918 118768 213974 118824
rect 214102 119448 214158 119504
rect 213918 118088 213974 118144
rect 213182 117408 213238 117464
rect 211894 91568 211950 91624
rect 214010 116728 214066 116784
rect 213918 116068 213974 116104
rect 213918 116048 213920 116068
rect 213920 116048 213972 116068
rect 213972 116048 213974 116068
rect 214010 115368 214066 115424
rect 213918 114824 213974 114880
rect 214010 114144 214066 114200
rect 213918 113464 213974 113520
rect 214010 112784 214066 112840
rect 213918 112104 213974 112160
rect 214010 111424 214066 111480
rect 213918 110744 213974 110800
rect 213918 110200 213974 110256
rect 214010 108840 214066 108896
rect 213918 108160 213974 108216
rect 213918 107480 213974 107536
rect 214010 106120 214066 106176
rect 213918 105576 213974 105632
rect 213918 104216 213974 104272
rect 213918 102196 213974 102232
rect 213918 102176 213920 102196
rect 213920 102176 213972 102196
rect 213972 102176 213974 102196
rect 214010 101496 214066 101552
rect 213918 100952 213974 101008
rect 214010 100272 214066 100328
rect 213918 99592 213974 99648
rect 213918 98912 213974 98968
rect 213918 97552 213974 97608
rect 214654 106800 214710 106856
rect 214562 96328 214618 96384
rect 214838 98232 214894 98288
rect 214746 96872 214802 96928
rect 250166 166640 250222 166696
rect 251178 159568 251234 159624
rect 251362 164328 251418 164384
rect 251362 162968 251418 163024
rect 251822 173304 251878 173360
rect 252466 172388 252468 172408
rect 252468 172388 252520 172408
rect 252520 172388 252522 172408
rect 252466 172352 252522 172388
rect 252006 171400 252062 171456
rect 251822 170448 251878 170504
rect 252466 170892 252468 170912
rect 252468 170892 252520 170912
rect 252520 170892 252522 170912
rect 252466 170856 252522 170892
rect 252098 170040 252154 170096
rect 252466 169088 252522 169144
rect 252006 168544 252062 168600
rect 251914 168172 251916 168192
rect 251916 168172 251968 168192
rect 251968 168172 251970 168192
rect 251914 168136 251970 168172
rect 252466 167592 252522 167648
rect 252098 167184 252154 167240
rect 251822 166232 251878 166288
rect 252466 165280 252522 165336
rect 252374 164736 252430 164792
rect 252466 163920 252522 163976
rect 252466 162424 252522 162480
rect 252098 161472 252154 161528
rect 251270 158752 251326 158808
rect 250442 152904 250498 152960
rect 249982 150728 250038 150784
rect 249890 138896 249946 138952
rect 249890 138080 249946 138136
rect 251178 152088 251234 152144
rect 251270 151136 251326 151192
rect 251270 148860 251272 148880
rect 251272 148860 251324 148880
rect 251324 148860 251326 148880
rect 251270 148824 251326 148860
rect 252098 161064 252154 161120
rect 252466 160520 252522 160576
rect 252006 160112 252062 160168
rect 252466 159160 252522 159216
rect 252466 158208 252522 158264
rect 252374 157800 252430 157856
rect 252466 157276 252522 157312
rect 252466 157256 252468 157276
rect 252468 157256 252520 157276
rect 252520 157256 252522 157276
rect 252374 156848 252430 156904
rect 252466 155896 252522 155952
rect 252374 154944 252430 155000
rect 252650 169496 252706 169552
rect 252742 165688 252798 165744
rect 252558 154400 252614 154456
rect 252466 153992 252522 154048
rect 252374 153448 252430 153504
rect 252466 153040 252522 153096
rect 252466 151716 252468 151736
rect 252468 151716 252520 151736
rect 252520 151716 252522 151736
rect 252466 151680 252522 151716
rect 252282 149776 252338 149832
rect 251730 149268 251732 149288
rect 251732 149268 251784 149288
rect 251784 149268 251786 149288
rect 251730 149232 251786 149268
rect 251914 148280 251970 148336
rect 252466 147872 252522 147928
rect 252466 147464 252522 147520
rect 251730 146920 251786 146976
rect 251730 146512 251786 146568
rect 251914 145968 251970 146024
rect 251730 145560 251786 145616
rect 252098 145016 252154 145072
rect 251270 140800 251326 140856
rect 251362 139884 251364 139904
rect 251364 139884 251416 139904
rect 251416 139884 251418 139904
rect 251362 139848 251418 139884
rect 251362 137944 251418 138000
rect 250442 136584 250498 136640
rect 251546 136176 251602 136232
rect 251638 134680 251694 134736
rect 251454 133320 251510 133376
rect 251362 132368 251418 132424
rect 251730 130464 251786 130520
rect 251730 129104 251786 129160
rect 251546 127608 251602 127664
rect 251270 124344 251326 124400
rect 251362 119584 251418 119640
rect 252006 131416 252062 131472
rect 252006 130056 252062 130112
rect 252466 144608 252522 144664
rect 252374 144064 252430 144120
rect 252466 143656 252522 143712
rect 252466 143112 252522 143168
rect 252466 141344 252522 141400
rect 252466 138488 252522 138544
rect 252466 136992 252522 137048
rect 252466 135632 252522 135688
rect 252374 135224 252430 135280
rect 252466 134272 252522 134328
rect 252466 132776 252522 132832
rect 252282 131824 252338 131880
rect 252466 130872 252522 130928
rect 252006 129512 252062 129568
rect 252098 128560 252154 128616
rect 252466 128188 252468 128208
rect 252468 128188 252520 128208
rect 252520 128188 252522 128208
rect 252466 128152 252522 128188
rect 252006 127200 252062 127256
rect 251914 126248 251970 126304
rect 252466 126656 252522 126712
rect 252098 125704 252154 125760
rect 252466 125296 252522 125352
rect 252374 124752 252430 124808
rect 252282 123936 252338 123992
rect 252006 122984 252062 123040
rect 252466 123392 252522 123448
rect 251914 120128 251970 120184
rect 251822 119176 251878 119232
rect 251178 117272 251234 117328
rect 251822 117816 251878 117872
rect 251914 116320 251970 116376
rect 251638 114416 251694 114472
rect 252466 122440 252522 122496
rect 252374 122032 252430 122088
rect 252466 121488 252522 121544
rect 252466 121080 252522 121136
rect 252374 120536 252430 120592
rect 252466 118768 252522 118824
rect 253386 142704 253442 142760
rect 253386 142296 253442 142352
rect 252466 118224 252522 118280
rect 252466 116864 252522 116920
rect 252374 115912 252430 115968
rect 252466 115368 252522 115424
rect 252374 114960 252430 115016
rect 252466 114008 252522 114064
rect 252374 113464 252430 113520
rect 252098 113056 252154 113112
rect 252006 112648 252062 112704
rect 252282 111716 252338 111752
rect 252282 111696 252284 111716
rect 252284 111696 252336 111716
rect 252336 111696 252338 111716
rect 251546 110744 251602 110800
rect 252466 112104 252522 112160
rect 252466 111152 252522 111208
rect 252466 110200 252522 110256
rect 252374 109792 252430 109848
rect 251914 109284 251916 109304
rect 251916 109284 251968 109304
rect 251968 109284 251970 109304
rect 251914 109248 251970 109284
rect 252466 108876 252468 108896
rect 252468 108876 252520 108896
rect 252520 108876 252522 108896
rect 252466 108840 252522 108876
rect 251730 108296 251786 108352
rect 251362 107888 251418 107944
rect 251270 107480 251326 107536
rect 252466 106936 252522 106992
rect 251362 106528 251418 106584
rect 252006 105984 252062 106040
rect 252282 105576 252338 105632
rect 252006 104624 252062 104680
rect 251178 103672 251234 103728
rect 216034 102856 216090 102912
rect 251178 102756 251180 102776
rect 251180 102756 251232 102776
rect 251232 102756 251234 102776
rect 251178 102720 251234 102756
rect 252466 104080 252522 104136
rect 252466 103128 252522 103184
rect 251546 102176 251602 102232
rect 252466 101768 252522 101824
rect 252374 101360 252430 101416
rect 252098 100816 252154 100872
rect 251178 99864 251234 99920
rect 252466 100408 252522 100464
rect 252098 99456 252154 99512
rect 251178 98504 251234 98560
rect 252282 98912 252338 98968
rect 252190 97960 252246 98016
rect 252466 97552 252522 97608
rect 251178 97008 251234 97064
rect 249154 96600 249210 96656
rect 249522 96600 249578 96656
rect 248418 95648 248474 95704
rect 125874 3304 125930 3360
rect 255962 144064 256018 144120
rect 256974 175888 257030 175944
rect 269946 133048 270002 133104
rect 274086 138624 274142 138680
rect 300122 181328 300178 181384
rect 305642 178744 305698 178800
rect 307114 178608 307170 178664
rect 307022 175208 307078 175264
rect 306746 174800 306802 174856
rect 282182 155216 282238 155272
rect 306930 173168 306986 173224
rect 306930 170992 306986 171048
rect 306562 165008 306618 165064
rect 293498 142704 293554 142760
rect 292118 141344 292174 141400
rect 306562 160792 306618 160848
rect 306930 159976 306986 160032
rect 306930 158616 306986 158672
rect 306746 156984 306802 157040
rect 306654 153176 306710 153232
rect 305826 146376 305882 146432
rect 305734 118904 305790 118960
rect 305642 105440 305698 105496
rect 306930 150592 306986 150648
rect 306930 150184 306986 150240
rect 307666 174392 307722 174448
rect 307574 173984 307630 174040
rect 307666 173576 307722 173632
rect 307298 172660 307300 172680
rect 307300 172660 307352 172680
rect 307352 172660 307354 172680
rect 307298 172624 307354 172660
rect 307482 172216 307538 172272
rect 307574 171808 307630 171864
rect 307666 171400 307722 171456
rect 307482 170584 307538 170640
rect 307666 170176 307722 170232
rect 307206 169768 307262 169824
rect 307482 169224 307538 169280
rect 307666 168816 307722 168872
rect 307298 168408 307354 168464
rect 307482 168000 307538 168056
rect 307574 167592 307630 167648
rect 307666 167204 307722 167240
rect 307666 167184 307668 167204
rect 307668 167184 307720 167204
rect 307720 167184 307722 167204
rect 307666 166776 307722 166832
rect 307482 166368 307538 166424
rect 307298 165824 307354 165880
rect 307482 165416 307538 165472
rect 307666 164600 307722 164656
rect 307574 164192 307630 164248
rect 307482 163784 307538 163840
rect 307666 163376 307722 163432
rect 307298 162968 307354 163024
rect 307482 162424 307538 162480
rect 307298 162016 307354 162072
rect 307666 161608 307722 161664
rect 307666 161200 307722 161256
rect 307114 160384 307170 160440
rect 306930 148824 306986 148880
rect 307022 148416 307078 148472
rect 306746 147192 306802 147248
rect 306562 144608 306618 144664
rect 306746 142976 306802 143032
rect 306930 137808 306986 137864
rect 306746 134816 306802 134872
rect 306746 131416 306802 131472
rect 306746 131008 306802 131064
rect 306930 130192 306986 130248
rect 306746 125840 306802 125896
rect 306746 125432 306802 125488
rect 306562 123800 306618 123856
rect 306746 119992 306802 120048
rect 306746 116592 306802 116648
rect 306746 115640 306802 115696
rect 306746 114416 306802 114472
rect 307482 159568 307538 159624
rect 307666 159024 307722 159080
rect 307482 158208 307538 158264
rect 307298 157800 307354 157856
rect 307390 157392 307446 157448
rect 307206 154400 307262 154456
rect 307574 156576 307630 156632
rect 307666 156168 307722 156224
rect 307482 155624 307538 155680
rect 307574 155216 307630 155272
rect 307666 154808 307722 154864
rect 307482 153992 307538 154048
rect 307666 153584 307722 153640
rect 307482 152632 307538 152688
rect 307666 152224 307722 152280
rect 307666 151836 307722 151872
rect 307666 151816 307668 151836
rect 307668 151816 307720 151836
rect 307720 151816 307722 151836
rect 307482 151408 307538 151464
rect 307666 151000 307722 151056
rect 307666 149776 307722 149832
rect 307574 149232 307630 149288
rect 307666 148008 307722 148064
rect 307390 147600 307446 147656
rect 307666 146784 307722 146840
rect 307482 145832 307538 145888
rect 307298 142024 307354 142080
rect 307206 140392 307262 140448
rect 307114 136992 307170 137048
rect 306746 108840 306802 108896
rect 306010 108432 306066 108488
rect 305826 104216 305882 104272
rect 306562 105848 306618 105904
rect 306746 103400 306802 103456
rect 306930 102448 306986 102504
rect 306746 97824 306802 97880
rect 307022 97008 307078 97064
rect 307390 141616 307446 141672
rect 307574 145424 307630 145480
rect 307666 145036 307722 145072
rect 307666 145016 307668 145036
rect 307668 145016 307720 145036
rect 307720 145016 307722 145036
rect 307666 144200 307722 144256
rect 307666 143384 307722 143440
rect 307666 141208 307722 141264
rect 307574 139984 307630 140040
rect 307666 139576 307722 139632
rect 307482 139032 307538 139088
rect 307574 138624 307630 138680
rect 307666 138216 307722 138272
rect 307482 137400 307538 137456
rect 307390 136584 307446 136640
rect 307666 136176 307722 136232
rect 307482 135632 307538 135688
rect 307574 135224 307630 135280
rect 307574 134408 307630 134464
rect 307666 134036 307668 134056
rect 307668 134036 307720 134056
rect 307720 134036 307722 134056
rect 307666 134000 307722 134036
rect 307666 133592 307722 133648
rect 307482 133184 307538 133240
rect 307482 132232 307538 132288
rect 307666 131824 307722 131880
rect 307666 129804 307722 129840
rect 307666 129784 307668 129804
rect 307668 129784 307720 129804
rect 307720 129784 307722 129804
rect 307482 129240 307538 129296
rect 307574 128832 307630 128888
rect 307666 128460 307668 128480
rect 307668 128460 307720 128480
rect 307720 128460 307722 128480
rect 307666 128424 307722 128460
rect 307482 128016 307538 128072
rect 307574 127608 307630 127664
rect 307666 127200 307722 127256
rect 307482 126792 307538 126848
rect 307666 126384 307722 126440
rect 307482 125024 307538 125080
rect 307298 124616 307354 124672
rect 307206 116184 307262 116240
rect 307666 124228 307722 124264
rect 307666 124208 307668 124228
rect 307668 124208 307720 124228
rect 307720 124208 307722 124228
rect 307574 123392 307630 123448
rect 307666 123004 307722 123040
rect 307666 122984 307668 123004
rect 307668 122984 307720 123004
rect 307720 122984 307722 123004
rect 307482 122440 307538 122496
rect 307574 122032 307630 122088
rect 307666 121644 307722 121680
rect 307666 121624 307668 121644
rect 307668 121624 307720 121644
rect 307720 121624 307722 121644
rect 307482 121216 307538 121272
rect 307574 120808 307630 120864
rect 307666 120400 307722 120456
rect 307574 119584 307630 119640
rect 307666 119040 307722 119096
rect 307574 118904 307630 118960
rect 307482 118632 307538 118688
rect 307574 117816 307630 117872
rect 307666 117428 307722 117464
rect 307666 117408 307668 117428
rect 307668 117408 307720 117428
rect 307720 117408 307722 117428
rect 307666 117000 307722 117056
rect 307666 114824 307722 114880
rect 307574 113600 307630 113656
rect 307666 113212 307722 113248
rect 307666 113192 307668 113212
rect 307668 113192 307720 113212
rect 307720 113192 307722 113212
rect 307574 112240 307630 112296
rect 307666 111852 307722 111888
rect 307666 111832 307668 111852
rect 307668 111832 307720 111852
rect 307720 111832 307722 111852
rect 307482 111424 307538 111480
rect 307574 111016 307630 111072
rect 307666 110608 307722 110664
rect 307482 110200 307538 110256
rect 307574 109792 307630 109848
rect 307666 109248 307722 109304
rect 307574 108024 307630 108080
rect 307666 107616 307722 107672
rect 307482 107208 307538 107264
rect 307574 106800 307630 106856
rect 307666 106392 307722 106448
rect 307666 105052 307722 105088
rect 307666 105032 307668 105052
rect 307668 105032 307720 105052
rect 307720 105032 307722 105052
rect 307574 104624 307630 104680
rect 307666 103808 307722 103864
rect 307482 102992 307538 103048
rect 307574 102040 307630 102096
rect 307482 101632 307538 101688
rect 307666 100836 307722 100872
rect 307666 100816 307668 100836
rect 307668 100816 307720 100836
rect 307720 100816 307722 100836
rect 307482 100408 307538 100464
rect 307666 100000 307722 100056
rect 307482 99048 307538 99104
rect 307666 98640 307722 98696
rect 307574 98232 307630 98288
rect 307482 97416 307538 97472
rect 307666 96192 307722 96248
rect 308494 95920 308550 95976
rect 313922 177248 313978 177304
rect 316038 176704 316094 176760
rect 312542 175888 312598 175944
rect 325698 290536 325754 290592
rect 320178 176704 320234 176760
rect 319442 176568 319498 176624
rect 321466 176024 321522 176080
rect 321466 175208 321522 175264
rect 321374 173712 321430 173768
rect 321282 165008 321338 165064
rect 321834 172624 321890 172680
rect 321650 165688 321706 165744
rect 322938 153176 322994 153232
rect 321742 151272 321798 151328
rect 324318 169360 324374 169416
rect 324410 168544 324466 168600
rect 324318 167728 324374 167784
rect 324410 167048 324466 167104
rect 324318 166232 324374 166288
rect 324318 163920 324374 163976
rect 324410 163104 324466 163160
rect 324318 162424 324374 162480
rect 324410 161608 324466 161664
rect 324318 160112 324374 160168
rect 324318 159296 324374 159352
rect 324318 158480 324374 158536
rect 324410 157800 324466 157856
rect 324318 156984 324374 157040
rect 324410 156304 324466 156360
rect 324318 155488 324374 155544
rect 324502 154672 324558 154728
rect 324318 153992 324374 154048
rect 324318 152360 324374 152416
rect 324318 151716 324320 151736
rect 324320 151716 324372 151736
rect 324372 151716 324374 151736
rect 324318 151680 324374 151716
rect 324318 150048 324374 150104
rect 324410 149368 324466 149424
rect 324318 148552 324374 148608
rect 324410 147736 324466 147792
rect 324318 147056 324374 147112
rect 324318 146240 324374 146296
rect 324410 145424 324466 145480
rect 324318 144744 324374 144800
rect 324410 143928 324466 143984
rect 324318 142432 324374 142488
rect 324318 141616 324374 141672
rect 324318 139340 324320 139360
rect 324320 139340 324372 139360
rect 324372 139340 324374 139360
rect 324318 139304 324374 139340
rect 324318 137808 324374 137864
rect 324318 136312 324374 136368
rect 324318 133184 324374 133240
rect 324318 132388 324374 132424
rect 324318 132368 324320 132388
rect 324320 132368 324372 132388
rect 324372 132368 324374 132388
rect 324502 140800 324558 140856
rect 324502 138488 324558 138544
rect 324502 136992 324558 137048
rect 324502 135496 324558 135552
rect 324502 131688 324558 131744
rect 324318 130872 324374 130928
rect 324410 130056 324466 130112
rect 324318 128560 324374 128616
rect 324318 127744 324374 127800
rect 324318 126248 324374 126304
rect 324502 125432 324558 125488
rect 324318 123936 324374 123992
rect 324318 121624 324374 121680
rect 324318 120808 324374 120864
rect 324410 120128 324466 120184
rect 324502 119312 324558 119368
rect 324318 118532 324320 118552
rect 324320 118532 324372 118552
rect 324372 118532 324374 118552
rect 324318 118496 324374 118532
rect 324410 117816 324466 117872
rect 324318 117000 324374 117056
rect 324410 116320 324466 116376
rect 324318 115504 324374 115560
rect 324318 114008 324374 114064
rect 324410 113192 324466 113248
rect 324318 112376 324374 112432
rect 324318 111732 324320 111752
rect 324320 111732 324372 111752
rect 324372 111732 324374 111752
rect 324318 111696 324374 111732
rect 324410 108568 324466 108624
rect 324318 107752 324374 107808
rect 323490 106528 323546 106584
rect 323490 106256 323546 106312
rect 321558 105984 321614 106040
rect 324318 103128 324374 103184
rect 321742 98096 321798 98152
rect 321558 97280 321614 97336
rect 321466 96620 321522 96656
rect 321466 96600 321468 96620
rect 321468 96600 321520 96620
rect 321520 96600 321522 96620
rect 321650 96600 321706 96656
rect 321650 95104 321706 95160
rect 324686 160792 324742 160848
rect 324686 142704 324742 142760
rect 324686 140120 324742 140176
rect 325606 124752 325662 124808
rect 325882 176568 325938 176624
rect 325882 171672 325938 171728
rect 325790 134000 325846 134056
rect 324962 123120 325018 123176
rect 324686 122440 324742 122496
rect 346398 292576 346454 292632
rect 345110 291252 345112 291272
rect 345112 291252 345164 291272
rect 345164 291252 345166 291272
rect 345110 291216 345166 291252
rect 345294 182824 345350 182880
rect 324594 100816 324650 100872
rect 580906 697176 580962 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 582378 590960 582434 591016
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580262 511264 580318 511320
rect 580170 484608 580226 484664
rect 580170 471416 580226 471472
rect 580170 458088 580226 458144
rect 579894 431568 579950 431624
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 579618 365064 579674 365120
rect 580170 351908 580172 351928
rect 580172 351908 580224 351928
rect 580224 351908 580226 351928
rect 580170 351872 580226 351908
rect 580170 325216 580226 325272
rect 580170 312024 580226 312080
rect 579618 258848 579674 258904
rect 579894 245520 579950 245576
rect 580170 205672 580226 205728
rect 579986 179152 580042 179208
rect 580354 279656 580410 279712
rect 580446 272176 580502 272232
rect 580446 264152 580502 264208
rect 582470 537784 582526 537840
rect 582746 298696 582802 298752
rect 580446 232328 580502 232384
rect 580354 219000 580410 219056
rect 580262 152632 580318 152688
rect 580170 125976 580226 126032
rect 324502 100136 324558 100192
rect 580170 99456 580226 99512
rect 580170 59608 580226 59664
rect 582470 46280 582526 46336
rect 582838 231104 582894 231160
rect 582654 112784 582710 112840
rect 582838 86128 582894 86184
rect 582746 33088 582802 33144
rect 582562 19760 582618 19816
rect 582378 6568 582434 6624
<< obsm2 >>
rect 68800 95100 164756 174600
<< metal3 >>
rect -960 697220 480 697460
rect 580901 697234 580967 697237
rect 583520 697234 584960 697324
rect 580901 697232 584960 697234
rect 580901 697176 580906 697232
rect 580962 697176 584960 697232
rect 580901 697174 584960 697176
rect 580901 697171 580967 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3509 658202 3575 658205
rect -960 658200 3575 658202
rect -960 658144 3514 658200
rect 3570 658144 3575 658200
rect -960 658142 3575 658144
rect -960 658052 480 658142
rect 3509 658139 3575 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 644058 584960 644148
rect 583342 643998 584960 644058
rect 583342 643922 583402 643998
rect 583520 643922 584960 643998
rect 583342 643908 584960 643922
rect 583342 643862 583586 643908
rect 120574 643180 120580 643244
rect 120644 643242 120650 643244
rect 583526 643242 583586 643862
rect 120644 643182 583586 643242
rect 120644 643180 120650 643182
rect -960 632090 480 632180
rect 3509 632090 3575 632093
rect -960 632088 3575 632090
rect -960 632032 3514 632088
rect 3570 632032 3575 632088
rect -960 632030 3575 632032
rect -960 631940 480 632030
rect 3509 632027 3575 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 2773 606114 2839 606117
rect -960 606112 2839 606114
rect -960 606056 2778 606112
rect 2834 606056 2839 606112
rect -960 606054 2839 606056
rect -960 605964 480 606054
rect 2773 606051 2839 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 582373 591018 582439 591021
rect 583520 591018 584960 591108
rect 582373 591016 584960 591018
rect 582373 590960 582378 591016
rect 582434 590960 584960 591016
rect 582373 590958 584960 590960
rect 582373 590955 582439 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3233 566946 3299 566949
rect -960 566944 3299 566946
rect -960 566888 3238 566944
rect 3294 566888 3299 566944
rect -960 566886 3299 566888
rect -960 566796 480 566886
rect 3233 566883 3299 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 582465 537842 582531 537845
rect 583520 537842 584960 537932
rect 582465 537840 584960 537842
rect 582465 537784 582470 537840
rect 582526 537784 584960 537840
rect 582465 537782 584960 537784
rect 582465 537779 582531 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 2957 527914 3023 527917
rect -960 527912 3023 527914
rect -960 527856 2962 527912
rect 3018 527856 3023 527912
rect -960 527854 3023 527856
rect -960 527764 480 527854
rect 2957 527851 3023 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3509 514858 3575 514861
rect -960 514856 3575 514858
rect -960 514800 3514 514856
rect 3570 514800 3575 514856
rect -960 514798 3575 514800
rect -960 514708 480 514798
rect 3509 514795 3575 514798
rect 580257 511322 580323 511325
rect 583520 511322 584960 511412
rect 580257 511320 584960 511322
rect 580257 511264 580262 511320
rect 580318 511264 584960 511320
rect 580257 511262 584960 511264
rect 580257 511259 580323 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3325 501802 3391 501805
rect -960 501800 3391 501802
rect -960 501744 3330 501800
rect 3386 501744 3391 501800
rect -960 501742 3391 501744
rect -960 501652 480 501742
rect 3325 501739 3391 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3049 475690 3115 475693
rect -960 475688 3115 475690
rect -960 475632 3054 475688
rect 3110 475632 3115 475688
rect -960 475630 3115 475632
rect -960 475540 480 475630
rect 3049 475627 3115 475630
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3325 462634 3391 462637
rect -960 462632 3391 462634
rect -960 462576 3330 462632
rect 3386 462576 3391 462632
rect -960 462574 3391 462576
rect -960 462484 480 462574
rect 3325 462571 3391 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3325 449578 3391 449581
rect -960 449576 3391 449578
rect -960 449520 3330 449576
rect 3386 449520 3391 449576
rect -960 449518 3391 449520
rect -960 449428 480 449518
rect 3325 449515 3391 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 579889 431626 579955 431629
rect 583520 431626 584960 431716
rect 579889 431624 584960 431626
rect 579889 431568 579894 431624
rect 579950 431568 584960 431624
rect 579889 431566 584960 431568
rect 579889 431563 579955 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3325 423602 3391 423605
rect -960 423600 3391 423602
rect -960 423544 3330 423600
rect 3386 423544 3391 423600
rect -960 423542 3391 423544
rect -960 423452 480 423542
rect 3325 423539 3391 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3325 410546 3391 410549
rect -960 410544 3391 410546
rect -960 410488 3330 410544
rect 3386 410488 3391 410544
rect -960 410486 3391 410488
rect -960 410396 480 410486
rect 3325 410483 3391 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 579613 365122 579679 365125
rect 583520 365122 584960 365212
rect 579613 365120 584960 365122
rect 579613 365064 579618 365120
rect 579674 365064 584960 365120
rect 579613 365062 584960 365064
rect 579613 365059 579679 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3417 306234 3483 306237
rect -960 306232 3483 306234
rect -960 306176 3422 306232
rect 3478 306176 3483 306232
rect -960 306174 3483 306176
rect -960 306084 480 306174
rect 3417 306171 3483 306174
rect 75361 302290 75427 302293
rect 331254 302290 331260 302292
rect 75361 302288 331260 302290
rect 75361 302232 75366 302288
rect 75422 302232 331260 302288
rect 75361 302230 331260 302232
rect 75361 302227 75427 302230
rect 331254 302228 331260 302230
rect 331324 302228 331330 302292
rect 80513 299570 80579 299573
rect 265014 299570 265020 299572
rect 80513 299568 265020 299570
rect 80513 299512 80518 299568
rect 80574 299512 265020 299568
rect 80513 299510 265020 299512
rect 80513 299507 80579 299510
rect 265014 299508 265020 299510
rect 265084 299508 265090 299572
rect 582741 298754 582807 298757
rect 583520 298754 584960 298844
rect 582741 298752 584960 298754
rect 582741 298696 582746 298752
rect 582802 298696 584960 298752
rect 582741 298694 584960 298696
rect 582741 298691 582807 298694
rect 583520 298604 584960 298694
rect 68829 296850 68895 296853
rect 252502 296850 252508 296852
rect 68829 296848 252508 296850
rect 68829 296792 68834 296848
rect 68890 296792 252508 296848
rect 68829 296790 252508 296792
rect 68829 296787 68895 296790
rect 252502 296788 252508 296790
rect 252572 296788 252578 296852
rect 99649 295490 99715 295493
rect 256734 295490 256740 295492
rect 99649 295488 256740 295490
rect 99649 295432 99654 295488
rect 99710 295432 256740 295488
rect 99649 295430 256740 295432
rect 99649 295427 99715 295430
rect 256734 295428 256740 295430
rect 256804 295428 256810 295492
rect 111793 295354 111859 295357
rect 340822 295354 340828 295356
rect 111793 295352 340828 295354
rect 111793 295296 111798 295352
rect 111854 295296 340828 295352
rect 111793 295294 340828 295296
rect 111793 295291 111859 295294
rect 340822 295292 340828 295294
rect 340892 295292 340898 295356
rect 95785 294266 95851 294269
rect 180057 294266 180123 294269
rect 95785 294264 180123 294266
rect 95785 294208 95790 294264
rect 95846 294208 180062 294264
rect 180118 294208 180123 294264
rect 95785 294206 180123 294208
rect 95785 294203 95851 294206
rect 180057 294203 180123 294206
rect 80329 294130 80395 294133
rect 119654 294130 119660 294132
rect 80329 294128 119660 294130
rect 80329 294072 80334 294128
rect 80390 294072 119660 294128
rect 80329 294070 119660 294072
rect 80329 294067 80395 294070
rect 119654 294068 119660 294070
rect 119724 294068 119730 294132
rect 113173 293994 113239 293997
rect 120717 293994 120783 293997
rect 113173 293992 120783 293994
rect 113173 293936 113178 293992
rect 113234 293936 120722 293992
rect 120778 293936 120783 293992
rect 113173 293934 120783 293936
rect 113173 293931 113239 293934
rect 120717 293931 120783 293934
rect -960 293178 480 293268
rect 2773 293178 2839 293181
rect -960 293176 2839 293178
rect -960 293120 2778 293176
rect 2834 293120 2839 293176
rect -960 293118 2839 293120
rect -960 293028 480 293118
rect 2773 293115 2839 293118
rect 116577 293178 116643 293181
rect 126973 293178 127039 293181
rect 116577 293176 127039 293178
rect 116577 293120 116582 293176
rect 116638 293120 126978 293176
rect 127034 293120 127039 293176
rect 116577 293118 127039 293120
rect 116577 293115 116643 293118
rect 126973 293115 127039 293118
rect 105445 292770 105511 292773
rect 125041 292770 125107 292773
rect 105445 292768 125107 292770
rect 105445 292712 105450 292768
rect 105506 292712 125046 292768
rect 125102 292712 125107 292768
rect 105445 292710 125107 292712
rect 105445 292707 105511 292710
rect 125041 292707 125107 292710
rect 62614 292572 62620 292636
rect 62684 292634 62690 292636
rect 101581 292634 101647 292637
rect 62684 292632 101647 292634
rect 62684 292576 101586 292632
rect 101642 292576 101647 292632
rect 62684 292574 101647 292576
rect 62684 292572 62690 292574
rect 101581 292571 101647 292574
rect 104157 292634 104223 292637
rect 346393 292634 346459 292637
rect 104157 292632 346459 292634
rect 104157 292576 104162 292632
rect 104218 292576 346398 292632
rect 346454 292576 346459 292632
rect 104157 292574 346459 292576
rect 104157 292571 104223 292574
rect 346393 292571 346459 292574
rect 108205 291954 108271 291957
rect 335670 291954 335676 291956
rect 108205 291952 335676 291954
rect 108205 291896 108210 291952
rect 108266 291896 335676 291952
rect 108205 291894 335676 291896
rect 108205 291891 108271 291894
rect 335670 291892 335676 291894
rect 335740 291892 335746 291956
rect 121637 291818 121703 291821
rect 119876 291816 121703 291818
rect 69749 291274 69815 291277
rect 70166 291274 70226 291788
rect 119876 291760 121642 291816
rect 121698 291760 121703 291816
rect 119876 291758 121703 291760
rect 121637 291755 121703 291758
rect 69749 291272 70226 291274
rect 69749 291216 69754 291272
rect 69810 291216 70226 291272
rect 69749 291214 70226 291216
rect 345105 291274 345171 291277
rect 346158 291274 346164 291276
rect 345105 291272 346164 291274
rect 345105 291216 345110 291272
rect 345166 291216 346164 291272
rect 345105 291214 346164 291216
rect 69749 291211 69815 291214
rect 345105 291211 345171 291214
rect 346158 291212 346164 291214
rect 346228 291212 346234 291276
rect 67633 291138 67699 291141
rect 121729 291138 121795 291141
rect 67633 291136 70196 291138
rect 67633 291080 67638 291136
rect 67694 291080 70196 291136
rect 67633 291078 70196 291080
rect 119876 291136 121795 291138
rect 119876 291080 121734 291136
rect 121790 291080 121795 291136
rect 119876 291078 121795 291080
rect 67633 291075 67699 291078
rect 121729 291075 121795 291078
rect 119889 290594 119955 290597
rect 325693 290594 325759 290597
rect 119889 290592 325759 290594
rect 119889 290536 119894 290592
rect 119950 290536 325698 290592
rect 325754 290536 325759 290592
rect 119889 290534 325759 290536
rect 119889 290531 119955 290534
rect 325693 290531 325759 290534
rect 68829 290458 68895 290461
rect 121637 290458 121703 290461
rect 68829 290456 70196 290458
rect 68829 290400 68834 290456
rect 68890 290400 70196 290456
rect 68829 290398 70196 290400
rect 119876 290456 121703 290458
rect 119876 290400 121642 290456
rect 121698 290400 121703 290456
rect 119876 290398 121703 290400
rect 68829 290395 68895 290398
rect 121637 290395 121703 290398
rect 68737 289778 68803 289781
rect 121637 289778 121703 289781
rect 68737 289776 70196 289778
rect 68737 289720 68742 289776
rect 68798 289720 70196 289776
rect 68737 289718 70196 289720
rect 119876 289776 121703 289778
rect 119876 289720 121642 289776
rect 121698 289720 121703 289776
rect 119876 289718 121703 289720
rect 68737 289715 68803 289718
rect 121637 289715 121703 289718
rect 68185 289098 68251 289101
rect 121637 289098 121703 289101
rect 68185 289096 70196 289098
rect 68185 289040 68190 289096
rect 68246 289040 70196 289096
rect 68185 289038 70196 289040
rect 119876 289096 121703 289098
rect 119876 289040 121642 289096
rect 121698 289040 121703 289096
rect 119876 289038 121703 289040
rect 68185 289035 68251 289038
rect 121637 289035 121703 289038
rect 69105 288418 69171 288421
rect 121821 288418 121887 288421
rect 69105 288416 70196 288418
rect 69105 288360 69110 288416
rect 69166 288360 70196 288416
rect 69105 288358 70196 288360
rect 119876 288416 121887 288418
rect 119876 288360 121826 288416
rect 121882 288360 121887 288416
rect 119876 288358 121887 288360
rect 69105 288355 69171 288358
rect 121821 288355 121887 288358
rect 67633 287738 67699 287741
rect 122189 287738 122255 287741
rect 67633 287736 70196 287738
rect 67633 287680 67638 287736
rect 67694 287680 70196 287736
rect 67633 287678 70196 287680
rect 119876 287736 122255 287738
rect 119876 287680 122194 287736
rect 122250 287680 122255 287736
rect 119876 287678 122255 287680
rect 67633 287675 67699 287678
rect 122189 287675 122255 287678
rect 67725 287058 67791 287061
rect 121637 287058 121703 287061
rect 67725 287056 70196 287058
rect 67725 287000 67730 287056
rect 67786 287000 70196 287056
rect 67725 286998 70196 287000
rect 119876 287056 121703 287058
rect 119876 287000 121642 287056
rect 121698 287000 121703 287056
rect 119876 286998 121703 287000
rect 67725 286995 67791 286998
rect 121637 286995 121703 286998
rect 119797 286786 119863 286789
rect 119797 286784 119906 286786
rect 119797 286728 119802 286784
rect 119858 286728 119906 286784
rect 119797 286723 119906 286728
rect 67633 286378 67699 286381
rect 67633 286376 70196 286378
rect 67633 286320 67638 286376
rect 67694 286320 70196 286376
rect 119846 286348 119906 286723
rect 67633 286318 70196 286320
rect 67633 286315 67699 286318
rect 67449 285698 67515 285701
rect 121545 285698 121611 285701
rect 67449 285696 70196 285698
rect 67449 285640 67454 285696
rect 67510 285640 70196 285696
rect 67449 285638 70196 285640
rect 119876 285696 121611 285698
rect 119876 285640 121550 285696
rect 121606 285640 121611 285696
rect 119876 285638 121611 285640
rect 67449 285635 67515 285638
rect 121545 285635 121611 285638
rect 583520 285276 584960 285516
rect 121545 285018 121611 285021
rect 119876 285016 121611 285018
rect 64638 284412 64644 284476
rect 64708 284474 64714 284476
rect 70166 284474 70226 284988
rect 119876 284960 121550 285016
rect 121606 284960 121611 285016
rect 119876 284958 121611 284960
rect 121545 284955 121611 284958
rect 64708 284414 70226 284474
rect 64708 284412 64714 284414
rect 67633 284338 67699 284341
rect 121637 284338 121703 284341
rect 67633 284336 70196 284338
rect 67633 284280 67638 284336
rect 67694 284280 70196 284336
rect 67633 284278 70196 284280
rect 119876 284336 121703 284338
rect 119876 284280 121642 284336
rect 121698 284280 121703 284336
rect 119876 284278 121703 284280
rect 67633 284275 67699 284278
rect 121637 284275 121703 284278
rect 68829 283658 68895 283661
rect 121545 283658 121611 283661
rect 68829 283656 70196 283658
rect 68829 283600 68834 283656
rect 68890 283600 70196 283656
rect 68829 283598 70196 283600
rect 119876 283656 121611 283658
rect 119876 283600 121550 283656
rect 121606 283600 121611 283656
rect 119876 283598 121611 283600
rect 68829 283595 68895 283598
rect 121545 283595 121611 283598
rect 67541 282978 67607 282981
rect 121545 282978 121611 282981
rect 67541 282976 70196 282978
rect 67541 282920 67546 282976
rect 67602 282920 70196 282976
rect 67541 282918 70196 282920
rect 119876 282976 121611 282978
rect 119876 282920 121550 282976
rect 121606 282920 121611 282976
rect 119876 282918 121611 282920
rect 67541 282915 67607 282918
rect 121545 282915 121611 282918
rect 121545 282298 121611 282301
rect 119876 282296 121611 282298
rect 119876 282240 121550 282296
rect 121606 282240 121611 282296
rect 119876 282238 121611 282240
rect 121545 282235 121611 282238
rect 68553 281618 68619 281621
rect 122097 281618 122163 281621
rect 68553 281616 70196 281618
rect 68553 281560 68558 281616
rect 68614 281560 70196 281616
rect 68553 281558 70196 281560
rect 119876 281616 122163 281618
rect 119876 281560 122102 281616
rect 122158 281560 122163 281616
rect 119876 281558 122163 281560
rect 68553 281555 68619 281558
rect 122097 281555 122163 281558
rect 67633 280938 67699 280941
rect 121637 280938 121703 280941
rect 67633 280936 70196 280938
rect 67633 280880 67638 280936
rect 67694 280880 70196 280936
rect 67633 280878 70196 280880
rect 119876 280936 121703 280938
rect 119876 280880 121642 280936
rect 121698 280880 121703 280936
rect 119876 280878 121703 280880
rect 67633 280875 67699 280878
rect 121637 280875 121703 280878
rect 68369 280258 68435 280261
rect 121545 280258 121611 280261
rect 68369 280256 70196 280258
rect -960 279972 480 280212
rect 68369 280200 68374 280256
rect 68430 280200 70196 280256
rect 68369 280198 70196 280200
rect 119876 280256 121611 280258
rect 119876 280200 121550 280256
rect 121606 280200 121611 280256
rect 119876 280198 121611 280200
rect 68369 280195 68435 280198
rect 121545 280195 121611 280198
rect 120022 279652 120028 279716
rect 120092 279714 120098 279716
rect 580349 279714 580415 279717
rect 120092 279712 580415 279714
rect 120092 279656 580354 279712
rect 580410 279656 580415 279712
rect 120092 279654 580415 279656
rect 120092 279652 120098 279654
rect 580349 279651 580415 279654
rect 67633 279578 67699 279581
rect 121637 279578 121703 279581
rect 67633 279576 70196 279578
rect 67633 279520 67638 279576
rect 67694 279520 70196 279576
rect 67633 279518 70196 279520
rect 119876 279576 121703 279578
rect 119876 279520 121642 279576
rect 121698 279520 121703 279576
rect 119876 279518 121703 279520
rect 67633 279515 67699 279518
rect 121637 279515 121703 279518
rect 69013 278898 69079 278901
rect 121545 278898 121611 278901
rect 69013 278896 70196 278898
rect 69013 278840 69018 278896
rect 69074 278840 70196 278896
rect 69013 278838 70196 278840
rect 119876 278896 121611 278898
rect 119876 278840 121550 278896
rect 121606 278840 121611 278896
rect 119876 278838 121611 278840
rect 69013 278835 69079 278838
rect 121545 278835 121611 278838
rect 67725 278218 67791 278221
rect 121637 278218 121703 278221
rect 67725 278216 70196 278218
rect 67725 278160 67730 278216
rect 67786 278160 70196 278216
rect 67725 278158 70196 278160
rect 119876 278216 121703 278218
rect 119876 278160 121642 278216
rect 121698 278160 121703 278216
rect 119876 278158 121703 278160
rect 67725 278155 67791 278158
rect 121637 278155 121703 278158
rect 67633 277538 67699 277541
rect 121545 277538 121611 277541
rect 67633 277536 70196 277538
rect 67633 277480 67638 277536
rect 67694 277480 70196 277536
rect 67633 277478 70196 277480
rect 119876 277536 121611 277538
rect 119876 277480 121550 277536
rect 121606 277480 121611 277536
rect 119876 277478 121611 277480
rect 67633 277475 67699 277478
rect 121545 277475 121611 277478
rect 67725 276858 67791 276861
rect 121637 276858 121703 276861
rect 67725 276856 70196 276858
rect 67725 276800 67730 276856
rect 67786 276800 70196 276856
rect 67725 276798 70196 276800
rect 119876 276856 121703 276858
rect 119876 276800 121642 276856
rect 121698 276800 121703 276856
rect 119876 276798 121703 276800
rect 67725 276795 67791 276798
rect 121637 276795 121703 276798
rect 67633 276178 67699 276181
rect 121545 276178 121611 276181
rect 67633 276176 70196 276178
rect 67633 276120 67638 276176
rect 67694 276120 70196 276176
rect 67633 276118 70196 276120
rect 119876 276176 121611 276178
rect 119876 276120 121550 276176
rect 121606 276120 121611 276176
rect 119876 276118 121611 276120
rect 67633 276115 67699 276118
rect 121545 276115 121611 276118
rect 67725 275498 67791 275501
rect 121729 275498 121795 275501
rect 67725 275496 70196 275498
rect 67725 275440 67730 275496
rect 67786 275440 70196 275496
rect 67725 275438 70196 275440
rect 119876 275496 121795 275498
rect 119876 275440 121734 275496
rect 121790 275440 121795 275496
rect 119876 275438 121795 275440
rect 67725 275435 67791 275438
rect 121729 275435 121795 275438
rect 67633 274818 67699 274821
rect 121545 274818 121611 274821
rect 67633 274816 70196 274818
rect 67633 274760 67638 274816
rect 67694 274760 70196 274816
rect 67633 274758 70196 274760
rect 119876 274816 121611 274818
rect 119876 274760 121550 274816
rect 121606 274760 121611 274816
rect 119876 274758 121611 274760
rect 67633 274755 67699 274758
rect 121545 274755 121611 274758
rect 67633 274138 67699 274141
rect 121637 274138 121703 274141
rect 67633 274136 70196 274138
rect 67633 274080 67638 274136
rect 67694 274080 70196 274136
rect 67633 274078 70196 274080
rect 119876 274136 121703 274138
rect 119876 274080 121642 274136
rect 121698 274080 121703 274136
rect 119876 274078 121703 274080
rect 67633 274075 67699 274078
rect 121637 274075 121703 274078
rect 68001 273458 68067 273461
rect 121545 273458 121611 273461
rect 68001 273456 70196 273458
rect 68001 273400 68006 273456
rect 68062 273400 70196 273456
rect 68001 273398 70196 273400
rect 119876 273456 121611 273458
rect 119876 273400 121550 273456
rect 121606 273400 121611 273456
rect 119876 273398 121611 273400
rect 68001 273395 68067 273398
rect 121545 273395 121611 273398
rect 67817 272778 67883 272781
rect 121637 272778 121703 272781
rect 67817 272776 70196 272778
rect 67817 272720 67822 272776
rect 67878 272720 70196 272776
rect 67817 272718 70196 272720
rect 119876 272776 121703 272778
rect 119876 272720 121642 272776
rect 121698 272720 121703 272776
rect 119876 272718 121703 272720
rect 67817 272715 67883 272718
rect 121637 272715 121703 272718
rect 580441 272234 580507 272237
rect 583520 272234 584960 272324
rect 580441 272232 584960 272234
rect 580441 272176 580446 272232
rect 580502 272176 584960 272232
rect 580441 272174 584960 272176
rect 580441 272171 580507 272174
rect 67633 272098 67699 272101
rect 67633 272096 70196 272098
rect 67633 272040 67638 272096
rect 67694 272040 70196 272096
rect 67633 272038 70196 272040
rect 119876 272038 122850 272098
rect 583520 272084 584960 272174
rect 67633 272035 67699 272038
rect 122790 271962 122850 272038
rect 173934 271962 173940 271964
rect 122790 271902 173940 271962
rect 173934 271900 173940 271902
rect 174004 271900 174010 271964
rect 67633 271418 67699 271421
rect 121545 271418 121611 271421
rect 67633 271416 70196 271418
rect 67633 271360 67638 271416
rect 67694 271360 70196 271416
rect 67633 271358 70196 271360
rect 119876 271416 121611 271418
rect 119876 271360 121550 271416
rect 121606 271360 121611 271416
rect 119876 271358 121611 271360
rect 67633 271355 67699 271358
rect 121545 271355 121611 271358
rect 67725 270738 67791 270741
rect 67725 270736 70196 270738
rect 67725 270680 67730 270736
rect 67786 270680 70196 270736
rect 67725 270678 70196 270680
rect 67725 270675 67791 270678
rect 67633 270058 67699 270061
rect 121637 270058 121703 270061
rect 67633 270056 70196 270058
rect 67633 270000 67638 270056
rect 67694 270000 70196 270056
rect 67633 269998 70196 270000
rect 119876 270056 121703 270058
rect 119876 270000 121642 270056
rect 121698 270000 121703 270056
rect 119876 269998 121703 270000
rect 67633 269995 67699 269998
rect 121637 269995 121703 269998
rect 68277 269378 68343 269381
rect 121545 269378 121611 269381
rect 68277 269376 70196 269378
rect 68277 269320 68282 269376
rect 68338 269320 70196 269376
rect 68277 269318 70196 269320
rect 119876 269376 121611 269378
rect 119876 269320 121550 269376
rect 121606 269320 121611 269376
rect 119876 269318 121611 269320
rect 68277 269315 68343 269318
rect 121545 269315 121611 269318
rect 67541 268698 67607 268701
rect 121821 268698 121887 268701
rect 67541 268696 70196 268698
rect 67541 268640 67546 268696
rect 67602 268640 70196 268696
rect 67541 268638 70196 268640
rect 119876 268696 121887 268698
rect 119876 268640 121826 268696
rect 121882 268640 121887 268696
rect 119876 268638 121887 268640
rect 67541 268635 67607 268638
rect 121821 268635 121887 268638
rect 67633 268018 67699 268021
rect 121545 268018 121611 268021
rect 67633 268016 70196 268018
rect 67633 267960 67638 268016
rect 67694 267960 70196 268016
rect 67633 267958 70196 267960
rect 119876 268016 121611 268018
rect 119876 267960 121550 268016
rect 121606 267960 121611 268016
rect 119876 267958 121611 267960
rect 67633 267955 67699 267958
rect 121545 267955 121611 267958
rect 67633 267338 67699 267341
rect 121453 267338 121519 267341
rect 67633 267336 70196 267338
rect -960 267202 480 267292
rect 67633 267280 67638 267336
rect 67694 267280 70196 267336
rect 67633 267278 70196 267280
rect 119876 267336 121519 267338
rect 119876 267280 121458 267336
rect 121514 267280 121519 267336
rect 119876 267278 121519 267280
rect 67633 267275 67699 267278
rect 121453 267275 121519 267278
rect 3509 267202 3575 267205
rect -960 267200 3575 267202
rect -960 267144 3514 267200
rect 3570 267144 3575 267200
rect -960 267142 3575 267144
rect -960 267052 480 267142
rect 3509 267139 3575 267142
rect 67725 266658 67791 266661
rect 122189 266658 122255 266661
rect 67725 266656 70196 266658
rect 67725 266600 67730 266656
rect 67786 266600 70196 266656
rect 67725 266598 70196 266600
rect 119876 266656 122255 266658
rect 119876 266600 122194 266656
rect 122250 266600 122255 266656
rect 119876 266598 122255 266600
rect 67725 266595 67791 266598
rect 122189 266595 122255 266598
rect 67817 265978 67883 265981
rect 121545 265978 121611 265981
rect 67817 265976 70196 265978
rect 67817 265920 67822 265976
rect 67878 265920 70196 265976
rect 67817 265918 70196 265920
rect 119876 265976 121611 265978
rect 119876 265920 121550 265976
rect 121606 265920 121611 265976
rect 119876 265918 121611 265920
rect 67817 265915 67883 265918
rect 121545 265915 121611 265918
rect 67633 265298 67699 265301
rect 121453 265298 121519 265301
rect 67633 265296 70196 265298
rect 67633 265240 67638 265296
rect 67694 265240 70196 265296
rect 67633 265238 70196 265240
rect 119876 265296 121519 265298
rect 119876 265240 121458 265296
rect 121514 265240 121519 265296
rect 119876 265238 121519 265240
rect 67633 265235 67699 265238
rect 121453 265235 121519 265238
rect 67725 264618 67791 264621
rect 121453 264618 121519 264621
rect 67725 264616 70196 264618
rect 67725 264560 67730 264616
rect 67786 264560 70196 264616
rect 67725 264558 70196 264560
rect 119876 264616 121519 264618
rect 119876 264560 121458 264616
rect 121514 264560 121519 264616
rect 119876 264558 121519 264560
rect 67725 264555 67791 264558
rect 121453 264555 121519 264558
rect 120022 264148 120028 264212
rect 120092 264210 120098 264212
rect 580441 264210 580507 264213
rect 120092 264208 580507 264210
rect 120092 264152 580446 264208
rect 580502 264152 580507 264208
rect 120092 264150 580507 264152
rect 120092 264148 120098 264150
rect 580441 264147 580507 264150
rect 67633 263938 67699 263941
rect 121453 263938 121519 263941
rect 67633 263936 70196 263938
rect 67633 263880 67638 263936
rect 67694 263880 70196 263936
rect 67633 263878 70196 263880
rect 119876 263936 121519 263938
rect 119876 263880 121458 263936
rect 121514 263880 121519 263936
rect 119876 263878 121519 263880
rect 67633 263875 67699 263878
rect 121453 263875 121519 263878
rect 67633 263258 67699 263261
rect 121637 263258 121703 263261
rect 67633 263256 70196 263258
rect 67633 263200 67638 263256
rect 67694 263200 70196 263256
rect 67633 263198 70196 263200
rect 119876 263256 121703 263258
rect 119876 263200 121642 263256
rect 121698 263200 121703 263256
rect 119876 263198 121703 263200
rect 67633 263195 67699 263198
rect 121637 263195 121703 263198
rect 67633 262578 67699 262581
rect 121453 262578 121519 262581
rect 67633 262576 70196 262578
rect 67633 262520 67638 262576
rect 67694 262520 70196 262576
rect 67633 262518 70196 262520
rect 119876 262576 121519 262578
rect 119876 262520 121458 262576
rect 121514 262520 121519 262576
rect 119876 262518 121519 262520
rect 67633 262515 67699 262518
rect 121453 262515 121519 262518
rect 67725 261898 67791 261901
rect 121453 261898 121519 261901
rect 67725 261896 70196 261898
rect 67725 261840 67730 261896
rect 67786 261840 70196 261896
rect 67725 261838 70196 261840
rect 119876 261896 121519 261898
rect 119876 261840 121458 261896
rect 121514 261840 121519 261896
rect 119876 261838 121519 261840
rect 67725 261835 67791 261838
rect 121453 261835 121519 261838
rect 67357 261218 67423 261221
rect 120165 261218 120231 261221
rect 67357 261216 70196 261218
rect 67357 261160 67362 261216
rect 67418 261160 70196 261216
rect 67357 261158 70196 261160
rect 119876 261216 120231 261218
rect 119876 261160 120170 261216
rect 120226 261160 120231 261216
rect 119876 261158 120231 261160
rect 67357 261155 67423 261158
rect 120165 261155 120231 261158
rect 67633 260538 67699 260541
rect 67633 260536 70196 260538
rect 67633 260480 67638 260536
rect 67694 260480 70196 260536
rect 67633 260478 70196 260480
rect 67633 260475 67699 260478
rect 119846 259994 119906 260508
rect 119846 259934 122850 259994
rect 67633 259858 67699 259861
rect 121453 259858 121519 259861
rect 67633 259856 70196 259858
rect 67633 259800 67638 259856
rect 67694 259800 70196 259856
rect 67633 259798 70196 259800
rect 119876 259856 121519 259858
rect 119876 259800 121458 259856
rect 121514 259800 121519 259856
rect 119876 259798 121519 259800
rect 67633 259795 67699 259798
rect 121453 259795 121519 259798
rect 122790 259586 122850 259934
rect 337326 259586 337332 259588
rect 122790 259526 337332 259586
rect 337326 259524 337332 259526
rect 337396 259524 337402 259588
rect 67725 259178 67791 259181
rect 122097 259178 122163 259181
rect 67725 259176 70196 259178
rect 67725 259120 67730 259176
rect 67786 259120 70196 259176
rect 67725 259118 70196 259120
rect 119876 259176 122163 259178
rect 119876 259120 122102 259176
rect 122158 259120 122163 259176
rect 119876 259118 122163 259120
rect 67725 259115 67791 259118
rect 122097 259115 122163 259118
rect 579613 258906 579679 258909
rect 583520 258906 584960 258996
rect 579613 258904 584960 258906
rect 579613 258848 579618 258904
rect 579674 258848 584960 258904
rect 579613 258846 584960 258848
rect 579613 258843 579679 258846
rect 583520 258756 584960 258846
rect 67633 258498 67699 258501
rect 121453 258498 121519 258501
rect 67633 258496 70196 258498
rect 67633 258440 67638 258496
rect 67694 258440 70196 258496
rect 67633 258438 70196 258440
rect 119876 258496 121519 258498
rect 119876 258440 121458 258496
rect 121514 258440 121519 258496
rect 119876 258438 121519 258440
rect 67633 258435 67699 258438
rect 121453 258435 121519 258438
rect 67725 257818 67791 257821
rect 121637 257818 121703 257821
rect 67725 257816 70196 257818
rect 67725 257760 67730 257816
rect 67786 257760 70196 257816
rect 67725 257758 70196 257760
rect 119876 257816 121703 257818
rect 119876 257760 121642 257816
rect 121698 257760 121703 257816
rect 119876 257758 121703 257760
rect 67725 257755 67791 257758
rect 121637 257755 121703 257758
rect 67633 257138 67699 257141
rect 121453 257138 121519 257141
rect 67633 257136 70196 257138
rect 67633 257080 67638 257136
rect 67694 257080 70196 257136
rect 67633 257078 70196 257080
rect 119876 257136 121519 257138
rect 119876 257080 121458 257136
rect 121514 257080 121519 257136
rect 119876 257078 121519 257080
rect 67633 257075 67699 257078
rect 121453 257075 121519 257078
rect 67633 256458 67699 256461
rect 121453 256458 121519 256461
rect 67633 256456 70196 256458
rect 67633 256400 67638 256456
rect 67694 256400 70196 256456
rect 67633 256398 70196 256400
rect 119876 256456 121519 256458
rect 119876 256400 121458 256456
rect 121514 256400 121519 256456
rect 119876 256398 121519 256400
rect 67633 256395 67699 256398
rect 121453 256395 121519 256398
rect 67725 255778 67791 255781
rect 121545 255778 121611 255781
rect 67725 255776 70196 255778
rect 67725 255720 67730 255776
rect 67786 255720 70196 255776
rect 67725 255718 70196 255720
rect 119876 255776 121611 255778
rect 119876 255720 121550 255776
rect 121606 255720 121611 255776
rect 119876 255718 121611 255720
rect 67725 255715 67791 255718
rect 121545 255715 121611 255718
rect 67633 255098 67699 255101
rect 121545 255098 121611 255101
rect 67633 255096 70196 255098
rect 67633 255040 67638 255096
rect 67694 255040 70196 255096
rect 67633 255038 70196 255040
rect 119876 255096 121611 255098
rect 119876 255040 121550 255096
rect 121606 255040 121611 255096
rect 119876 255038 121611 255040
rect 67633 255035 67699 255038
rect 121545 255035 121611 255038
rect 121453 254418 121519 254421
rect 119876 254416 121519 254418
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 64454 254084 64460 254148
rect 64524 254146 64530 254148
rect 70166 254146 70226 254388
rect 119876 254360 121458 254416
rect 121514 254360 121519 254416
rect 119876 254358 121519 254360
rect 121453 254355 121519 254358
rect 64524 254086 70226 254146
rect 64524 254084 64530 254086
rect 67633 253738 67699 253741
rect 121545 253738 121611 253741
rect 67633 253736 70196 253738
rect 67633 253680 67638 253736
rect 67694 253680 70196 253736
rect 67633 253678 70196 253680
rect 119876 253736 121611 253738
rect 119876 253680 121550 253736
rect 121606 253680 121611 253736
rect 119876 253678 121611 253680
rect 67633 253675 67699 253678
rect 121545 253675 121611 253678
rect 68093 253058 68159 253061
rect 121453 253058 121519 253061
rect 68093 253056 70196 253058
rect 68093 253000 68098 253056
rect 68154 253000 70196 253056
rect 68093 252998 70196 253000
rect 119876 253056 121519 253058
rect 119876 253000 121458 253056
rect 121514 253000 121519 253056
rect 119876 252998 121519 253000
rect 68093 252995 68159 252998
rect 121453 252995 121519 252998
rect 121637 252378 121703 252381
rect 119876 252376 121703 252378
rect 70166 251834 70226 252348
rect 119876 252320 121642 252376
rect 121698 252320 121703 252376
rect 119876 252318 121703 252320
rect 121637 252315 121703 252318
rect 64830 251774 70226 251834
rect 63350 251364 63356 251428
rect 63420 251426 63426 251428
rect 64830 251426 64890 251774
rect 67449 251698 67515 251701
rect 121453 251698 121519 251701
rect 67449 251696 70196 251698
rect 67449 251640 67454 251696
rect 67510 251640 70196 251696
rect 67449 251638 70196 251640
rect 119876 251696 121519 251698
rect 119876 251640 121458 251696
rect 121514 251640 121519 251696
rect 119876 251638 121519 251640
rect 67449 251635 67515 251638
rect 121453 251635 121519 251638
rect 63420 251366 64890 251426
rect 63420 251364 63426 251366
rect 67633 251018 67699 251021
rect 120165 251018 120231 251021
rect 67633 251016 70196 251018
rect 67633 250960 67638 251016
rect 67694 250960 70196 251016
rect 67633 250958 70196 250960
rect 119876 251016 120231 251018
rect 119876 250960 120170 251016
rect 120226 250960 120231 251016
rect 119876 250958 120231 250960
rect 67633 250955 67699 250958
rect 120165 250955 120231 250958
rect 67725 250338 67791 250341
rect 121545 250338 121611 250341
rect 67725 250336 70196 250338
rect 67725 250280 67730 250336
rect 67786 250280 70196 250336
rect 67725 250278 70196 250280
rect 119876 250336 121611 250338
rect 119876 250280 121550 250336
rect 121606 250280 121611 250336
rect 119876 250278 121611 250280
rect 67725 250275 67791 250278
rect 121545 250275 121611 250278
rect 67633 249658 67699 249661
rect 121453 249658 121519 249661
rect 67633 249656 70196 249658
rect 67633 249600 67638 249656
rect 67694 249600 70196 249656
rect 67633 249598 70196 249600
rect 119876 249656 121519 249658
rect 119876 249600 121458 249656
rect 121514 249600 121519 249656
rect 119876 249598 121519 249600
rect 67633 249595 67699 249598
rect 121453 249595 121519 249598
rect 67633 248978 67699 248981
rect 121453 248978 121519 248981
rect 67633 248976 70196 248978
rect 67633 248920 67638 248976
rect 67694 248920 70196 248976
rect 67633 248918 70196 248920
rect 119876 248976 121519 248978
rect 119876 248920 121458 248976
rect 121514 248920 121519 248976
rect 119876 248918 121519 248920
rect 67633 248915 67699 248918
rect 121453 248915 121519 248918
rect 67633 248298 67699 248301
rect 121453 248298 121519 248301
rect 67633 248296 70196 248298
rect 67633 248240 67638 248296
rect 67694 248240 70196 248296
rect 67633 248238 70196 248240
rect 119876 248296 121519 248298
rect 119876 248240 121458 248296
rect 121514 248240 121519 248296
rect 119876 248238 121519 248240
rect 67633 248235 67699 248238
rect 121453 248235 121519 248238
rect 67725 247618 67791 247621
rect 120073 247618 120139 247621
rect 67725 247616 70196 247618
rect 67725 247560 67730 247616
rect 67786 247560 70196 247616
rect 67725 247558 70196 247560
rect 119876 247616 120139 247618
rect 119876 247560 120078 247616
rect 120134 247560 120139 247616
rect 119876 247558 120139 247560
rect 67725 247555 67791 247558
rect 120073 247555 120139 247558
rect 67633 246938 67699 246941
rect 121545 246938 121611 246941
rect 67633 246936 70196 246938
rect 67633 246880 67638 246936
rect 67694 246880 70196 246936
rect 67633 246878 70196 246880
rect 119876 246936 121611 246938
rect 119876 246880 121550 246936
rect 121606 246880 121611 246936
rect 119876 246878 121611 246880
rect 67633 246875 67699 246878
rect 121545 246875 121611 246878
rect 120717 246394 120783 246397
rect 120717 246392 122850 246394
rect 120717 246336 120722 246392
rect 120778 246336 122850 246392
rect 120717 246334 122850 246336
rect 120717 246331 120783 246334
rect 69013 246258 69079 246261
rect 121637 246258 121703 246261
rect 69013 246256 70196 246258
rect 69013 246200 69018 246256
rect 69074 246200 70196 246256
rect 69013 246198 70196 246200
rect 119876 246256 121703 246258
rect 119876 246200 121642 246256
rect 121698 246200 121703 246256
rect 119876 246198 121703 246200
rect 122790 246258 122850 246334
rect 580206 246258 580212 246260
rect 122790 246198 580212 246258
rect 69013 246195 69079 246198
rect 121637 246195 121703 246198
rect 580206 246196 580212 246198
rect 580276 246196 580282 246260
rect 66110 245652 66116 245716
rect 66180 245714 66186 245716
rect 68277 245714 68343 245717
rect 66180 245712 68343 245714
rect 66180 245656 68282 245712
rect 68338 245656 68343 245712
rect 66180 245654 68343 245656
rect 66180 245652 66186 245654
rect 68277 245651 68343 245654
rect 67633 245578 67699 245581
rect 121545 245578 121611 245581
rect 67633 245576 70196 245578
rect 67633 245520 67638 245576
rect 67694 245520 70196 245576
rect 67633 245518 70196 245520
rect 119876 245576 121611 245578
rect 119876 245520 121550 245576
rect 121606 245520 121611 245576
rect 119876 245518 121611 245520
rect 67633 245515 67699 245518
rect 121545 245515 121611 245518
rect 579889 245578 579955 245581
rect 583520 245578 584960 245668
rect 579889 245576 584960 245578
rect 579889 245520 579894 245576
rect 579950 245520 584960 245576
rect 579889 245518 584960 245520
rect 579889 245515 579955 245518
rect 583520 245428 584960 245518
rect 67633 244898 67699 244901
rect 121453 244898 121519 244901
rect 67633 244896 70196 244898
rect 67633 244840 67638 244896
rect 67694 244840 70196 244896
rect 67633 244838 70196 244840
rect 119876 244896 121519 244898
rect 119876 244840 121458 244896
rect 121514 244840 121519 244896
rect 119876 244838 121519 244840
rect 67633 244835 67699 244838
rect 121453 244835 121519 244838
rect 67817 244218 67883 244221
rect 121545 244218 121611 244221
rect 67817 244216 70196 244218
rect 67817 244160 67822 244216
rect 67878 244160 70196 244216
rect 67817 244158 70196 244160
rect 119876 244216 121611 244218
rect 119876 244160 121550 244216
rect 121606 244160 121611 244216
rect 119876 244158 121611 244160
rect 67817 244155 67883 244158
rect 121545 244155 121611 244158
rect 67725 243538 67791 243541
rect 121453 243538 121519 243541
rect 67725 243536 70196 243538
rect 67725 243480 67730 243536
rect 67786 243480 70196 243536
rect 67725 243478 70196 243480
rect 119876 243536 121519 243538
rect 119876 243480 121458 243536
rect 121514 243480 121519 243536
rect 119876 243478 121519 243480
rect 67725 243475 67791 243478
rect 121453 243475 121519 243478
rect 121637 243538 121703 243541
rect 260966 243538 260972 243540
rect 121637 243536 260972 243538
rect 121637 243480 121642 243536
rect 121698 243480 260972 243536
rect 121637 243478 260972 243480
rect 121637 243475 121703 243478
rect 260966 243476 260972 243478
rect 261036 243476 261042 243540
rect 67633 242858 67699 242861
rect 121453 242858 121519 242861
rect 67633 242856 70196 242858
rect 67633 242800 67638 242856
rect 67694 242800 70196 242856
rect 67633 242798 70196 242800
rect 119876 242856 121519 242858
rect 119876 242800 121458 242856
rect 121514 242800 121519 242856
rect 119876 242798 121519 242800
rect 67633 242795 67699 242798
rect 121453 242795 121519 242798
rect 67725 242178 67791 242181
rect 121545 242178 121611 242181
rect 67725 242176 70196 242178
rect 67725 242120 67730 242176
rect 67786 242120 70196 242176
rect 67725 242118 70196 242120
rect 119876 242176 121611 242178
rect 119876 242120 121550 242176
rect 121606 242120 121611 242176
rect 119876 242118 121611 242120
rect 67725 242115 67791 242118
rect 121545 242115 121611 242118
rect 67633 241498 67699 241501
rect 121453 241498 121519 241501
rect 67633 241496 70196 241498
rect 67633 241440 67638 241496
rect 67694 241440 70196 241496
rect 67633 241438 70196 241440
rect 119876 241496 121519 241498
rect 119876 241440 121458 241496
rect 121514 241440 121519 241496
rect 119876 241438 121519 241440
rect 67633 241435 67699 241438
rect 121453 241435 121519 241438
rect -960 241090 480 241180
rect 3049 241090 3115 241093
rect -960 241088 3115 241090
rect -960 241032 3054 241088
rect 3110 241032 3115 241088
rect -960 241030 3115 241032
rect -960 240940 480 241030
rect 3049 241027 3115 241030
rect 122097 240818 122163 240821
rect 119876 240816 122163 240818
rect 70534 239869 70594 240788
rect 119876 240760 122102 240816
rect 122158 240760 122163 240816
rect 119876 240758 122163 240760
rect 122097 240755 122163 240758
rect 121545 240138 121611 240141
rect 119876 240136 121611 240138
rect 119876 240080 121550 240136
rect 121606 240080 121611 240136
rect 119876 240078 121611 240080
rect 121545 240075 121611 240078
rect 70534 239864 70643 239869
rect 70534 239808 70582 239864
rect 70638 239808 70643 239864
rect 70534 239806 70643 239808
rect 70577 239803 70643 239806
rect 118325 238642 118391 238645
rect 120574 238642 120580 238644
rect 118325 238640 120580 238642
rect 118325 238584 118330 238640
rect 118386 238584 120580 238640
rect 118325 238582 120580 238584
rect 118325 238579 118391 238582
rect 120574 238580 120580 238582
rect 120644 238580 120650 238644
rect 91277 238506 91343 238509
rect 119654 238506 119660 238508
rect 91277 238504 119660 238506
rect 91277 238448 91282 238504
rect 91338 238448 119660 238504
rect 91277 238446 119660 238448
rect 91277 238443 91343 238446
rect 119654 238444 119660 238446
rect 119724 238444 119730 238508
rect 63350 236540 63356 236604
rect 63420 236602 63426 236604
rect 166257 236602 166323 236605
rect 63420 236600 166323 236602
rect 63420 236544 166262 236600
rect 166318 236544 166323 236600
rect 63420 236542 166323 236544
rect 63420 236540 63426 236542
rect 166257 236539 166323 236542
rect 54937 232522 55003 232525
rect 332542 232522 332548 232524
rect 54937 232520 332548 232522
rect 54937 232464 54942 232520
rect 54998 232464 332548 232520
rect 54937 232462 332548 232464
rect 54937 232459 55003 232462
rect 332542 232460 332548 232462
rect 332612 232460 332618 232524
rect 580441 232386 580507 232389
rect 583520 232386 584960 232476
rect 580441 232384 584960 232386
rect 580441 232328 580446 232384
rect 580502 232328 584960 232384
rect 580441 232326 584960 232328
rect 580441 232323 580507 232326
rect 583520 232236 584960 232326
rect 64454 231100 64460 231164
rect 64524 231162 64530 231164
rect 582833 231162 582899 231165
rect 64524 231160 582899 231162
rect 64524 231104 582838 231160
rect 582894 231104 582899 231160
rect 64524 231102 582899 231104
rect 64524 231100 64530 231102
rect 582833 231099 582899 231102
rect -960 227884 480 228124
rect 77109 224226 77175 224229
rect 329782 224226 329788 224228
rect 77109 224224 329788 224226
rect 77109 224168 77114 224224
rect 77170 224168 329788 224224
rect 77109 224166 329788 224168
rect 77109 224163 77175 224166
rect 329782 224164 329788 224166
rect 329852 224164 329858 224228
rect 84377 221506 84443 221509
rect 328494 221506 328500 221508
rect 84377 221504 328500 221506
rect 84377 221448 84382 221504
rect 84438 221448 328500 221504
rect 84377 221446 328500 221448
rect 84377 221443 84443 221446
rect 328494 221444 328500 221446
rect 328564 221444 328570 221508
rect 580349 219058 580415 219061
rect 583520 219058 584960 219148
rect 580349 219056 584960 219058
rect 580349 219000 580354 219056
rect 580410 219000 584960 219056
rect 580349 218998 584960 219000
rect 580349 218995 580415 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3509 214978 3575 214981
rect -960 214976 3575 214978
rect -960 214920 3514 214976
rect 3570 214920 3575 214976
rect -960 214918 3575 214920
rect -960 214828 480 214918
rect 3509 214915 3575 214918
rect 110413 214570 110479 214573
rect 248638 214570 248644 214572
rect 110413 214568 248644 214570
rect 110413 214512 110418 214568
rect 110474 214512 248644 214568
rect 110413 214510 248644 214512
rect 110413 214507 110479 214510
rect 248638 214508 248644 214510
rect 248708 214508 248714 214572
rect 55029 208994 55095 208997
rect 263726 208994 263732 208996
rect 55029 208992 263732 208994
rect 55029 208936 55034 208992
rect 55090 208936 263732 208992
rect 55029 208934 263732 208936
rect 55029 208931 55095 208934
rect 263726 208932 263732 208934
rect 263796 208932 263802 208996
rect 57789 207634 57855 207637
rect 265198 207634 265204 207636
rect 57789 207632 265204 207634
rect 57789 207576 57794 207632
rect 57850 207576 265204 207632
rect 57789 207574 265204 207576
rect 57789 207571 57855 207574
rect 265198 207572 265204 207574
rect 265268 207572 265274 207636
rect 46841 206274 46907 206277
rect 335670 206274 335676 206276
rect 46841 206272 335676 206274
rect 46841 206216 46846 206272
rect 46902 206216 335676 206272
rect 46841 206214 335676 206216
rect 46841 206211 46907 206214
rect 335670 206212 335676 206214
rect 335740 206212 335746 206276
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect 103605 204914 103671 204917
rect 327022 204914 327028 204916
rect 103605 204912 327028 204914
rect 103605 204856 103610 204912
rect 103666 204856 327028 204912
rect 103605 204854 327028 204856
rect 103605 204851 103671 204854
rect 327022 204852 327028 204854
rect 327092 204852 327098 204916
rect -960 201922 480 202012
rect 3049 201922 3115 201925
rect -960 201920 3115 201922
rect -960 201864 3054 201920
rect 3110 201864 3115 201920
rect -960 201862 3115 201864
rect -960 201772 480 201862
rect 3049 201859 3115 201862
rect 52361 197978 52427 197981
rect 338246 197978 338252 197980
rect 52361 197976 338252 197978
rect 52361 197920 52366 197976
rect 52422 197920 338252 197976
rect 52361 197918 338252 197920
rect 52361 197915 52427 197918
rect 338246 197916 338252 197918
rect 338316 197916 338322 197980
rect 152457 196618 152523 196621
rect 342294 196618 342300 196620
rect 152457 196616 342300 196618
rect 152457 196560 152462 196616
rect 152518 196560 342300 196616
rect 152457 196558 342300 196560
rect 152457 196555 152523 196558
rect 342294 196556 342300 196558
rect 342364 196556 342370 196620
rect 61837 193898 61903 193901
rect 263542 193898 263548 193900
rect 61837 193896 263548 193898
rect 61837 193840 61842 193896
rect 61898 193840 263548 193896
rect 61837 193838 263548 193840
rect 61837 193835 61903 193838
rect 263542 193836 263548 193838
rect 263612 193836 263618 193900
rect 583520 192538 584960 192628
rect 583342 192478 584960 192538
rect 583342 192402 583402 192478
rect 583520 192402 584960 192478
rect 583342 192388 584960 192402
rect 583342 192342 583586 192388
rect 64638 191796 64644 191860
rect 64708 191858 64714 191860
rect 583526 191858 583586 192342
rect 64708 191798 583586 191858
rect 64708 191796 64714 191798
rect 77293 189682 77359 189685
rect 327206 189682 327212 189684
rect 77293 189680 327212 189682
rect 77293 189624 77298 189680
rect 77354 189624 327212 189680
rect 77293 189622 327212 189624
rect 77293 189619 77359 189622
rect 327206 189620 327212 189622
rect 327276 189620 327282 189684
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 214557 188322 214623 188325
rect 259494 188322 259500 188324
rect 214557 188320 259500 188322
rect 214557 188264 214562 188320
rect 214618 188264 259500 188320
rect 214557 188262 259500 188264
rect 214557 188259 214623 188262
rect 259494 188260 259500 188262
rect 259564 188260 259570 188324
rect 73245 186962 73311 186965
rect 320214 186962 320220 186964
rect 73245 186960 320220 186962
rect 73245 186904 73250 186960
rect 73306 186904 320220 186960
rect 73245 186902 320220 186904
rect 73245 186899 73311 186902
rect 320214 186900 320220 186902
rect 320284 186900 320290 186964
rect 178677 184378 178743 184381
rect 256918 184378 256924 184380
rect 178677 184376 256924 184378
rect 178677 184320 178682 184376
rect 178738 184320 256924 184376
rect 178677 184318 256924 184320
rect 178677 184315 178743 184318
rect 256918 184316 256924 184318
rect 256988 184316 256994 184380
rect 60641 184242 60707 184245
rect 262254 184242 262260 184244
rect 60641 184240 262260 184242
rect 60641 184184 60646 184240
rect 60702 184184 262260 184240
rect 60641 184182 262260 184184
rect 60641 184179 60707 184182
rect 262254 184180 262260 184182
rect 262324 184180 262330 184244
rect 66110 182820 66116 182884
rect 66180 182882 66186 182884
rect 345289 182882 345355 182885
rect 66180 182880 345355 182882
rect 66180 182824 345294 182880
rect 345350 182824 345355 182880
rect 66180 182822 345355 182824
rect 66180 182820 66186 182822
rect 345289 182819 345355 182822
rect 300117 181386 300183 181389
rect 334014 181386 334020 181388
rect 300117 181384 334020 181386
rect 300117 181328 300122 181384
rect 300178 181328 334020 181384
rect 300117 181326 334020 181328
rect 300117 181323 300183 181326
rect 334014 181324 334020 181326
rect 334084 181324 334090 181388
rect 224309 180162 224375 180165
rect 257838 180162 257844 180164
rect 224309 180160 257844 180162
rect 224309 180104 224314 180160
rect 224370 180104 257844 180160
rect 224309 180102 257844 180104
rect 224309 180099 224375 180102
rect 257838 180100 257844 180102
rect 257908 180100 257914 180164
rect 189717 180026 189783 180029
rect 255262 180026 255268 180028
rect 189717 180024 255268 180026
rect 189717 179968 189722 180024
rect 189778 179968 255268 180024
rect 189717 179966 255268 179968
rect 189717 179963 189783 179966
rect 255262 179964 255268 179966
rect 255332 179964 255338 180028
rect 97349 179482 97415 179485
rect 167494 179482 167500 179484
rect 97349 179480 167500 179482
rect 97349 179424 97354 179480
rect 97410 179424 167500 179480
rect 97349 179422 167500 179424
rect 97349 179419 97415 179422
rect 167494 179420 167500 179422
rect 167564 179420 167570 179484
rect 579981 179210 580047 179213
rect 583520 179210 584960 179300
rect 579981 179208 584960 179210
rect 579981 179152 579986 179208
rect 580042 179152 584960 179208
rect 579981 179150 584960 179152
rect 579981 179147 580047 179150
rect 583520 179060 584960 179150
rect 305637 178802 305703 178805
rect 332726 178802 332732 178804
rect 305637 178800 332732 178802
rect 305637 178744 305642 178800
rect 305698 178744 332732 178800
rect 305637 178742 332732 178744
rect 305637 178739 305703 178742
rect 332726 178740 332732 178742
rect 332796 178740 332802 178804
rect 307109 178666 307175 178669
rect 336774 178666 336780 178668
rect 307109 178664 336780 178666
rect 307109 178608 307114 178664
rect 307170 178608 336780 178664
rect 307109 178606 336780 178608
rect 307109 178603 307175 178606
rect 336774 178604 336780 178606
rect 336844 178604 336850 178668
rect 99414 177516 99420 177580
rect 99484 177578 99490 177580
rect 100661 177578 100727 177581
rect 99484 177576 100727 177578
rect 99484 177520 100666 177576
rect 100722 177520 100727 177576
rect 99484 177518 100727 177520
rect 99484 177516 99490 177518
rect 100661 177515 100727 177518
rect 106038 177516 106044 177580
rect 106108 177578 106114 177580
rect 106181 177578 106247 177581
rect 106108 177576 106247 177578
rect 106108 177520 106186 177576
rect 106242 177520 106247 177576
rect 106108 177518 106247 177520
rect 106108 177516 106114 177518
rect 106181 177515 106247 177518
rect 106958 177516 106964 177580
rect 107028 177578 107034 177580
rect 107561 177578 107627 177581
rect 110689 177580 110755 177581
rect 112161 177580 112227 177581
rect 110638 177578 110644 177580
rect 107028 177576 107627 177578
rect 107028 177520 107566 177576
rect 107622 177520 107627 177576
rect 107028 177518 107627 177520
rect 110598 177518 110644 177578
rect 110708 177576 110755 177580
rect 112110 177578 112116 177580
rect 110750 177520 110755 177576
rect 107028 177516 107034 177518
rect 107561 177515 107627 177518
rect 110638 177516 110644 177518
rect 110708 177516 110755 177520
rect 112070 177518 112116 177578
rect 112180 177576 112227 177580
rect 112222 177520 112227 177576
rect 112110 177516 112116 177518
rect 112180 177516 112227 177520
rect 114134 177516 114140 177580
rect 114204 177578 114210 177580
rect 114369 177578 114435 177581
rect 114204 177576 114435 177578
rect 114204 177520 114374 177576
rect 114430 177520 114435 177576
rect 114204 177518 114435 177520
rect 114204 177516 114210 177518
rect 110689 177515 110755 177516
rect 112161 177515 112227 177516
rect 114369 177515 114435 177518
rect 116894 177516 116900 177580
rect 116964 177578 116970 177580
rect 117221 177578 117287 177581
rect 116964 177576 117287 177578
rect 116964 177520 117226 177576
rect 117282 177520 117287 177576
rect 116964 177518 117287 177520
rect 116964 177516 116970 177518
rect 117221 177515 117287 177518
rect 118366 177516 118372 177580
rect 118436 177578 118442 177580
rect 118601 177578 118667 177581
rect 118436 177576 118667 177578
rect 118436 177520 118606 177576
rect 118662 177520 118667 177576
rect 118436 177518 118667 177520
rect 118436 177516 118442 177518
rect 118601 177515 118667 177518
rect 122966 177516 122972 177580
rect 123036 177578 123042 177580
rect 124121 177578 124187 177581
rect 123036 177576 124187 177578
rect 123036 177520 124126 177576
rect 124182 177520 124187 177576
rect 123036 177518 124187 177520
rect 123036 177516 123042 177518
rect 124121 177515 124187 177518
rect 124438 177516 124444 177580
rect 124508 177578 124514 177580
rect 125041 177578 125107 177581
rect 124508 177576 125107 177578
rect 124508 177520 125046 177576
rect 125102 177520 125107 177576
rect 124508 177518 125107 177520
rect 124508 177516 124514 177518
rect 125041 177515 125107 177518
rect 125726 177516 125732 177580
rect 125796 177578 125802 177580
rect 126789 177578 126855 177581
rect 125796 177576 126855 177578
rect 125796 177520 126794 177576
rect 126850 177520 126855 177576
rect 125796 177518 126855 177520
rect 125796 177516 125802 177518
rect 126789 177515 126855 177518
rect 248413 177578 248479 177581
rect 249374 177578 249380 177580
rect 248413 177576 249380 177578
rect 248413 177520 248418 177576
rect 248474 177520 249380 177576
rect 248413 177518 249380 177520
rect 248413 177515 248479 177518
rect 249374 177516 249380 177518
rect 249444 177516 249450 177580
rect 313917 177306 313983 177309
rect 331438 177306 331444 177308
rect 313917 177304 331444 177306
rect 313917 177248 313922 177304
rect 313978 177248 331444 177304
rect 313917 177246 331444 177248
rect 313917 177243 313983 177246
rect 331438 177244 331444 177246
rect 331508 177244 331514 177308
rect 120758 177108 120764 177172
rect 120828 177170 120834 177172
rect 121177 177170 121243 177173
rect 133137 177172 133203 177173
rect 133086 177170 133092 177172
rect 120828 177168 121243 177170
rect 120828 177112 121182 177168
rect 121238 177112 121243 177168
rect 120828 177110 121243 177112
rect 133046 177110 133092 177170
rect 133156 177168 133203 177172
rect 133198 177112 133203 177168
rect 120828 177108 120834 177110
rect 121177 177107 121243 177110
rect 133086 177108 133092 177110
rect 133156 177108 133203 177112
rect 133137 177107 133203 177108
rect 103278 176972 103284 177036
rect 103348 177034 103354 177036
rect 167678 177034 167684 177036
rect 103348 176974 167684 177034
rect 103348 176972 103354 176974
rect 167678 176972 167684 176974
rect 167748 176972 167754 177036
rect 97022 176836 97028 176900
rect 97092 176898 97098 176900
rect 97349 176898 97415 176901
rect 97092 176896 97415 176898
rect 97092 176840 97354 176896
rect 97410 176840 97415 176896
rect 97092 176838 97415 176840
rect 97092 176836 97098 176838
rect 97349 176835 97415 176838
rect 104566 176836 104572 176900
rect 104636 176898 104642 176900
rect 166206 176898 166212 176900
rect 104636 176838 166212 176898
rect 104636 176836 104642 176838
rect 166206 176836 166212 176838
rect 166276 176836 166282 176900
rect 98310 176700 98316 176764
rect 98380 176762 98386 176764
rect 99097 176762 99163 176765
rect 102041 176764 102107 176765
rect 108113 176764 108179 176765
rect 101990 176762 101996 176764
rect 98380 176760 99163 176762
rect 98380 176704 99102 176760
rect 99158 176704 99163 176760
rect 98380 176702 99163 176704
rect 101950 176702 101996 176762
rect 102060 176760 102107 176764
rect 108062 176762 108068 176764
rect 102102 176704 102107 176760
rect 98380 176700 98386 176702
rect 99097 176699 99163 176702
rect 101990 176700 101996 176702
rect 102060 176700 102107 176704
rect 108022 176702 108068 176762
rect 108132 176760 108179 176764
rect 108174 176704 108179 176760
rect 108062 176700 108068 176702
rect 108132 176700 108179 176704
rect 109534 176700 109540 176764
rect 109604 176762 109610 176764
rect 110045 176762 110111 176765
rect 115841 176764 115907 176765
rect 127065 176764 127131 176765
rect 115790 176762 115796 176764
rect 109604 176760 110111 176762
rect 109604 176704 110050 176760
rect 110106 176704 110111 176760
rect 109604 176702 110111 176704
rect 115750 176702 115796 176762
rect 115860 176760 115907 176764
rect 127014 176762 127020 176764
rect 115902 176704 115907 176760
rect 109604 176700 109610 176702
rect 102041 176699 102107 176700
rect 108113 176699 108179 176700
rect 110045 176699 110111 176702
rect 115790 176700 115796 176702
rect 115860 176700 115907 176704
rect 126974 176702 127020 176762
rect 127084 176760 127131 176764
rect 128169 176762 128235 176765
rect 129457 176764 129523 176765
rect 132033 176764 132099 176765
rect 129406 176762 129412 176764
rect 127126 176704 127131 176760
rect 127014 176700 127020 176702
rect 127084 176700 127131 176704
rect 115841 176699 115907 176700
rect 127065 176699 127131 176700
rect 128126 176760 128235 176762
rect 128126 176704 128174 176760
rect 128230 176704 128235 176760
rect 128126 176699 128235 176704
rect 129366 176702 129412 176762
rect 129476 176760 129523 176764
rect 131982 176762 131988 176764
rect 129518 176704 129523 176760
rect 129406 176700 129412 176702
rect 129476 176700 129523 176704
rect 131942 176702 131988 176762
rect 132052 176760 132099 176764
rect 132094 176704 132099 176760
rect 131982 176700 131988 176702
rect 132052 176700 132099 176704
rect 134374 176700 134380 176764
rect 134444 176762 134450 176764
rect 134701 176762 134767 176765
rect 135713 176764 135779 176765
rect 148225 176764 148291 176765
rect 135662 176762 135668 176764
rect 134444 176760 134767 176762
rect 134444 176704 134706 176760
rect 134762 176704 134767 176760
rect 134444 176702 134767 176704
rect 135622 176702 135668 176762
rect 135732 176760 135779 176764
rect 148174 176762 148180 176764
rect 135774 176704 135779 176760
rect 134444 176700 134450 176702
rect 129457 176699 129523 176700
rect 132033 176699 132099 176700
rect 134701 176699 134767 176702
rect 135662 176700 135668 176702
rect 135732 176700 135779 176704
rect 148134 176702 148180 176762
rect 148244 176760 148291 176764
rect 148286 176704 148291 176760
rect 148174 176700 148180 176702
rect 148244 176700 148291 176704
rect 260046 176700 260052 176764
rect 260116 176762 260122 176764
rect 316033 176762 316099 176765
rect 260116 176760 316099 176762
rect 260116 176704 316038 176760
rect 316094 176704 316099 176760
rect 260116 176702 316099 176704
rect 260116 176700 260122 176702
rect 135713 176699 135779 176700
rect 148225 176699 148291 176700
rect 316033 176699 316099 176702
rect 320173 176762 320239 176765
rect 321318 176762 321324 176764
rect 320173 176760 321324 176762
rect 320173 176704 320178 176760
rect 320234 176704 321324 176760
rect 320173 176702 321324 176704
rect 320173 176699 320239 176702
rect 321318 176700 321324 176702
rect 321388 176700 321394 176764
rect 128126 176492 128186 176699
rect 319437 176626 319503 176629
rect 325877 176626 325943 176629
rect 319437 176624 325943 176626
rect 319437 176568 319442 176624
rect 319498 176568 325882 176624
rect 325938 176568 325943 176624
rect 319437 176566 325943 176568
rect 319437 176563 319503 176566
rect 325877 176563 325943 176566
rect 128118 176428 128124 176492
rect 128188 176428 128194 176492
rect 321502 176218 321508 176220
rect 315990 176158 321508 176218
rect 240777 176082 240843 176085
rect 249742 176082 249748 176084
rect 240777 176080 249748 176082
rect -960 175796 480 176036
rect 240777 176024 240782 176080
rect 240838 176024 249748 176080
rect 240777 176022 249748 176024
rect 240777 176019 240843 176022
rect 249742 176020 249748 176022
rect 249812 176020 249818 176084
rect 210417 175946 210483 175949
rect 256969 175946 257035 175949
rect 210417 175944 257035 175946
rect 210417 175888 210422 175944
rect 210478 175888 256974 175944
rect 257030 175888 257035 175944
rect 210417 175886 257035 175888
rect 210417 175883 210483 175886
rect 256969 175883 257035 175886
rect 312537 175946 312603 175949
rect 315990 175946 316050 176158
rect 321502 176156 321508 176158
rect 321572 176156 321578 176220
rect 321461 176082 321527 176085
rect 321461 176080 321570 176082
rect 321461 176024 321466 176080
rect 321522 176024 321570 176080
rect 321461 176019 321570 176024
rect 312537 175944 316050 175946
rect 312537 175888 312542 175944
rect 312598 175888 316050 175944
rect 312537 175886 316050 175888
rect 312537 175883 312603 175886
rect 248045 175810 248111 175813
rect 248045 175808 248338 175810
rect 248045 175752 248050 175808
rect 248106 175752 248338 175808
rect 248045 175750 248338 175752
rect 248045 175747 248111 175750
rect 213913 175674 213979 175677
rect 213913 175672 217212 175674
rect 213913 175616 213918 175672
rect 213974 175616 217212 175672
rect 248278 175644 248338 175750
rect 213913 175614 217212 175616
rect 213913 175611 213979 175614
rect 306966 175612 306972 175676
rect 307036 175674 307042 175676
rect 307036 175614 310132 175674
rect 307036 175612 307042 175614
rect 130745 175540 130811 175541
rect 158897 175540 158963 175541
rect 113214 175476 113220 175540
rect 113284 175538 113290 175540
rect 130694 175538 130700 175540
rect 113284 175478 122850 175538
rect 130654 175478 130700 175538
rect 130764 175536 130811 175540
rect 158846 175538 158852 175540
rect 130806 175480 130811 175536
rect 113284 175476 113290 175478
rect 100753 175404 100819 175405
rect 121913 175404 121979 175405
rect 100702 175402 100708 175404
rect 100662 175342 100708 175402
rect 100772 175400 100819 175404
rect 121862 175402 121868 175404
rect 100814 175344 100819 175400
rect 100702 175340 100708 175342
rect 100772 175340 100819 175344
rect 121822 175342 121868 175402
rect 121932 175400 121979 175404
rect 121974 175344 121979 175400
rect 121862 175340 121868 175342
rect 121932 175340 121979 175344
rect 122790 175402 122850 175478
rect 130694 175476 130700 175478
rect 130764 175476 130811 175480
rect 158806 175478 158852 175538
rect 158916 175536 158963 175540
rect 158958 175480 158963 175536
rect 321510 175508 321570 176019
rect 158846 175476 158852 175478
rect 158916 175476 158963 175480
rect 130745 175475 130811 175476
rect 158897 175475 158963 175476
rect 166390 175402 166396 175404
rect 122790 175342 166396 175402
rect 166390 175340 166396 175342
rect 166460 175340 166466 175404
rect 100753 175339 100819 175340
rect 121913 175339 121979 175340
rect 249241 175266 249307 175269
rect 248860 175264 249307 175266
rect 248860 175208 249246 175264
rect 249302 175208 249307 175264
rect 248860 175206 249307 175208
rect 249241 175203 249307 175206
rect 307017 175266 307083 175269
rect 321461 175266 321527 175269
rect 307017 175264 310132 175266
rect 307017 175208 307022 175264
rect 307078 175208 310132 175264
rect 307017 175206 310132 175208
rect 321461 175264 321570 175266
rect 321461 175208 321466 175264
rect 321522 175208 321570 175264
rect 307017 175203 307083 175206
rect 321461 175203 321570 175208
rect 119429 174996 119495 174997
rect 119392 174994 119398 174996
rect 119338 174934 119398 174994
rect 119462 174992 119495 174996
rect 119490 174936 119495 174992
rect 119392 174932 119398 174934
rect 119462 174932 119495 174936
rect 119429 174931 119495 174932
rect 213913 174994 213979 174997
rect 213913 174992 217212 174994
rect 213913 174936 213918 174992
rect 213974 174936 217212 174992
rect 213913 174934 217212 174936
rect 213913 174931 213979 174934
rect 306741 174858 306807 174861
rect 306741 174856 310132 174858
rect 306741 174800 306746 174856
rect 306802 174800 310132 174856
rect 306741 174798 310132 174800
rect 306741 174795 306807 174798
rect 249149 174722 249215 174725
rect 248860 174720 249215 174722
rect 248860 174664 249154 174720
rect 249210 174664 249215 174720
rect 321510 174692 321570 175203
rect 248860 174662 249215 174664
rect 249149 174659 249215 174662
rect 307661 174450 307727 174453
rect 307661 174448 310132 174450
rect 307661 174392 307666 174448
rect 307722 174392 310132 174448
rect 307661 174390 310132 174392
rect 307661 174387 307727 174390
rect 321502 174388 321508 174452
rect 321572 174388 321578 174452
rect 214005 174314 214071 174317
rect 249374 174314 249380 174316
rect 214005 174312 217212 174314
rect 214005 174256 214010 174312
rect 214066 174256 217212 174312
rect 214005 174254 217212 174256
rect 248860 174254 249380 174314
rect 214005 174251 214071 174254
rect 249374 174252 249380 174254
rect 249444 174252 249450 174316
rect 307569 174042 307635 174045
rect 307569 174040 310132 174042
rect 307569 173984 307574 174040
rect 307630 173984 310132 174040
rect 321510 174012 321570 174388
rect 307569 173982 310132 173984
rect 307569 173979 307635 173982
rect 249742 173770 249748 173772
rect 248860 173710 249748 173770
rect 249742 173708 249748 173710
rect 249812 173708 249818 173772
rect 321369 173770 321435 173773
rect 321369 173768 321570 173770
rect 321369 173712 321374 173768
rect 321430 173712 321570 173768
rect 321369 173710 321570 173712
rect 321369 173707 321435 173710
rect 213913 173634 213979 173637
rect 307661 173634 307727 173637
rect 213913 173632 217212 173634
rect 213913 173576 213918 173632
rect 213974 173576 217212 173632
rect 213913 173574 217212 173576
rect 307661 173632 310132 173634
rect 307661 173576 307666 173632
rect 307722 173576 310132 173632
rect 307661 173574 310132 173576
rect 213913 173571 213979 173574
rect 307661 173571 307727 173574
rect 251817 173362 251883 173365
rect 248860 173360 251883 173362
rect 248860 173304 251822 173360
rect 251878 173304 251883 173360
rect 248860 173302 251883 173304
rect 251817 173299 251883 173302
rect 306925 173226 306991 173229
rect 306925 173224 310132 173226
rect 306925 173168 306930 173224
rect 306986 173168 310132 173224
rect 321510 173196 321570 173710
rect 306925 173166 310132 173168
rect 306925 173163 306991 173166
rect 214097 172954 214163 172957
rect 214097 172952 217212 172954
rect 214097 172896 214102 172952
rect 214158 172896 217212 172952
rect 214097 172894 217212 172896
rect 214097 172891 214163 172894
rect 249149 172818 249215 172821
rect 248860 172816 249215 172818
rect 248860 172760 249154 172816
rect 249210 172760 249215 172816
rect 248860 172758 249215 172760
rect 249149 172755 249215 172758
rect 307293 172682 307359 172685
rect 321829 172682 321895 172685
rect 307293 172680 310132 172682
rect 307293 172624 307298 172680
rect 307354 172624 310132 172680
rect 307293 172622 310132 172624
rect 321829 172680 321938 172682
rect 321829 172624 321834 172680
rect 321890 172624 321938 172680
rect 307293 172619 307359 172622
rect 321829 172619 321938 172624
rect 252461 172410 252527 172413
rect 248860 172408 252527 172410
rect 248860 172352 252466 172408
rect 252522 172352 252527 172408
rect 321878 172380 321938 172619
rect 248860 172350 252527 172352
rect 252461 172347 252527 172350
rect 213913 172274 213979 172277
rect 307477 172274 307543 172277
rect 213913 172272 217212 172274
rect 213913 172216 213918 172272
rect 213974 172216 217212 172272
rect 213913 172214 217212 172216
rect 307477 172272 310132 172274
rect 307477 172216 307482 172272
rect 307538 172216 310132 172272
rect 307477 172214 310132 172216
rect 213913 172211 213979 172214
rect 307477 172211 307543 172214
rect 249793 171866 249859 171869
rect 248860 171864 249859 171866
rect 248860 171808 249798 171864
rect 249854 171808 249859 171864
rect 248860 171806 249859 171808
rect 249793 171803 249859 171806
rect 307569 171866 307635 171869
rect 307569 171864 310132 171866
rect 307569 171808 307574 171864
rect 307630 171808 310132 171864
rect 307569 171806 310132 171808
rect 307569 171803 307635 171806
rect 325877 171730 325943 171733
rect 321908 171728 325943 171730
rect 321908 171672 325882 171728
rect 325938 171672 325943 171728
rect 321908 171670 325943 171672
rect 325877 171667 325943 171670
rect 167637 171594 167703 171597
rect 164694 171592 167703 171594
rect 164694 171536 167642 171592
rect 167698 171536 167703 171592
rect 164694 171534 167703 171536
rect -960 162890 480 162980
rect 3233 162890 3299 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect -960 136778 480 136868
rect 3233 136778 3299 136781
rect -960 136776 3299 136778
rect -960 136720 3238 136776
rect 3294 136720 3299 136776
rect -960 136718 3299 136720
rect -960 136628 480 136718
rect 3233 136715 3299 136718
rect 167637 171531 167703 171534
rect 214005 171594 214071 171597
rect 214005 171592 217212 171594
rect 214005 171536 214010 171592
rect 214066 171536 217212 171592
rect 214005 171534 217212 171536
rect 214005 171531 214071 171534
rect 252001 171458 252067 171461
rect 248860 171456 252067 171458
rect 248860 171400 252006 171456
rect 252062 171400 252067 171456
rect 248860 171398 252067 171400
rect 252001 171395 252067 171398
rect 307661 171458 307727 171461
rect 307661 171456 310132 171458
rect 307661 171400 307666 171456
rect 307722 171400 310132 171456
rect 307661 171398 310132 171400
rect 307661 171395 307727 171398
rect 214005 171050 214071 171053
rect 306925 171050 306991 171053
rect 214005 171048 217212 171050
rect 214005 170992 214010 171048
rect 214066 170992 217212 171048
rect 214005 170990 217212 170992
rect 306925 171048 310132 171050
rect 306925 170992 306930 171048
rect 306986 170992 310132 171048
rect 306925 170990 310132 170992
rect 214005 170987 214071 170990
rect 306925 170987 306991 170990
rect 321318 170988 321324 171052
rect 321388 170988 321394 171052
rect 252461 170914 252527 170917
rect 248860 170912 252527 170914
rect 248860 170856 252466 170912
rect 252522 170856 252527 170912
rect 321326 170884 321386 170988
rect 248860 170854 252527 170856
rect 252461 170851 252527 170854
rect 307477 170642 307543 170645
rect 307477 170640 310132 170642
rect 307477 170584 307482 170640
rect 307538 170584 310132 170640
rect 307477 170582 310132 170584
rect 307477 170579 307543 170582
rect 251817 170506 251883 170509
rect 248860 170504 251883 170506
rect 248860 170448 251822 170504
rect 251878 170448 251883 170504
rect 248860 170446 251883 170448
rect 251817 170443 251883 170446
rect 213913 170370 213979 170373
rect 213913 170368 217212 170370
rect 213913 170312 213918 170368
rect 213974 170312 217212 170368
rect 213913 170310 217212 170312
rect 213913 170307 213979 170310
rect 321318 170308 321324 170372
rect 321388 170308 321394 170372
rect 307661 170234 307727 170237
rect 307661 170232 310132 170234
rect 307661 170176 307666 170232
rect 307722 170176 310132 170232
rect 307661 170174 310132 170176
rect 307661 170171 307727 170174
rect 252093 170098 252159 170101
rect 248860 170096 252159 170098
rect 248860 170040 252098 170096
rect 252154 170040 252159 170096
rect 321326 170068 321386 170308
rect 248860 170038 252159 170040
rect 252093 170035 252159 170038
rect 307201 169826 307267 169829
rect 307201 169824 310132 169826
rect 307201 169768 307206 169824
rect 307262 169768 310132 169824
rect 307201 169766 310132 169768
rect 307201 169763 307267 169766
rect 214005 169690 214071 169693
rect 214005 169688 217212 169690
rect 214005 169632 214010 169688
rect 214066 169632 217212 169688
rect 214005 169630 217212 169632
rect 214005 169627 214071 169630
rect 252645 169554 252711 169557
rect 248860 169552 252711 169554
rect 248860 169496 252650 169552
rect 252706 169496 252711 169552
rect 248860 169494 252711 169496
rect 252645 169491 252711 169494
rect 324313 169418 324379 169421
rect 321908 169416 324379 169418
rect 321908 169360 324318 169416
rect 324374 169360 324379 169416
rect 321908 169358 324379 169360
rect 324313 169355 324379 169358
rect 307477 169282 307543 169285
rect 307477 169280 310132 169282
rect 307477 169224 307482 169280
rect 307538 169224 310132 169280
rect 307477 169222 310132 169224
rect 307477 169219 307543 169222
rect 252461 169146 252527 169149
rect 248860 169144 252527 169146
rect 248860 169088 252466 169144
rect 252522 169088 252527 169144
rect 248860 169086 252527 169088
rect 252461 169083 252527 169086
rect 213913 169010 213979 169013
rect 213913 169008 217212 169010
rect 213913 168952 213918 169008
rect 213974 168952 217212 169008
rect 213913 168950 217212 168952
rect 213913 168947 213979 168950
rect 307661 168874 307727 168877
rect 307661 168872 310132 168874
rect 307661 168816 307666 168872
rect 307722 168816 310132 168872
rect 307661 168814 310132 168816
rect 307661 168811 307727 168814
rect 252001 168602 252067 168605
rect 324405 168602 324471 168605
rect 248860 168600 252067 168602
rect 248860 168544 252006 168600
rect 252062 168544 252067 168600
rect 248860 168542 252067 168544
rect 321908 168600 324471 168602
rect 321908 168544 324410 168600
rect 324466 168544 324471 168600
rect 321908 168542 324471 168544
rect 252001 168539 252067 168542
rect 324405 168539 324471 168542
rect 307293 168466 307359 168469
rect 307293 168464 310132 168466
rect 307293 168408 307298 168464
rect 307354 168408 310132 168464
rect 307293 168406 310132 168408
rect 307293 168403 307359 168406
rect 213913 168330 213979 168333
rect 213913 168328 217212 168330
rect 213913 168272 213918 168328
rect 213974 168272 217212 168328
rect 213913 168270 217212 168272
rect 213913 168267 213979 168270
rect 251909 168194 251975 168197
rect 248860 168192 251975 168194
rect 248860 168136 251914 168192
rect 251970 168136 251975 168192
rect 248860 168134 251975 168136
rect 251909 168131 251975 168134
rect 307477 168058 307543 168061
rect 307477 168056 310132 168058
rect 307477 168000 307482 168056
rect 307538 168000 310132 168056
rect 307477 167998 310132 168000
rect 307477 167995 307543 167998
rect 324313 167786 324379 167789
rect 321908 167784 324379 167786
rect 321908 167728 324318 167784
rect 324374 167728 324379 167784
rect 321908 167726 324379 167728
rect 324313 167723 324379 167726
rect 214005 167650 214071 167653
rect 252461 167650 252527 167653
rect 214005 167648 217212 167650
rect 214005 167592 214010 167648
rect 214066 167592 217212 167648
rect 214005 167590 217212 167592
rect 248860 167648 252527 167650
rect 248860 167592 252466 167648
rect 252522 167592 252527 167648
rect 248860 167590 252527 167592
rect 214005 167587 214071 167590
rect 252461 167587 252527 167590
rect 307569 167650 307635 167653
rect 307569 167648 310132 167650
rect 307569 167592 307574 167648
rect 307630 167592 310132 167648
rect 307569 167590 310132 167592
rect 307569 167587 307635 167590
rect 252093 167242 252159 167245
rect 248860 167240 252159 167242
rect 248860 167184 252098 167240
rect 252154 167184 252159 167240
rect 248860 167182 252159 167184
rect 252093 167179 252159 167182
rect 307661 167242 307727 167245
rect 307661 167240 310132 167242
rect 307661 167184 307666 167240
rect 307722 167184 310132 167240
rect 307661 167182 310132 167184
rect 307661 167179 307727 167182
rect 324405 167106 324471 167109
rect 321908 167104 324471 167106
rect 321908 167048 324410 167104
rect 324466 167048 324471 167104
rect 321908 167046 324471 167048
rect 324405 167043 324471 167046
rect 213913 166970 213979 166973
rect 213913 166968 217212 166970
rect 213913 166912 213918 166968
rect 213974 166912 217212 166968
rect 213913 166910 217212 166912
rect 213913 166907 213979 166910
rect 307661 166834 307727 166837
rect 307661 166832 310132 166834
rect 307661 166776 307666 166832
rect 307722 166776 310132 166832
rect 307661 166774 310132 166776
rect 307661 166771 307727 166774
rect 250161 166698 250227 166701
rect 248860 166696 250227 166698
rect 248860 166640 250166 166696
rect 250222 166640 250227 166696
rect 248860 166638 250227 166640
rect 250161 166635 250227 166638
rect 214005 166426 214071 166429
rect 307477 166426 307543 166429
rect 214005 166424 217212 166426
rect 214005 166368 214010 166424
rect 214066 166368 217212 166424
rect 214005 166366 217212 166368
rect 307477 166424 310132 166426
rect 307477 166368 307482 166424
rect 307538 166368 310132 166424
rect 307477 166366 310132 166368
rect 214005 166363 214071 166366
rect 307477 166363 307543 166366
rect 251817 166290 251883 166293
rect 324313 166290 324379 166293
rect 248860 166288 251883 166290
rect 248860 166232 251822 166288
rect 251878 166232 251883 166288
rect 248860 166230 251883 166232
rect 321908 166288 324379 166290
rect 321908 166232 324318 166288
rect 324374 166232 324379 166288
rect 321908 166230 324379 166232
rect 251817 166227 251883 166230
rect 324313 166227 324379 166230
rect 307293 165882 307359 165885
rect 583520 165882 584960 165972
rect 307293 165880 310132 165882
rect 307293 165824 307298 165880
rect 307354 165824 310132 165880
rect 307293 165822 310132 165824
rect 567150 165822 584960 165882
rect 307293 165819 307359 165822
rect 214649 165746 214715 165749
rect 252737 165746 252803 165749
rect 214649 165744 217212 165746
rect 214649 165688 214654 165744
rect 214710 165688 217212 165744
rect 214649 165686 217212 165688
rect 248860 165744 252803 165746
rect 248860 165688 252742 165744
rect 252798 165688 252803 165744
rect 248860 165686 252803 165688
rect 214649 165683 214715 165686
rect 252737 165683 252803 165686
rect 321645 165746 321711 165749
rect 321645 165744 321754 165746
rect 321645 165688 321650 165744
rect 321706 165688 321754 165744
rect 321645 165683 321754 165688
rect 337326 165684 337332 165748
rect 337396 165746 337402 165748
rect 567150 165746 567210 165822
rect 337396 165686 567210 165746
rect 583520 165732 584960 165822
rect 337396 165684 337402 165686
rect 307477 165474 307543 165477
rect 307477 165472 310132 165474
rect 307477 165416 307482 165472
rect 307538 165416 310132 165472
rect 321694 165444 321754 165683
rect 307477 165414 310132 165416
rect 307477 165411 307543 165414
rect 252461 165338 252527 165341
rect 248860 165336 252527 165338
rect 248860 165280 252466 165336
rect 252522 165280 252527 165336
rect 248860 165278 252527 165280
rect 252461 165275 252527 165278
rect 213913 165066 213979 165069
rect 306557 165066 306623 165069
rect 321277 165066 321343 165069
rect 213913 165064 217212 165066
rect 213913 165008 213918 165064
rect 213974 165008 217212 165064
rect 213913 165006 217212 165008
rect 306557 165064 310132 165066
rect 306557 165008 306562 165064
rect 306618 165008 310132 165064
rect 306557 165006 310132 165008
rect 321277 165064 321386 165066
rect 321277 165008 321282 165064
rect 321338 165008 321386 165064
rect 213913 165003 213979 165006
rect 306557 165003 306623 165006
rect 321277 165003 321386 165008
rect 252369 164794 252435 164797
rect 248860 164792 252435 164794
rect 248860 164736 252374 164792
rect 252430 164736 252435 164792
rect 321326 164764 321386 165003
rect 248860 164734 252435 164736
rect 252369 164731 252435 164734
rect 307661 164658 307727 164661
rect 307661 164656 310132 164658
rect 307661 164600 307666 164656
rect 307722 164600 310132 164656
rect 307661 164598 310132 164600
rect 307661 164595 307727 164598
rect 214005 164386 214071 164389
rect 251357 164386 251423 164389
rect 214005 164384 217212 164386
rect 214005 164328 214010 164384
rect 214066 164328 217212 164384
rect 214005 164326 217212 164328
rect 248860 164384 251423 164386
rect 248860 164328 251362 164384
rect 251418 164328 251423 164384
rect 248860 164326 251423 164328
rect 214005 164323 214071 164326
rect 251357 164323 251423 164326
rect 307569 164250 307635 164253
rect 307569 164248 310132 164250
rect 307569 164192 307574 164248
rect 307630 164192 310132 164248
rect 307569 164190 310132 164192
rect 307569 164187 307635 164190
rect 252461 163978 252527 163981
rect 324313 163978 324379 163981
rect 248860 163976 252527 163978
rect 248860 163920 252466 163976
rect 252522 163920 252527 163976
rect 248860 163918 252527 163920
rect 321908 163976 324379 163978
rect 321908 163920 324318 163976
rect 324374 163920 324379 163976
rect 321908 163918 324379 163920
rect 252461 163915 252527 163918
rect 324313 163915 324379 163918
rect 307477 163842 307543 163845
rect 307477 163840 310132 163842
rect 307477 163784 307482 163840
rect 307538 163784 310132 163840
rect 307477 163782 310132 163784
rect 307477 163779 307543 163782
rect 166390 163100 166396 163164
rect 166460 163162 166466 163164
rect 217182 163162 217242 163676
rect 263726 163434 263732 163436
rect 248860 163374 263732 163434
rect 263726 163372 263732 163374
rect 263796 163372 263802 163436
rect 307661 163434 307727 163437
rect 307661 163432 310132 163434
rect 307661 163376 307666 163432
rect 307722 163376 310132 163432
rect 307661 163374 310132 163376
rect 307661 163371 307727 163374
rect 324405 163162 324471 163165
rect 166460 163102 217242 163162
rect 321908 163160 324471 163162
rect 321908 163104 324410 163160
rect 324466 163104 324471 163160
rect 321908 163102 324471 163104
rect 166460 163100 166466 163102
rect 324405 163099 324471 163102
rect 213913 163026 213979 163029
rect 251357 163026 251423 163029
rect 213913 163024 217212 163026
rect 213913 162968 213918 163024
rect 213974 162968 217212 163024
rect 213913 162966 217212 162968
rect 248860 163024 251423 163026
rect 248860 162968 251362 163024
rect 251418 162968 251423 163024
rect 248860 162966 251423 162968
rect 213913 162963 213979 162966
rect 251357 162963 251423 162966
rect 307293 163026 307359 163029
rect 307293 163024 310132 163026
rect 307293 162968 307298 163024
rect 307354 162968 310132 163024
rect 307293 162966 310132 162968
rect 307293 162963 307359 162966
rect 252461 162482 252527 162485
rect 248860 162480 252527 162482
rect 248860 162424 252466 162480
rect 252522 162424 252527 162480
rect 248860 162422 252527 162424
rect 252461 162419 252527 162422
rect 307477 162482 307543 162485
rect 324313 162482 324379 162485
rect 307477 162480 310132 162482
rect 307477 162424 307482 162480
rect 307538 162424 310132 162480
rect 307477 162422 310132 162424
rect 321908 162480 324379 162482
rect 321908 162424 324318 162480
rect 324374 162424 324379 162480
rect 321908 162422 324379 162424
rect 307477 162419 307543 162422
rect 324313 162419 324379 162422
rect 213913 162346 213979 162349
rect 213913 162344 217212 162346
rect 213913 162288 213918 162344
rect 213974 162288 217212 162344
rect 213913 162286 217212 162288
rect 213913 162283 213979 162286
rect 265198 162074 265204 162076
rect 248860 162014 265204 162074
rect 265198 162012 265204 162014
rect 265268 162012 265274 162076
rect 307293 162074 307359 162077
rect 307293 162072 310132 162074
rect 307293 162016 307298 162072
rect 307354 162016 310132 162072
rect 307293 162014 310132 162016
rect 307293 162011 307359 162014
rect 214741 161802 214807 161805
rect 214741 161800 217212 161802
rect 214741 161744 214746 161800
rect 214802 161744 217212 161800
rect 214741 161742 217212 161744
rect 214741 161739 214807 161742
rect 307661 161666 307727 161669
rect 324405 161666 324471 161669
rect 307661 161664 310132 161666
rect 307661 161608 307666 161664
rect 307722 161608 310132 161664
rect 307661 161606 310132 161608
rect 321908 161664 324471 161666
rect 321908 161608 324410 161664
rect 324466 161608 324471 161664
rect 321908 161606 324471 161608
rect 307661 161603 307727 161606
rect 324405 161603 324471 161606
rect 252093 161530 252159 161533
rect 248860 161528 252159 161530
rect 248860 161472 252098 161528
rect 252154 161472 252159 161528
rect 248860 161470 252159 161472
rect 252093 161467 252159 161470
rect 307661 161258 307727 161261
rect 307661 161256 310132 161258
rect 307661 161200 307666 161256
rect 307722 161200 310132 161256
rect 307661 161198 310132 161200
rect 307661 161195 307727 161198
rect 213913 161122 213979 161125
rect 252093 161122 252159 161125
rect 213913 161120 217212 161122
rect 213913 161064 213918 161120
rect 213974 161064 217212 161120
rect 213913 161062 217212 161064
rect 248860 161120 252159 161122
rect 248860 161064 252098 161120
rect 252154 161064 252159 161120
rect 248860 161062 252159 161064
rect 213913 161059 213979 161062
rect 252093 161059 252159 161062
rect 306557 160850 306623 160853
rect 324681 160850 324747 160853
rect 306557 160848 310132 160850
rect 306557 160792 306562 160848
rect 306618 160792 310132 160848
rect 306557 160790 310132 160792
rect 321908 160848 324747 160850
rect 321908 160792 324686 160848
rect 324742 160792 324747 160848
rect 321908 160790 324747 160792
rect 306557 160787 306623 160790
rect 324681 160787 324747 160790
rect 252461 160578 252527 160581
rect 248860 160576 252527 160578
rect 248860 160520 252466 160576
rect 252522 160520 252527 160576
rect 248860 160518 252527 160520
rect 252461 160515 252527 160518
rect 214005 160442 214071 160445
rect 307109 160442 307175 160445
rect 214005 160440 217212 160442
rect 214005 160384 214010 160440
rect 214066 160384 217212 160440
rect 214005 160382 217212 160384
rect 307109 160440 310132 160442
rect 307109 160384 307114 160440
rect 307170 160384 310132 160440
rect 307109 160382 310132 160384
rect 214005 160379 214071 160382
rect 307109 160379 307175 160382
rect 252001 160170 252067 160173
rect 324313 160170 324379 160173
rect 248860 160168 252067 160170
rect 248860 160112 252006 160168
rect 252062 160112 252067 160168
rect 248860 160110 252067 160112
rect 321908 160168 324379 160170
rect 321908 160112 324318 160168
rect 324374 160112 324379 160168
rect 321908 160110 324379 160112
rect 252001 160107 252067 160110
rect 324313 160107 324379 160110
rect 306925 160034 306991 160037
rect 306925 160032 310132 160034
rect 306925 159976 306930 160032
rect 306986 159976 310132 160032
rect 306925 159974 310132 159976
rect 306925 159971 306991 159974
rect 214465 159762 214531 159765
rect 214465 159760 217212 159762
rect 214465 159704 214470 159760
rect 214526 159704 217212 159760
rect 214465 159702 217212 159704
rect 214465 159699 214531 159702
rect 251173 159626 251239 159629
rect 248860 159624 251239 159626
rect 248860 159568 251178 159624
rect 251234 159568 251239 159624
rect 248860 159566 251239 159568
rect 251173 159563 251239 159566
rect 307477 159626 307543 159629
rect 307477 159624 310132 159626
rect 307477 159568 307482 159624
rect 307538 159568 310132 159624
rect 307477 159566 310132 159568
rect 307477 159563 307543 159566
rect 324313 159354 324379 159357
rect 321908 159352 324379 159354
rect 321908 159296 324318 159352
rect 324374 159296 324379 159352
rect 321908 159294 324379 159296
rect 324313 159291 324379 159294
rect 252461 159218 252527 159221
rect 248860 159216 252527 159218
rect 248860 159160 252466 159216
rect 252522 159160 252527 159216
rect 248860 159158 252527 159160
rect 252461 159155 252527 159158
rect 307661 159082 307727 159085
rect 200070 159022 217212 159082
rect 307661 159080 310132 159082
rect 307661 159024 307666 159080
rect 307722 159024 310132 159080
rect 307661 159022 310132 159024
rect 166206 158884 166212 158948
rect 166276 158946 166282 158948
rect 200070 158946 200130 159022
rect 307661 159019 307727 159022
rect 166276 158886 200130 158946
rect 166276 158884 166282 158886
rect 251265 158810 251331 158813
rect 248860 158808 251331 158810
rect 248860 158752 251270 158808
rect 251326 158752 251331 158808
rect 248860 158750 251331 158752
rect 251265 158747 251331 158750
rect 306925 158674 306991 158677
rect 306925 158672 310132 158674
rect 306925 158616 306930 158672
rect 306986 158616 310132 158672
rect 306925 158614 310132 158616
rect 306925 158611 306991 158614
rect 324313 158538 324379 158541
rect 321908 158536 324379 158538
rect 321908 158480 324318 158536
rect 324374 158480 324379 158536
rect 321908 158478 324379 158480
rect 324313 158475 324379 158478
rect 217182 157858 217242 158372
rect 252461 158266 252527 158269
rect 248860 158264 252527 158266
rect 248860 158208 252466 158264
rect 252522 158208 252527 158264
rect 248860 158206 252527 158208
rect 252461 158203 252527 158206
rect 307477 158266 307543 158269
rect 307477 158264 310132 158266
rect 307477 158208 307482 158264
rect 307538 158208 310132 158264
rect 307477 158206 310132 158208
rect 307477 158203 307543 158206
rect 252369 157858 252435 157861
rect 200070 157798 217242 157858
rect 248860 157856 252435 157858
rect 248860 157800 252374 157856
rect 252430 157800 252435 157856
rect 248860 157798 252435 157800
rect 167678 157388 167684 157452
rect 167748 157450 167754 157452
rect 200070 157450 200130 157798
rect 252369 157795 252435 157798
rect 307293 157858 307359 157861
rect 324405 157858 324471 157861
rect 307293 157856 310132 157858
rect 307293 157800 307298 157856
rect 307354 157800 310132 157856
rect 307293 157798 310132 157800
rect 321908 157856 324471 157858
rect 321908 157800 324410 157856
rect 324466 157800 324471 157856
rect 321908 157798 324471 157800
rect 307293 157795 307359 157798
rect 324405 157795 324471 157798
rect 213913 157722 213979 157725
rect 213913 157720 217212 157722
rect 213913 157664 213918 157720
rect 213974 157664 217212 157720
rect 213913 157662 217212 157664
rect 213913 157659 213979 157662
rect 167748 157390 200130 157450
rect 307385 157450 307451 157453
rect 307385 157448 310132 157450
rect 307385 157392 307390 157448
rect 307446 157392 310132 157448
rect 307385 157390 310132 157392
rect 167748 157388 167754 157390
rect 307385 157387 307451 157390
rect 252461 157314 252527 157317
rect 248860 157312 252527 157314
rect 248860 157256 252466 157312
rect 252522 157256 252527 157312
rect 248860 157254 252527 157256
rect 252461 157251 252527 157254
rect 214005 157178 214071 157181
rect 214005 157176 217212 157178
rect 214005 157120 214010 157176
rect 214066 157120 217212 157176
rect 214005 157118 217212 157120
rect 214005 157115 214071 157118
rect 306741 157042 306807 157045
rect 324313 157042 324379 157045
rect 306741 157040 310132 157042
rect 306741 156984 306746 157040
rect 306802 156984 310132 157040
rect 306741 156982 310132 156984
rect 321908 157040 324379 157042
rect 321908 156984 324318 157040
rect 324374 156984 324379 157040
rect 321908 156982 324379 156984
rect 306741 156979 306807 156982
rect 324313 156979 324379 156982
rect 252369 156906 252435 156909
rect 248860 156904 252435 156906
rect 248860 156848 252374 156904
rect 252430 156848 252435 156904
rect 248860 156846 252435 156848
rect 252369 156843 252435 156846
rect 307569 156634 307635 156637
rect 307569 156632 310132 156634
rect 307569 156576 307574 156632
rect 307630 156576 310132 156632
rect 307569 156574 310132 156576
rect 307569 156571 307635 156574
rect 213913 156498 213979 156501
rect 213913 156496 217212 156498
rect 213913 156440 213918 156496
rect 213974 156440 217212 156496
rect 213913 156438 217212 156440
rect 213913 156435 213979 156438
rect 259494 156362 259500 156364
rect 248860 156302 259500 156362
rect 259494 156300 259500 156302
rect 259564 156300 259570 156364
rect 324405 156362 324471 156365
rect 321908 156360 324471 156362
rect 321908 156304 324410 156360
rect 324466 156304 324471 156360
rect 321908 156302 324471 156304
rect 324405 156299 324471 156302
rect 307661 156226 307727 156229
rect 307661 156224 310132 156226
rect 307661 156168 307666 156224
rect 307722 156168 310132 156224
rect 307661 156166 310132 156168
rect 307661 156163 307727 156166
rect 252461 155954 252527 155957
rect 248860 155952 252527 155954
rect 248860 155896 252466 155952
rect 252522 155896 252527 155952
rect 248860 155894 252527 155896
rect 252461 155891 252527 155894
rect 213913 155818 213979 155821
rect 213913 155816 217212 155818
rect 213913 155760 213918 155816
rect 213974 155760 217212 155816
rect 213913 155758 217212 155760
rect 213913 155755 213979 155758
rect 307477 155682 307543 155685
rect 307477 155680 310132 155682
rect 307477 155624 307482 155680
rect 307538 155624 310132 155680
rect 307477 155622 310132 155624
rect 307477 155619 307543 155622
rect 324313 155546 324379 155549
rect 321908 155544 324379 155546
rect 321908 155488 324318 155544
rect 324374 155488 324379 155544
rect 321908 155486 324379 155488
rect 324313 155483 324379 155486
rect 249793 155410 249859 155413
rect 248860 155408 249859 155410
rect 248860 155352 249798 155408
rect 249854 155352 249859 155408
rect 248860 155350 249859 155352
rect 249793 155347 249859 155350
rect 251950 155212 251956 155276
rect 252020 155274 252026 155276
rect 282177 155274 282243 155277
rect 252020 155272 282243 155274
rect 252020 155216 282182 155272
rect 282238 155216 282243 155272
rect 252020 155214 282243 155216
rect 252020 155212 252026 155214
rect 282177 155211 282243 155214
rect 307569 155274 307635 155277
rect 307569 155272 310132 155274
rect 307569 155216 307574 155272
rect 307630 155216 310132 155272
rect 307569 155214 310132 155216
rect 307569 155211 307635 155214
rect 167494 154532 167500 154596
rect 167564 154594 167570 154596
rect 217182 154594 217242 155108
rect 252369 155002 252435 155005
rect 248860 155000 252435 155002
rect 248860 154944 252374 155000
rect 252430 154944 252435 155000
rect 248860 154942 252435 154944
rect 252369 154939 252435 154942
rect 307661 154866 307727 154869
rect 307661 154864 310132 154866
rect 307661 154808 307666 154864
rect 307722 154808 310132 154864
rect 307661 154806 310132 154808
rect 307661 154803 307727 154806
rect 324497 154730 324563 154733
rect 321908 154728 324563 154730
rect 321908 154672 324502 154728
rect 324558 154672 324563 154728
rect 321908 154670 324563 154672
rect 324497 154667 324563 154670
rect 167564 154534 217242 154594
rect 167564 154532 167570 154534
rect 213913 154458 213979 154461
rect 252553 154458 252619 154461
rect 213913 154456 217212 154458
rect 213913 154400 213918 154456
rect 213974 154400 217212 154456
rect 213913 154398 217212 154400
rect 248860 154456 252619 154458
rect 248860 154400 252558 154456
rect 252614 154400 252619 154456
rect 248860 154398 252619 154400
rect 213913 154395 213979 154398
rect 252553 154395 252619 154398
rect 307201 154458 307267 154461
rect 307201 154456 310132 154458
rect 307201 154400 307206 154456
rect 307262 154400 310132 154456
rect 307201 154398 310132 154400
rect 307201 154395 307267 154398
rect 252461 154050 252527 154053
rect 248860 154048 252527 154050
rect 248860 153992 252466 154048
rect 252522 153992 252527 154048
rect 248860 153990 252527 153992
rect 252461 153987 252527 153990
rect 307477 154050 307543 154053
rect 324313 154050 324379 154053
rect 307477 154048 310132 154050
rect 307477 153992 307482 154048
rect 307538 153992 310132 154048
rect 307477 153990 310132 153992
rect 321908 154048 324379 154050
rect 321908 153992 324318 154048
rect 324374 153992 324379 154048
rect 321908 153990 324379 153992
rect 307477 153987 307543 153990
rect 324313 153987 324379 153990
rect 215937 153778 216003 153781
rect 215937 153776 217212 153778
rect 215937 153720 215942 153776
rect 215998 153720 217212 153776
rect 215937 153718 217212 153720
rect 215937 153715 216003 153718
rect 307661 153642 307727 153645
rect 307661 153640 310132 153642
rect 307661 153584 307666 153640
rect 307722 153584 310132 153640
rect 307661 153582 310132 153584
rect 307661 153579 307727 153582
rect 252369 153506 252435 153509
rect 248860 153504 252435 153506
rect 248860 153448 252374 153504
rect 252430 153448 252435 153504
rect 248860 153446 252435 153448
rect 252369 153443 252435 153446
rect 306649 153234 306715 153237
rect 322933 153234 322999 153237
rect 306649 153232 310132 153234
rect 306649 153176 306654 153232
rect 306710 153176 310132 153232
rect 306649 153174 310132 153176
rect 321908 153232 322999 153234
rect 321908 153176 322938 153232
rect 322994 153176 322999 153232
rect 321908 153174 322999 153176
rect 306649 153171 306715 153174
rect 322933 153171 322999 153174
rect 214005 153098 214071 153101
rect 252461 153098 252527 153101
rect 214005 153096 217212 153098
rect 214005 153040 214010 153096
rect 214066 153040 217212 153096
rect 214005 153038 217212 153040
rect 248860 153096 252527 153098
rect 248860 153040 252466 153096
rect 252522 153040 252527 153096
rect 248860 153038 252527 153040
rect 214005 153035 214071 153038
rect 252461 153035 252527 153038
rect 250437 152962 250503 152965
rect 257838 152962 257844 152964
rect 250437 152960 257844 152962
rect 250437 152904 250442 152960
rect 250498 152904 257844 152960
rect 250437 152902 257844 152904
rect 250437 152899 250503 152902
rect 257838 152900 257844 152902
rect 257908 152900 257914 152964
rect 252502 152690 252508 152692
rect 248860 152630 252508 152690
rect 252502 152628 252508 152630
rect 252572 152628 252578 152692
rect 307477 152690 307543 152693
rect 580257 152690 580323 152693
rect 583520 152690 584960 152780
rect 307477 152688 310132 152690
rect 307477 152632 307482 152688
rect 307538 152632 310132 152688
rect 307477 152630 310132 152632
rect 580257 152688 584960 152690
rect 580257 152632 580262 152688
rect 580318 152632 584960 152688
rect 580257 152630 584960 152632
rect 307477 152627 307543 152630
rect 580257 152627 580323 152630
rect 213913 152554 213979 152557
rect 213913 152552 217212 152554
rect 213913 152496 213918 152552
rect 213974 152496 217212 152552
rect 583520 152540 584960 152630
rect 213913 152494 217212 152496
rect 213913 152491 213979 152494
rect 324313 152418 324379 152421
rect 321908 152416 324379 152418
rect 321908 152360 324318 152416
rect 324374 152360 324379 152416
rect 321908 152358 324379 152360
rect 324313 152355 324379 152358
rect 307661 152282 307727 152285
rect 307661 152280 310132 152282
rect 307661 152224 307666 152280
rect 307722 152224 310132 152280
rect 307661 152222 310132 152224
rect 307661 152219 307727 152222
rect 251173 152146 251239 152149
rect 248860 152144 251239 152146
rect 248860 152088 251178 152144
rect 251234 152088 251239 152144
rect 248860 152086 251239 152088
rect 251173 152083 251239 152086
rect 213269 151874 213335 151877
rect 307661 151874 307727 151877
rect 213269 151872 217212 151874
rect 213269 151816 213274 151872
rect 213330 151816 217212 151872
rect 213269 151814 217212 151816
rect 307661 151872 310132 151874
rect 307661 151816 307666 151872
rect 307722 151816 310132 151872
rect 307661 151814 310132 151816
rect 213269 151811 213335 151814
rect 307661 151811 307727 151814
rect 252461 151738 252527 151741
rect 324313 151738 324379 151741
rect 248860 151736 252527 151738
rect 248860 151680 252466 151736
rect 252522 151680 252527 151736
rect 248860 151678 252527 151680
rect 321908 151736 324379 151738
rect 321908 151680 324318 151736
rect 324374 151680 324379 151736
rect 321908 151678 324379 151680
rect 252461 151675 252527 151678
rect 324313 151675 324379 151678
rect 307477 151466 307543 151469
rect 307477 151464 310132 151466
rect 307477 151408 307482 151464
rect 307538 151408 310132 151464
rect 307477 151406 310132 151408
rect 307477 151403 307543 151406
rect 321737 151330 321803 151333
rect 321694 151328 321803 151330
rect 321694 151272 321742 151328
rect 321798 151272 321803 151328
rect 321694 151267 321803 151272
rect 214005 151194 214071 151197
rect 251265 151194 251331 151197
rect 214005 151192 217212 151194
rect 214005 151136 214010 151192
rect 214066 151136 217212 151192
rect 214005 151134 217212 151136
rect 248860 151192 251331 151194
rect 248860 151136 251270 151192
rect 251326 151136 251331 151192
rect 248860 151134 251331 151136
rect 214005 151131 214071 151134
rect 251265 151131 251331 151134
rect 307661 151058 307727 151061
rect 307661 151056 310132 151058
rect 307661 151000 307666 151056
rect 307722 151000 310132 151056
rect 307661 150998 310132 151000
rect 307661 150995 307727 150998
rect 321694 150892 321754 151267
rect 249977 150786 250043 150789
rect 248860 150784 250043 150786
rect 248860 150728 249982 150784
rect 250038 150728 250043 150784
rect 248860 150726 250043 150728
rect 249977 150723 250043 150726
rect 306925 150650 306991 150653
rect 306925 150648 310132 150650
rect 306925 150592 306930 150648
rect 306986 150592 310132 150648
rect 306925 150590 310132 150592
rect 306925 150587 306991 150590
rect 214649 150514 214715 150517
rect 214649 150512 217212 150514
rect 214649 150456 214654 150512
rect 214710 150456 217212 150512
rect 214649 150454 217212 150456
rect 214649 150451 214715 150454
rect 256918 150242 256924 150244
rect 248860 150182 256924 150242
rect 256918 150180 256924 150182
rect 256988 150180 256994 150244
rect 306925 150242 306991 150245
rect 306925 150240 310132 150242
rect 306925 150184 306930 150240
rect 306986 150184 310132 150240
rect 306925 150182 310132 150184
rect 306925 150179 306991 150182
rect 324313 150106 324379 150109
rect 321908 150104 324379 150106
rect 321908 150048 324318 150104
rect 324374 150048 324379 150104
rect 321908 150046 324379 150048
rect 324313 150043 324379 150046
rect 213913 149834 213979 149837
rect 252277 149834 252343 149837
rect 213913 149832 217212 149834
rect 213913 149776 213918 149832
rect 213974 149776 217212 149832
rect 213913 149774 217212 149776
rect 248860 149832 252343 149834
rect 248860 149776 252282 149832
rect 252338 149776 252343 149832
rect 248860 149774 252343 149776
rect 213913 149771 213979 149774
rect 252277 149771 252343 149774
rect 307661 149834 307727 149837
rect 307661 149832 310132 149834
rect 307661 149776 307666 149832
rect 307722 149776 310132 149832
rect 307661 149774 310132 149776
rect 307661 149771 307727 149774
rect 324405 149426 324471 149429
rect 321908 149424 324471 149426
rect 321908 149368 324410 149424
rect 324466 149368 324471 149424
rect 321908 149366 324471 149368
rect 324405 149363 324471 149366
rect 251725 149290 251791 149293
rect 248860 149288 251791 149290
rect 248860 149232 251730 149288
rect 251786 149232 251791 149288
rect 248860 149230 251791 149232
rect 251725 149227 251791 149230
rect 307569 149290 307635 149293
rect 307569 149288 310132 149290
rect 307569 149232 307574 149288
rect 307630 149232 310132 149288
rect 307569 149230 310132 149232
rect 307569 149227 307635 149230
rect 214005 149154 214071 149157
rect 214005 149152 217212 149154
rect 214005 149096 214010 149152
rect 214066 149096 217212 149152
rect 214005 149094 217212 149096
rect 214005 149091 214071 149094
rect 251265 148882 251331 148885
rect 248860 148880 251331 148882
rect 248860 148824 251270 148880
rect 251326 148824 251331 148880
rect 248860 148822 251331 148824
rect 251265 148819 251331 148822
rect 306925 148882 306991 148885
rect 306925 148880 310132 148882
rect 306925 148824 306930 148880
rect 306986 148824 310132 148880
rect 306925 148822 310132 148824
rect 306925 148819 306991 148822
rect 324313 148610 324379 148613
rect 321908 148608 324379 148610
rect 321908 148552 324318 148608
rect 324374 148552 324379 148608
rect 321908 148550 324379 148552
rect 324313 148547 324379 148550
rect 214557 148474 214623 148477
rect 307017 148474 307083 148477
rect 214557 148472 217212 148474
rect 214557 148416 214562 148472
rect 214618 148416 217212 148472
rect 214557 148414 217212 148416
rect 307017 148472 310132 148474
rect 307017 148416 307022 148472
rect 307078 148416 310132 148472
rect 307017 148414 310132 148416
rect 214557 148411 214623 148414
rect 307017 148411 307083 148414
rect 251909 148338 251975 148341
rect 248860 148336 251975 148338
rect 248860 148280 251914 148336
rect 251970 148280 251975 148336
rect 248860 148278 251975 148280
rect 251909 148275 251975 148278
rect 307661 148066 307727 148069
rect 307661 148064 310132 148066
rect 307661 148008 307666 148064
rect 307722 148008 310132 148064
rect 307661 148006 310132 148008
rect 307661 148003 307727 148006
rect 213913 147930 213979 147933
rect 252461 147930 252527 147933
rect 213913 147928 217212 147930
rect 213913 147872 213918 147928
rect 213974 147872 217212 147928
rect 213913 147870 217212 147872
rect 248860 147928 252527 147930
rect 248860 147872 252466 147928
rect 252522 147872 252527 147928
rect 248860 147870 252527 147872
rect 213913 147867 213979 147870
rect 252461 147867 252527 147870
rect 324405 147794 324471 147797
rect 321908 147792 324471 147794
rect 321908 147736 324410 147792
rect 324466 147736 324471 147792
rect 321908 147734 324471 147736
rect 324405 147731 324471 147734
rect 307385 147658 307451 147661
rect 307385 147656 310132 147658
rect 307385 147600 307390 147656
rect 307446 147600 310132 147656
rect 307385 147598 310132 147600
rect 307385 147595 307451 147598
rect 252461 147522 252527 147525
rect 248860 147520 252527 147522
rect 248860 147464 252466 147520
rect 252522 147464 252527 147520
rect 248860 147462 252527 147464
rect 252461 147459 252527 147462
rect 214005 147250 214071 147253
rect 306741 147250 306807 147253
rect 214005 147248 217212 147250
rect 214005 147192 214010 147248
rect 214066 147192 217212 147248
rect 214005 147190 217212 147192
rect 306741 147248 310132 147250
rect 306741 147192 306746 147248
rect 306802 147192 310132 147248
rect 306741 147190 310132 147192
rect 214005 147187 214071 147190
rect 306741 147187 306807 147190
rect 324313 147114 324379 147117
rect 321908 147112 324379 147114
rect 321908 147056 324318 147112
rect 324374 147056 324379 147112
rect 321908 147054 324379 147056
rect 324313 147051 324379 147054
rect 251725 146978 251791 146981
rect 248860 146976 251791 146978
rect 248860 146920 251730 146976
rect 251786 146920 251791 146976
rect 248860 146918 251791 146920
rect 251725 146915 251791 146918
rect 307661 146842 307727 146845
rect 307661 146840 310132 146842
rect 307661 146784 307666 146840
rect 307722 146784 310132 146840
rect 307661 146782 310132 146784
rect 307661 146779 307727 146782
rect 213913 146570 213979 146573
rect 251725 146570 251791 146573
rect 213913 146568 217212 146570
rect 213913 146512 213918 146568
rect 213974 146512 217212 146568
rect 213913 146510 217212 146512
rect 248860 146568 251791 146570
rect 248860 146512 251730 146568
rect 251786 146512 251791 146568
rect 248860 146510 251791 146512
rect 213913 146507 213979 146510
rect 251725 146507 251791 146510
rect 305821 146434 305887 146437
rect 305821 146432 310132 146434
rect 305821 146376 305826 146432
rect 305882 146376 310132 146432
rect 305821 146374 310132 146376
rect 305821 146371 305887 146374
rect 324313 146298 324379 146301
rect 321908 146296 324379 146298
rect 321908 146240 324318 146296
rect 324374 146240 324379 146296
rect 321908 146238 324379 146240
rect 324313 146235 324379 146238
rect 251909 146026 251975 146029
rect 248860 146024 251975 146026
rect 248860 145968 251914 146024
rect 251970 145968 251975 146024
rect 248860 145966 251975 145968
rect 251909 145963 251975 145966
rect 214005 145890 214071 145893
rect 307477 145890 307543 145893
rect 214005 145888 217212 145890
rect 214005 145832 214010 145888
rect 214066 145832 217212 145888
rect 214005 145830 217212 145832
rect 307477 145888 310132 145890
rect 307477 145832 307482 145888
rect 307538 145832 310132 145888
rect 307477 145830 310132 145832
rect 214005 145827 214071 145830
rect 307477 145827 307543 145830
rect 251725 145618 251791 145621
rect 248860 145616 251791 145618
rect 248860 145560 251730 145616
rect 251786 145560 251791 145616
rect 248860 145558 251791 145560
rect 251725 145555 251791 145558
rect 307569 145482 307635 145485
rect 324405 145482 324471 145485
rect 307569 145480 310132 145482
rect 307569 145424 307574 145480
rect 307630 145424 310132 145480
rect 307569 145422 310132 145424
rect 321908 145480 324471 145482
rect 321908 145424 324410 145480
rect 324466 145424 324471 145480
rect 321908 145422 324471 145424
rect 307569 145419 307635 145422
rect 324405 145419 324471 145422
rect 213913 145210 213979 145213
rect 213913 145208 217212 145210
rect 213913 145152 213918 145208
rect 213974 145152 217212 145208
rect 213913 145150 217212 145152
rect 213913 145147 213979 145150
rect 252093 145074 252159 145077
rect 248860 145072 252159 145074
rect 248860 145016 252098 145072
rect 252154 145016 252159 145072
rect 248860 145014 252159 145016
rect 252093 145011 252159 145014
rect 307661 145074 307727 145077
rect 307661 145072 310132 145074
rect 307661 145016 307666 145072
rect 307722 145016 310132 145072
rect 307661 145014 310132 145016
rect 307661 145011 307727 145014
rect 324313 144802 324379 144805
rect 321908 144800 324379 144802
rect 321908 144744 324318 144800
rect 324374 144744 324379 144800
rect 321908 144742 324379 144744
rect 324313 144739 324379 144742
rect 252461 144666 252527 144669
rect 248860 144664 252527 144666
rect 248860 144608 252466 144664
rect 252522 144608 252527 144664
rect 248860 144606 252527 144608
rect 252461 144603 252527 144606
rect 306557 144666 306623 144669
rect 306557 144664 310132 144666
rect 306557 144608 306562 144664
rect 306618 144608 310132 144664
rect 306557 144606 310132 144608
rect 306557 144603 306623 144606
rect 214005 144530 214071 144533
rect 214005 144528 217212 144530
rect 214005 144472 214010 144528
rect 214066 144472 217212 144528
rect 214005 144470 217212 144472
rect 214005 144467 214071 144470
rect 307661 144258 307727 144261
rect 307661 144256 310132 144258
rect 307661 144200 307666 144256
rect 307722 144200 310132 144256
rect 307661 144198 310132 144200
rect 307661 144195 307727 144198
rect 252369 144122 252435 144125
rect 248860 144120 252435 144122
rect 248860 144064 252374 144120
rect 252430 144064 252435 144120
rect 248860 144062 252435 144064
rect 252369 144059 252435 144062
rect 255957 144122 256023 144125
rect 306966 144122 306972 144124
rect 255957 144120 306972 144122
rect 255957 144064 255962 144120
rect 256018 144064 306972 144120
rect 255957 144062 306972 144064
rect 255957 144059 256023 144062
rect 306966 144060 306972 144062
rect 307036 144060 307042 144124
rect 324405 143986 324471 143989
rect 321908 143984 324471 143986
rect 321908 143928 324410 143984
rect 324466 143928 324471 143984
rect 321908 143926 324471 143928
rect 324405 143923 324471 143926
rect 213913 143850 213979 143853
rect 213913 143848 217212 143850
rect 213913 143792 213918 143848
rect 213974 143792 217212 143848
rect 213913 143790 217212 143792
rect 213913 143787 213979 143790
rect 307702 143788 307708 143852
rect 307772 143850 307778 143852
rect 307772 143790 310132 143850
rect 307772 143788 307778 143790
rect 252461 143714 252527 143717
rect 248860 143712 252527 143714
rect 248860 143656 252466 143712
rect 252522 143656 252527 143712
rect 248860 143654 252527 143656
rect 252461 143651 252527 143654
rect 307661 143442 307727 143445
rect 307661 143440 310132 143442
rect 307661 143384 307666 143440
rect 307722 143384 310132 143440
rect 307661 143382 310132 143384
rect 307661 143379 307727 143382
rect 214005 143306 214071 143309
rect 214005 143304 217212 143306
rect 214005 143248 214010 143304
rect 214066 143248 217212 143304
rect 214005 143246 217212 143248
rect 214005 143243 214071 143246
rect 252461 143170 252527 143173
rect 248860 143168 252527 143170
rect 248860 143112 252466 143168
rect 252522 143112 252527 143168
rect 248860 143110 252527 143112
rect 252461 143107 252527 143110
rect 306741 143034 306807 143037
rect 306741 143032 310132 143034
rect 306741 142976 306746 143032
rect 306802 142976 310132 143032
rect 306741 142974 310132 142976
rect 306741 142971 306807 142974
rect 253381 142762 253447 142765
rect 248860 142760 253447 142762
rect 248860 142704 253386 142760
rect 253442 142704 253447 142760
rect 248860 142702 253447 142704
rect 253381 142699 253447 142702
rect 293493 142762 293559 142765
rect 307702 142762 307708 142764
rect 293493 142760 307708 142762
rect 293493 142704 293498 142760
rect 293554 142704 307708 142760
rect 293493 142702 307708 142704
rect 293493 142699 293559 142702
rect 307702 142700 307708 142702
rect 307772 142700 307778 142764
rect 213913 142626 213979 142629
rect 321878 142626 321938 143140
rect 324681 142762 324747 142765
rect 331438 142762 331444 142764
rect 324681 142760 331444 142762
rect 324681 142704 324686 142760
rect 324742 142704 331444 142760
rect 324681 142702 331444 142704
rect 324681 142699 324747 142702
rect 331438 142700 331444 142702
rect 331508 142700 331514 142764
rect 213913 142624 217212 142626
rect 213913 142568 213918 142624
rect 213974 142568 217212 142624
rect 213913 142566 217212 142568
rect 321878 142566 325710 142626
rect 213913 142563 213979 142566
rect 265014 142490 265020 142492
rect 253246 142430 265020 142490
rect 253246 142218 253306 142430
rect 265014 142428 265020 142430
rect 265084 142428 265090 142492
rect 306414 142428 306420 142492
rect 306484 142490 306490 142492
rect 324313 142490 324379 142493
rect 306484 142430 310132 142490
rect 321908 142488 324379 142490
rect 321908 142432 324318 142488
rect 324374 142432 324379 142488
rect 321908 142430 324379 142432
rect 306484 142428 306490 142430
rect 324313 142427 324379 142430
rect 253381 142354 253447 142357
rect 260966 142354 260972 142356
rect 253381 142352 260972 142354
rect 253381 142296 253386 142352
rect 253442 142296 260972 142352
rect 253381 142294 260972 142296
rect 253381 142291 253447 142294
rect 260966 142292 260972 142294
rect 261036 142292 261042 142356
rect 248860 142158 253306 142218
rect 325650 142218 325710 142566
rect 335670 142218 335676 142220
rect 325650 142158 335676 142218
rect 335670 142156 335676 142158
rect 335740 142156 335746 142220
rect 307293 142082 307359 142085
rect 307293 142080 310132 142082
rect 307293 142024 307298 142080
rect 307354 142024 310132 142080
rect 307293 142022 310132 142024
rect 307293 142019 307359 142022
rect 213913 141946 213979 141949
rect 213913 141944 217212 141946
rect 213913 141888 213918 141944
rect 213974 141888 217212 141944
rect 213913 141886 217212 141888
rect 213913 141883 213979 141886
rect 262254 141810 262260 141812
rect 248860 141750 262260 141810
rect 262254 141748 262260 141750
rect 262324 141748 262330 141812
rect 307385 141674 307451 141677
rect 324313 141674 324379 141677
rect 307385 141672 310132 141674
rect 307385 141616 307390 141672
rect 307446 141616 310132 141672
rect 307385 141614 310132 141616
rect 321908 141672 324379 141674
rect 321908 141616 324318 141672
rect 324374 141616 324379 141672
rect 321908 141614 324379 141616
rect 307385 141611 307451 141614
rect 324313 141611 324379 141614
rect 252461 141402 252527 141405
rect 248860 141400 252527 141402
rect 248860 141344 252466 141400
rect 252522 141344 252527 141400
rect 248860 141342 252527 141344
rect 252461 141339 252527 141342
rect 292113 141402 292179 141405
rect 306414 141402 306420 141404
rect 292113 141400 306420 141402
rect 292113 141344 292118 141400
rect 292174 141344 306420 141400
rect 292113 141342 306420 141344
rect 292113 141339 292179 141342
rect 306414 141340 306420 141342
rect 306484 141340 306490 141404
rect 307661 141266 307727 141269
rect 307661 141264 310132 141266
rect 167494 140796 167500 140860
rect 167564 140858 167570 140860
rect 217182 140858 217242 141236
rect 307661 141208 307666 141264
rect 307722 141208 310132 141264
rect 307661 141206 310132 141208
rect 307661 141203 307727 141206
rect 251265 140858 251331 140861
rect 167564 140798 217242 140858
rect 248860 140856 251331 140858
rect 248860 140800 251270 140856
rect 251326 140800 251331 140856
rect 248860 140798 251331 140800
rect 167564 140796 167570 140798
rect 251265 140795 251331 140798
rect 307702 140796 307708 140860
rect 307772 140858 307778 140860
rect 324497 140858 324563 140861
rect 307772 140798 310132 140858
rect 321908 140856 324563 140858
rect 321908 140800 324502 140856
rect 324558 140800 324563 140856
rect 321908 140798 324563 140800
rect 307772 140796 307778 140798
rect 324497 140795 324563 140798
rect 213913 140586 213979 140589
rect 213913 140584 217212 140586
rect 213913 140528 213918 140584
rect 213974 140528 217212 140584
rect 213913 140526 217212 140528
rect 213913 140523 213979 140526
rect 255262 140450 255268 140452
rect 248860 140390 255268 140450
rect 255262 140388 255268 140390
rect 255332 140388 255338 140452
rect 307201 140450 307267 140453
rect 307201 140448 310132 140450
rect 307201 140392 307206 140448
rect 307262 140392 310132 140448
rect 307201 140390 310132 140392
rect 307201 140387 307267 140390
rect 324681 140178 324747 140181
rect 321908 140176 324747 140178
rect 321908 140120 324686 140176
rect 324742 140120 324747 140176
rect 321908 140118 324747 140120
rect 324681 140115 324747 140118
rect 307569 140042 307635 140045
rect 307569 140040 310132 140042
rect 307569 139984 307574 140040
rect 307630 139984 310132 140040
rect 307569 139982 310132 139984
rect 307569 139979 307635 139982
rect 251357 139906 251423 139909
rect 248860 139904 251423 139906
rect 166206 139436 166212 139500
rect 166276 139498 166282 139500
rect 217182 139498 217242 139876
rect 248860 139848 251362 139904
rect 251418 139848 251423 139904
rect 248860 139846 251423 139848
rect 251357 139843 251423 139846
rect 307661 139634 307727 139637
rect 307661 139632 310132 139634
rect 307661 139576 307666 139632
rect 307722 139576 310132 139632
rect 307661 139574 310132 139576
rect 307661 139571 307727 139574
rect 249190 139498 249196 139500
rect 166276 139438 217242 139498
rect 248860 139438 249196 139498
rect 166276 139436 166282 139438
rect 249190 139436 249196 139438
rect 249260 139436 249266 139500
rect 324313 139362 324379 139365
rect 583520 139362 584960 139452
rect 321908 139360 324379 139362
rect 321908 139304 324318 139360
rect 324374 139304 324379 139360
rect 321908 139302 324379 139304
rect 324313 139299 324379 139302
rect 583342 139302 584960 139362
rect 214649 139226 214715 139229
rect 583342 139226 583402 139302
rect 583520 139226 584960 139302
rect 214649 139224 217212 139226
rect 214649 139168 214654 139224
rect 214710 139168 217212 139224
rect 214649 139166 217212 139168
rect 583342 139212 584960 139226
rect 583342 139166 583586 139212
rect 214649 139163 214715 139166
rect 307477 139090 307543 139093
rect 307477 139088 310132 139090
rect 307477 139032 307482 139088
rect 307538 139032 310132 139088
rect 307477 139030 310132 139032
rect 307477 139027 307543 139030
rect 249885 138954 249951 138957
rect 248860 138952 249951 138954
rect 248860 138896 249890 138952
rect 249946 138896 249951 138952
rect 248860 138894 249951 138896
rect 249885 138891 249951 138894
rect 213913 138682 213979 138685
rect 213913 138680 217212 138682
rect 213913 138624 213918 138680
rect 213974 138624 217212 138680
rect 213913 138622 217212 138624
rect 213913 138619 213979 138622
rect 251766 138620 251772 138684
rect 251836 138682 251842 138684
rect 274081 138682 274147 138685
rect 251836 138680 274147 138682
rect 251836 138624 274086 138680
rect 274142 138624 274147 138680
rect 251836 138622 274147 138624
rect 251836 138620 251842 138622
rect 274081 138619 274147 138622
rect 307569 138682 307635 138685
rect 307569 138680 310132 138682
rect 307569 138624 307574 138680
rect 307630 138624 310132 138680
rect 307569 138622 310132 138624
rect 307569 138619 307635 138622
rect 252461 138546 252527 138549
rect 324497 138546 324563 138549
rect 248860 138544 252527 138546
rect 248860 138488 252466 138544
rect 252522 138488 252527 138544
rect 248860 138486 252527 138488
rect 321908 138544 324563 138546
rect 321908 138488 324502 138544
rect 324558 138488 324563 138544
rect 321908 138486 324563 138488
rect 252461 138483 252527 138486
rect 324497 138483 324563 138486
rect 307661 138274 307727 138277
rect 307661 138272 310132 138274
rect 307661 138216 307666 138272
rect 307722 138216 310132 138272
rect 307661 138214 310132 138216
rect 307661 138211 307727 138214
rect 249885 138138 249951 138141
rect 263542 138138 263548 138140
rect 249885 138136 263548 138138
rect 249885 138080 249890 138136
rect 249946 138080 263548 138136
rect 249885 138078 263548 138080
rect 249885 138075 249951 138078
rect 263542 138076 263548 138078
rect 263612 138076 263618 138140
rect 346158 138076 346164 138140
rect 346228 138138 346234 138140
rect 583526 138138 583586 139166
rect 346228 138078 583586 138138
rect 346228 138076 346234 138078
rect 214097 138002 214163 138005
rect 251357 138002 251423 138005
rect 214097 138000 217212 138002
rect 214097 137944 214102 138000
rect 214158 137944 217212 138000
rect 214097 137942 217212 137944
rect 248860 138000 251423 138002
rect 248860 137944 251362 138000
rect 251418 137944 251423 138000
rect 248860 137942 251423 137944
rect 214097 137939 214163 137942
rect 251357 137939 251423 137942
rect 306925 137866 306991 137869
rect 324313 137866 324379 137869
rect 306925 137864 310132 137866
rect 306925 137808 306930 137864
rect 306986 137808 310132 137864
rect 306925 137806 310132 137808
rect 321908 137864 324379 137866
rect 321908 137808 324318 137864
rect 324374 137808 324379 137864
rect 321908 137806 324379 137808
rect 306925 137803 306991 137806
rect 324313 137803 324379 137806
rect 256734 137594 256740 137596
rect 248860 137534 256740 137594
rect 256734 137532 256740 137534
rect 256804 137532 256810 137596
rect 307477 137458 307543 137461
rect 307477 137456 310132 137458
rect 307477 137400 307482 137456
rect 307538 137400 310132 137456
rect 307477 137398 310132 137400
rect 307477 137395 307543 137398
rect 213913 137322 213979 137325
rect 213913 137320 217212 137322
rect 213913 137264 213918 137320
rect 213974 137264 217212 137320
rect 213913 137262 217212 137264
rect 213913 137259 213979 137262
rect 252461 137050 252527 137053
rect 248860 137048 252527 137050
rect 248860 136992 252466 137048
rect 252522 136992 252527 137048
rect 248860 136990 252527 136992
rect 252461 136987 252527 136990
rect 307109 137050 307175 137053
rect 324497 137050 324563 137053
rect 307109 137048 310132 137050
rect 307109 136992 307114 137048
rect 307170 136992 310132 137048
rect 307109 136990 310132 136992
rect 321908 137048 324563 137050
rect 321908 136992 324502 137048
rect 324558 136992 324563 137048
rect 321908 136990 324563 136992
rect 307109 136987 307175 136990
rect 324497 136987 324563 136990
rect 214005 136642 214071 136645
rect 250437 136642 250503 136645
rect 214005 136640 217212 136642
rect 214005 136584 214010 136640
rect 214066 136584 217212 136640
rect 214005 136582 217212 136584
rect 248860 136640 250503 136642
rect 248860 136584 250442 136640
rect 250498 136584 250503 136640
rect 248860 136582 250503 136584
rect 214005 136579 214071 136582
rect 250437 136579 250503 136582
rect 307385 136642 307451 136645
rect 307385 136640 310132 136642
rect 307385 136584 307390 136640
rect 307446 136584 310132 136640
rect 307385 136582 310132 136584
rect 307385 136579 307451 136582
rect 324313 136370 324379 136373
rect 321908 136368 324379 136370
rect 321908 136312 324318 136368
rect 324374 136312 324379 136368
rect 321908 136310 324379 136312
rect 324313 136307 324379 136310
rect 251541 136234 251607 136237
rect 248860 136232 251607 136234
rect 248860 136176 251546 136232
rect 251602 136176 251607 136232
rect 248860 136174 251607 136176
rect 251541 136171 251607 136174
rect 307661 136234 307727 136237
rect 307661 136232 310132 136234
rect 307661 136176 307666 136232
rect 307722 136176 310132 136232
rect 307661 136174 310132 136176
rect 307661 136171 307727 136174
rect 170438 135492 170444 135556
rect 170508 135554 170514 135556
rect 217182 135554 217242 135932
rect 252461 135690 252527 135693
rect 248860 135688 252527 135690
rect 248860 135632 252466 135688
rect 252522 135632 252527 135688
rect 248860 135630 252527 135632
rect 252461 135627 252527 135630
rect 307477 135690 307543 135693
rect 307477 135688 310132 135690
rect 307477 135632 307482 135688
rect 307538 135632 310132 135688
rect 307477 135630 310132 135632
rect 307477 135627 307543 135630
rect 324497 135554 324563 135557
rect 170508 135494 217242 135554
rect 321908 135552 324563 135554
rect 321908 135496 324502 135552
rect 324558 135496 324563 135552
rect 321908 135494 324563 135496
rect 170508 135492 170514 135494
rect 324497 135491 324563 135494
rect 213913 135282 213979 135285
rect 252369 135282 252435 135285
rect 213913 135280 217212 135282
rect 213913 135224 213918 135280
rect 213974 135224 217212 135280
rect 213913 135222 217212 135224
rect 248860 135280 252435 135282
rect 248860 135224 252374 135280
rect 252430 135224 252435 135280
rect 248860 135222 252435 135224
rect 213913 135219 213979 135222
rect 252369 135219 252435 135222
rect 307569 135282 307635 135285
rect 307569 135280 310132 135282
rect 307569 135224 307574 135280
rect 307630 135224 310132 135280
rect 307569 135222 310132 135224
rect 307569 135219 307635 135222
rect 306741 134874 306807 134877
rect 306741 134872 310132 134874
rect 306741 134816 306746 134872
rect 306802 134816 310132 134872
rect 306741 134814 310132 134816
rect 306741 134811 306807 134814
rect 251633 134738 251699 134741
rect 248860 134736 251699 134738
rect 248860 134680 251638 134736
rect 251694 134680 251699 134736
rect 248860 134678 251699 134680
rect 251633 134675 251699 134678
rect 214005 134602 214071 134605
rect 214005 134600 217212 134602
rect 214005 134544 214010 134600
rect 214066 134544 217212 134600
rect 214005 134542 217212 134544
rect 214005 134539 214071 134542
rect 307569 134466 307635 134469
rect 307569 134464 310132 134466
rect 307569 134408 307574 134464
rect 307630 134408 310132 134464
rect 307569 134406 310132 134408
rect 307569 134403 307635 134406
rect 252461 134330 252527 134333
rect 248860 134328 252527 134330
rect 248860 134272 252466 134328
rect 252522 134272 252527 134328
rect 248860 134270 252527 134272
rect 252461 134267 252527 134270
rect 321878 134194 321938 134708
rect 340822 134194 340828 134196
rect 321878 134134 340828 134194
rect 340822 134132 340828 134134
rect 340892 134132 340898 134196
rect 307661 134058 307727 134061
rect 325785 134058 325851 134061
rect 307661 134056 310132 134058
rect 307661 134000 307666 134056
rect 307722 134000 310132 134056
rect 307661 133998 310132 134000
rect 321908 134056 325851 134058
rect 321908 134000 325790 134056
rect 325846 134000 325851 134056
rect 321908 133998 325851 134000
rect 307661 133995 307727 133998
rect 325785 133995 325851 133998
rect 213913 133922 213979 133925
rect 213913 133920 217212 133922
rect 213913 133864 213918 133920
rect 213974 133864 217212 133920
rect 213913 133862 217212 133864
rect 213913 133859 213979 133862
rect 251950 133786 251956 133788
rect 248860 133726 251956 133786
rect 251950 133724 251956 133726
rect 252020 133724 252026 133788
rect 307661 133650 307727 133653
rect 307661 133648 310132 133650
rect 307661 133592 307666 133648
rect 307722 133592 310132 133648
rect 307661 133590 310132 133592
rect 307661 133587 307727 133590
rect 213913 133378 213979 133381
rect 251449 133378 251515 133381
rect 213913 133376 217212 133378
rect 213913 133320 213918 133376
rect 213974 133320 217212 133376
rect 213913 133318 217212 133320
rect 248860 133376 251515 133378
rect 248860 133320 251454 133376
rect 251510 133320 251515 133376
rect 248860 133318 251515 133320
rect 213913 133315 213979 133318
rect 251449 133315 251515 133318
rect 307477 133242 307543 133245
rect 324313 133242 324379 133245
rect 307477 133240 310132 133242
rect 307477 133184 307482 133240
rect 307538 133184 310132 133240
rect 307477 133182 310132 133184
rect 321908 133240 324379 133242
rect 321908 133184 324318 133240
rect 324374 133184 324379 133240
rect 321908 133182 324379 133184
rect 307477 133179 307543 133182
rect 324313 133179 324379 133182
rect 269941 133106 270007 133109
rect 307702 133106 307708 133108
rect 269941 133104 307708 133106
rect 269941 133048 269946 133104
rect 270002 133048 307708 133104
rect 269941 133046 307708 133048
rect 269941 133043 270007 133046
rect 307702 133044 307708 133046
rect 307772 133044 307778 133108
rect 252461 132834 252527 132837
rect 248860 132832 252527 132834
rect 248860 132776 252466 132832
rect 252522 132776 252527 132832
rect 248860 132774 252527 132776
rect 252461 132771 252527 132774
rect 200070 132638 217212 132698
rect 170254 132500 170260 132564
rect 170324 132562 170330 132564
rect 200070 132562 200130 132638
rect 306966 132636 306972 132700
rect 307036 132698 307042 132700
rect 307036 132638 310132 132698
rect 307036 132636 307042 132638
rect 170324 132502 200130 132562
rect 170324 132500 170330 132502
rect 251357 132426 251423 132429
rect 324313 132426 324379 132429
rect 248860 132424 251423 132426
rect 248860 132368 251362 132424
rect 251418 132368 251423 132424
rect 248860 132366 251423 132368
rect 321908 132424 324379 132426
rect 321908 132368 324318 132424
rect 324374 132368 324379 132424
rect 321908 132366 324379 132368
rect 251357 132363 251423 132366
rect 324313 132363 324379 132366
rect 307477 132290 307543 132293
rect 307477 132288 310132 132290
rect 307477 132232 307482 132288
rect 307538 132232 310132 132288
rect 307477 132230 310132 132232
rect 307477 132227 307543 132230
rect 213913 132018 213979 132021
rect 213913 132016 217212 132018
rect 213913 131960 213918 132016
rect 213974 131960 217212 132016
rect 213913 131958 217212 131960
rect 213913 131955 213979 131958
rect 252277 131882 252343 131885
rect 248860 131880 252343 131882
rect 248860 131824 252282 131880
rect 252338 131824 252343 131880
rect 248860 131822 252343 131824
rect 252277 131819 252343 131822
rect 307661 131882 307727 131885
rect 307661 131880 310132 131882
rect 307661 131824 307666 131880
rect 307722 131824 310132 131880
rect 307661 131822 310132 131824
rect 307661 131819 307727 131822
rect 324497 131746 324563 131749
rect 321908 131744 324563 131746
rect 321908 131688 324502 131744
rect 324558 131688 324563 131744
rect 321908 131686 324563 131688
rect 324497 131683 324563 131686
rect 252001 131474 252067 131477
rect 248860 131472 252067 131474
rect 248860 131416 252006 131472
rect 252062 131416 252067 131472
rect 248860 131414 252067 131416
rect 252001 131411 252067 131414
rect 306741 131474 306807 131477
rect 306741 131472 310132 131474
rect 306741 131416 306746 131472
rect 306802 131416 310132 131472
rect 306741 131414 310132 131416
rect 306741 131411 306807 131414
rect 200070 131278 217212 131338
rect 166390 131140 166396 131204
rect 166460 131202 166466 131204
rect 200070 131202 200130 131278
rect 166460 131142 200130 131202
rect 166460 131140 166466 131142
rect 306741 131066 306807 131069
rect 306741 131064 310132 131066
rect 306741 131008 306746 131064
rect 306802 131008 310132 131064
rect 306741 131006 310132 131008
rect 306741 131003 306807 131006
rect 252461 130930 252527 130933
rect 324313 130930 324379 130933
rect 248860 130928 252527 130930
rect 248860 130872 252466 130928
rect 252522 130872 252527 130928
rect 248860 130870 252527 130872
rect 321908 130928 324379 130930
rect 321908 130872 324318 130928
rect 324374 130872 324379 130928
rect 321908 130870 324379 130872
rect 252461 130867 252527 130870
rect 324313 130867 324379 130870
rect 213913 130658 213979 130661
rect 213913 130656 217212 130658
rect 213913 130600 213918 130656
rect 213974 130600 217212 130656
rect 213913 130598 217212 130600
rect 213913 130595 213979 130598
rect 301446 130596 301452 130660
rect 301516 130658 301522 130660
rect 301516 130598 310132 130658
rect 301516 130596 301522 130598
rect 251725 130522 251791 130525
rect 248860 130520 251791 130522
rect 248860 130464 251730 130520
rect 251786 130464 251791 130520
rect 248860 130462 251791 130464
rect 251725 130459 251791 130462
rect 306925 130250 306991 130253
rect 306925 130248 310132 130250
rect 306925 130192 306930 130248
rect 306986 130192 310132 130248
rect 306925 130190 310132 130192
rect 306925 130187 306991 130190
rect 252001 130114 252067 130117
rect 324405 130114 324471 130117
rect 248860 130112 252067 130114
rect 248860 130056 252006 130112
rect 252062 130056 252067 130112
rect 248860 130054 252067 130056
rect 321908 130112 324471 130114
rect 321908 130056 324410 130112
rect 324466 130056 324471 130112
rect 321908 130054 324471 130056
rect 252001 130051 252067 130054
rect 324405 130051 324471 130054
rect 200070 129918 217212 129978
rect 171726 129780 171732 129844
rect 171796 129842 171802 129844
rect 200070 129842 200130 129918
rect 171796 129782 200130 129842
rect 307661 129842 307727 129845
rect 307661 129840 310132 129842
rect 307661 129784 307666 129840
rect 307722 129784 310132 129840
rect 307661 129782 310132 129784
rect 171796 129780 171802 129782
rect 307661 129779 307727 129782
rect 252001 129570 252067 129573
rect 248860 129568 252067 129570
rect 248860 129512 252006 129568
rect 252062 129512 252067 129568
rect 248860 129510 252067 129512
rect 252001 129507 252067 129510
rect 327206 129434 327212 129436
rect 321908 129374 327212 129434
rect 327206 129372 327212 129374
rect 327276 129372 327282 129436
rect 67357 129298 67423 129301
rect 68142 129298 68816 129304
rect 67357 129296 68816 129298
rect 67357 129240 67362 129296
rect 67418 129244 68816 129296
rect 67418 129240 68202 129244
rect 67357 129238 68202 129240
rect 67357 129235 67423 129238
rect 214005 129298 214071 129301
rect 307477 129298 307543 129301
rect 214005 129296 217212 129298
rect 214005 129240 214010 129296
rect 214066 129240 217212 129296
rect 214005 129238 217212 129240
rect 307477 129296 310132 129298
rect 307477 129240 307482 129296
rect 307538 129240 310132 129296
rect 307477 129238 310132 129240
rect 214005 129235 214071 129238
rect 307477 129235 307543 129238
rect 251725 129162 251791 129165
rect 248860 129160 251791 129162
rect 248860 129104 251730 129160
rect 251786 129104 251791 129160
rect 248860 129102 251791 129104
rect 251725 129099 251791 129102
rect 307569 128890 307635 128893
rect 307569 128888 310132 128890
rect 307569 128832 307574 128888
rect 307630 128832 310132 128888
rect 307569 128830 310132 128832
rect 307569 128827 307635 128830
rect 213913 128754 213979 128757
rect 213913 128752 217212 128754
rect 213913 128696 213918 128752
rect 213974 128696 217212 128752
rect 213913 128694 217212 128696
rect 213913 128691 213979 128694
rect 252093 128618 252159 128621
rect 324313 128618 324379 128621
rect 248860 128616 252159 128618
rect 248860 128560 252098 128616
rect 252154 128560 252159 128616
rect 248860 128558 252159 128560
rect 321908 128616 324379 128618
rect 321908 128560 324318 128616
rect 324374 128560 324379 128616
rect 321908 128558 324379 128560
rect 252093 128555 252159 128558
rect 324313 128555 324379 128558
rect 307661 128482 307727 128485
rect 307661 128480 310132 128482
rect 307661 128424 307666 128480
rect 307722 128424 310132 128480
rect 307661 128422 310132 128424
rect 307661 128419 307727 128422
rect 252461 128210 252527 128213
rect 248860 128208 252527 128210
rect 248860 128152 252466 128208
rect 252522 128152 252527 128208
rect 248860 128150 252527 128152
rect 252461 128147 252527 128150
rect 67633 128074 67699 128077
rect 68142 128074 68816 128080
rect 67633 128072 68816 128074
rect 67633 128016 67638 128072
rect 67694 128020 68816 128072
rect 67694 128016 68202 128020
rect 67633 128014 68202 128016
rect 67633 128011 67699 128014
rect 214005 128074 214071 128077
rect 307477 128074 307543 128077
rect 214005 128072 217212 128074
rect 214005 128016 214010 128072
rect 214066 128016 217212 128072
rect 214005 128014 217212 128016
rect 307477 128072 310132 128074
rect 307477 128016 307482 128072
rect 307538 128016 310132 128072
rect 307477 128014 310132 128016
rect 214005 128011 214071 128014
rect 307477 128011 307543 128014
rect 324313 127802 324379 127805
rect 321908 127800 324379 127802
rect 321908 127744 324318 127800
rect 324374 127744 324379 127800
rect 321908 127742 324379 127744
rect 324313 127739 324379 127742
rect 251541 127666 251607 127669
rect 248860 127664 251607 127666
rect 248860 127608 251546 127664
rect 251602 127608 251607 127664
rect 248860 127606 251607 127608
rect 251541 127603 251607 127606
rect 307569 127666 307635 127669
rect 307569 127664 310132 127666
rect 307569 127608 307574 127664
rect 307630 127608 310132 127664
rect 307569 127606 310132 127608
rect 307569 127603 307635 127606
rect 213913 127394 213979 127397
rect 213913 127392 217212 127394
rect 213913 127336 213918 127392
rect 213974 127336 217212 127392
rect 213913 127334 217212 127336
rect 213913 127331 213979 127334
rect 252001 127258 252067 127261
rect 248860 127256 252067 127258
rect 248860 127200 252006 127256
rect 252062 127200 252067 127256
rect 248860 127198 252067 127200
rect 252001 127195 252067 127198
rect 307661 127258 307727 127261
rect 307661 127256 310132 127258
rect 307661 127200 307666 127256
rect 307722 127200 310132 127256
rect 307661 127198 310132 127200
rect 307661 127195 307727 127198
rect 329782 127122 329788 127124
rect 321908 127062 329788 127122
rect 329782 127060 329788 127062
rect 329852 127060 329858 127124
rect 307477 126850 307543 126853
rect 307477 126848 310132 126850
rect 307477 126792 307482 126848
rect 307538 126792 310132 126848
rect 307477 126790 310132 126792
rect 307477 126787 307543 126790
rect 214005 126714 214071 126717
rect 252461 126714 252527 126717
rect 214005 126712 217212 126714
rect 214005 126656 214010 126712
rect 214066 126656 217212 126712
rect 214005 126654 217212 126656
rect 248860 126712 252527 126714
rect 248860 126656 252466 126712
rect 252522 126656 252527 126712
rect 248860 126654 252527 126656
rect 214005 126651 214071 126654
rect 252461 126651 252527 126654
rect 307661 126442 307727 126445
rect 307661 126440 310132 126442
rect 307661 126384 307666 126440
rect 307722 126384 310132 126440
rect 307661 126382 310132 126384
rect 307661 126379 307727 126382
rect 64965 126306 65031 126309
rect 68142 126306 68816 126312
rect 64965 126304 68816 126306
rect 64965 126248 64970 126304
rect 65026 126252 68816 126304
rect 251909 126306 251975 126309
rect 324313 126306 324379 126309
rect 65026 126248 68202 126252
rect 64965 126246 68202 126248
rect 64965 126243 65031 126246
rect 64689 125626 64755 125629
rect 64965 125626 65031 125629
rect 64689 125624 65031 125626
rect 64689 125568 64694 125624
rect 64750 125568 64970 125624
rect 65026 125568 65031 125624
rect 64689 125566 65031 125568
rect 64689 125563 64755 125566
rect 64965 125563 65031 125566
rect 248860 126304 251975 126306
rect 248860 126248 251914 126304
rect 251970 126248 251975 126304
rect 248860 126246 251975 126248
rect 321908 126304 324379 126306
rect 321908 126248 324318 126304
rect 324374 126248 324379 126304
rect 321908 126246 324379 126248
rect 251909 126243 251975 126246
rect 324313 126243 324379 126246
rect 213913 126034 213979 126037
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 213913 126032 217212 126034
rect 213913 125976 213918 126032
rect 213974 125976 217212 126032
rect 213913 125974 217212 125976
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 213913 125971 213979 125974
rect 580165 125971 580231 125974
rect 306741 125898 306807 125901
rect 306741 125896 310132 125898
rect 306741 125840 306746 125896
rect 306802 125840 310132 125896
rect 583520 125884 584960 125974
rect 306741 125838 310132 125840
rect 306741 125835 306807 125838
rect 252093 125762 252159 125765
rect 248860 125760 252159 125762
rect 248860 125704 252098 125760
rect 252154 125704 252159 125760
rect 248860 125702 252159 125704
rect 252093 125699 252159 125702
rect 306741 125490 306807 125493
rect 324497 125490 324563 125493
rect 306741 125488 310132 125490
rect 306741 125432 306746 125488
rect 306802 125432 310132 125488
rect 306741 125430 310132 125432
rect 321908 125488 324563 125490
rect 321908 125432 324502 125488
rect 324558 125432 324563 125488
rect 321908 125430 324563 125432
rect 306741 125427 306807 125430
rect 324497 125427 324563 125430
rect 214005 125354 214071 125357
rect 252461 125354 252527 125357
rect 214005 125352 217212 125354
rect 214005 125296 214010 125352
rect 214066 125296 217212 125352
rect 214005 125294 217212 125296
rect 248860 125352 252527 125354
rect 248860 125296 252466 125352
rect 252522 125296 252527 125352
rect 248860 125294 252527 125296
rect 214005 125291 214071 125294
rect 252461 125291 252527 125294
rect 66161 125218 66227 125221
rect 68142 125218 68816 125224
rect 66161 125216 68816 125218
rect 66161 125160 66166 125216
rect 66222 125164 68816 125216
rect 66222 125160 68202 125164
rect 66161 125158 68202 125160
rect 66161 125155 66227 125158
rect -960 123572 480 123812
rect 307477 125082 307543 125085
rect 307477 125080 310132 125082
rect 307477 125024 307482 125080
rect 307538 125024 310132 125080
rect 307477 125022 310132 125024
rect 307477 125019 307543 125022
rect 252369 124810 252435 124813
rect 325601 124810 325667 124813
rect 248860 124808 252435 124810
rect 248860 124752 252374 124808
rect 252430 124752 252435 124808
rect 248860 124750 252435 124752
rect 321908 124808 325667 124810
rect 321908 124752 325606 124808
rect 325662 124752 325667 124808
rect 321908 124750 325667 124752
rect 252369 124747 252435 124750
rect 325601 124747 325667 124750
rect 213913 124674 213979 124677
rect 307293 124674 307359 124677
rect 213913 124672 217212 124674
rect 213913 124616 213918 124672
rect 213974 124616 217212 124672
rect 213913 124614 217212 124616
rect 307293 124672 310132 124674
rect 307293 124616 307298 124672
rect 307354 124616 310132 124672
rect 307293 124614 310132 124616
rect 213913 124611 213979 124614
rect 307293 124611 307359 124614
rect 251265 124402 251331 124405
rect 248860 124400 251331 124402
rect 248860 124344 251270 124400
rect 251326 124344 251331 124400
rect 248860 124342 251331 124344
rect 251265 124339 251331 124342
rect 307661 124266 307727 124269
rect 307661 124264 310132 124266
rect 307661 124208 307666 124264
rect 307722 124208 310132 124264
rect 307661 124206 310132 124208
rect 307661 124203 307727 124206
rect 214005 124130 214071 124133
rect 214005 124128 217212 124130
rect 214005 124072 214010 124128
rect 214066 124072 217212 124128
rect 214005 124070 217212 124072
rect 214005 124067 214071 124070
rect 252277 123994 252343 123997
rect 324313 123994 324379 123997
rect 248860 123992 252343 123994
rect 248860 123936 252282 123992
rect 252338 123936 252343 123992
rect 248860 123934 252343 123936
rect 321908 123992 324379 123994
rect 321908 123936 324318 123992
rect 324374 123936 324379 123992
rect 321908 123934 324379 123936
rect 252277 123931 252343 123934
rect 324313 123931 324379 123934
rect 306557 123858 306623 123861
rect 306557 123856 310132 123858
rect 306557 123800 306562 123856
rect 306618 123800 310132 123856
rect 306557 123798 310132 123800
rect 306557 123795 306623 123798
rect 66069 123586 66135 123589
rect 68142 123586 68816 123592
rect 66069 123584 68816 123586
rect 66069 123528 66074 123584
rect 66130 123532 68816 123584
rect 66130 123528 68202 123532
rect 66069 123526 68202 123528
rect 66069 123523 66135 123526
rect 213913 123450 213979 123453
rect 252461 123450 252527 123453
rect 213913 123448 217212 123450
rect 213913 123392 213918 123448
rect 213974 123392 217212 123448
rect 213913 123390 217212 123392
rect 248860 123448 252527 123450
rect 248860 123392 252466 123448
rect 252522 123392 252527 123448
rect 248860 123390 252527 123392
rect 213913 123387 213979 123390
rect 252461 123387 252527 123390
rect 307569 123450 307635 123453
rect 307569 123448 310132 123450
rect 307569 123392 307574 123448
rect 307630 123392 310132 123448
rect 307569 123390 310132 123392
rect 307569 123387 307635 123390
rect 324957 123178 325023 123181
rect 321908 123176 325023 123178
rect 321908 123120 324962 123176
rect 325018 123120 325023 123176
rect 321908 123118 325023 123120
rect 324957 123115 325023 123118
rect 252001 123042 252067 123045
rect 248860 123040 252067 123042
rect 248860 122984 252006 123040
rect 252062 122984 252067 123040
rect 248860 122982 252067 122984
rect 252001 122979 252067 122982
rect 307661 123042 307727 123045
rect 307661 123040 310132 123042
rect 307661 122984 307666 123040
rect 307722 122984 310132 123040
rect 307661 122982 310132 122984
rect 307661 122979 307727 122982
rect 214005 122770 214071 122773
rect 214005 122768 217212 122770
rect 214005 122712 214010 122768
rect 214066 122712 217212 122768
rect 214005 122710 217212 122712
rect 214005 122707 214071 122710
rect 67449 122634 67515 122637
rect 68142 122634 68816 122640
rect 67449 122632 68816 122634
rect 67449 122576 67454 122632
rect 67510 122580 68816 122632
rect 67510 122576 68202 122580
rect 67449 122574 68202 122576
rect 67449 122571 67515 122574
rect 252461 122498 252527 122501
rect 248860 122496 252527 122498
rect 248860 122440 252466 122496
rect 252522 122440 252527 122496
rect 248860 122438 252527 122440
rect 252461 122435 252527 122438
rect 307477 122498 307543 122501
rect 324681 122498 324747 122501
rect 307477 122496 310132 122498
rect 307477 122440 307482 122496
rect 307538 122440 310132 122496
rect 307477 122438 310132 122440
rect 321908 122496 324747 122498
rect 321908 122440 324686 122496
rect 324742 122440 324747 122496
rect 321908 122438 324747 122440
rect 307477 122435 307543 122438
rect 324681 122435 324747 122438
rect 213913 122090 213979 122093
rect 252369 122090 252435 122093
rect 213913 122088 217212 122090
rect 213913 122032 213918 122088
rect 213974 122032 217212 122088
rect 213913 122030 217212 122032
rect 248860 122088 252435 122090
rect 248860 122032 252374 122088
rect 252430 122032 252435 122088
rect 248860 122030 252435 122032
rect 213913 122027 213979 122030
rect 252369 122027 252435 122030
rect 307569 122090 307635 122093
rect 307569 122088 310132 122090
rect 307569 122032 307574 122088
rect 307630 122032 310132 122088
rect 307569 122030 310132 122032
rect 307569 122027 307635 122030
rect 307661 121682 307727 121685
rect 324313 121682 324379 121685
rect 307661 121680 310132 121682
rect 307661 121624 307666 121680
rect 307722 121624 310132 121680
rect 307661 121622 310132 121624
rect 321908 121680 324379 121682
rect 321908 121624 324318 121680
rect 324374 121624 324379 121680
rect 321908 121622 324379 121624
rect 307661 121619 307727 121622
rect 324313 121619 324379 121622
rect 252461 121546 252527 121549
rect 248860 121544 252527 121546
rect 248860 121488 252466 121544
rect 252522 121488 252527 121544
rect 248860 121486 252527 121488
rect 252461 121483 252527 121486
rect 214005 121410 214071 121413
rect 214005 121408 217212 121410
rect 214005 121352 214010 121408
rect 214066 121352 217212 121408
rect 214005 121350 217212 121352
rect 214005 121347 214071 121350
rect 307477 121274 307543 121277
rect 307477 121272 310132 121274
rect 307477 121216 307482 121272
rect 307538 121216 310132 121272
rect 307477 121214 310132 121216
rect 307477 121211 307543 121214
rect 252461 121138 252527 121141
rect 248860 121136 252527 121138
rect 248860 121080 252466 121136
rect 252522 121080 252527 121136
rect 248860 121078 252527 121080
rect 252461 121075 252527 121078
rect 67541 120866 67607 120869
rect 68142 120866 68816 120872
rect 67541 120864 68816 120866
rect 67541 120808 67546 120864
rect 67602 120812 68816 120864
rect 67602 120808 68202 120812
rect 67541 120806 68202 120808
rect 67541 120803 67607 120806
rect 307569 120866 307635 120869
rect 324313 120866 324379 120869
rect 307569 120864 310132 120866
rect 307569 120808 307574 120864
rect 307630 120808 310132 120864
rect 307569 120806 310132 120808
rect 321908 120864 324379 120866
rect 321908 120808 324318 120864
rect 324374 120808 324379 120864
rect 321908 120806 324379 120808
rect 307569 120803 307635 120806
rect 324313 120803 324379 120806
rect 213913 120730 213979 120733
rect 213913 120728 217212 120730
rect 213913 120672 213918 120728
rect 213974 120672 217212 120728
rect 213913 120670 217212 120672
rect 213913 120667 213979 120670
rect 252369 120594 252435 120597
rect 248860 120592 252435 120594
rect 248860 120536 252374 120592
rect 252430 120536 252435 120592
rect 248860 120534 252435 120536
rect 252369 120531 252435 120534
rect 307661 120458 307727 120461
rect 307661 120456 310132 120458
rect 307661 120400 307666 120456
rect 307722 120400 310132 120456
rect 307661 120398 310132 120400
rect 307661 120395 307727 120398
rect 251909 120186 251975 120189
rect 324405 120186 324471 120189
rect 248860 120184 251975 120186
rect 248860 120128 251914 120184
rect 251970 120128 251975 120184
rect 248860 120126 251975 120128
rect 321908 120184 324471 120186
rect 321908 120128 324410 120184
rect 324466 120128 324471 120184
rect 321908 120126 324471 120128
rect 251909 120123 251975 120126
rect 324405 120123 324471 120126
rect 214005 120050 214071 120053
rect 306741 120050 306807 120053
rect 214005 120048 217212 120050
rect 214005 119992 214010 120048
rect 214066 119992 217212 120048
rect 214005 119990 217212 119992
rect 306741 120048 310132 120050
rect 306741 119992 306746 120048
rect 306802 119992 310132 120048
rect 306741 119990 310132 119992
rect 214005 119987 214071 119990
rect 306741 119987 306807 119990
rect 251357 119642 251423 119645
rect 248860 119640 251423 119642
rect 248860 119584 251362 119640
rect 251418 119584 251423 119640
rect 248860 119582 251423 119584
rect 251357 119579 251423 119582
rect 307569 119642 307635 119645
rect 307569 119640 310132 119642
rect 307569 119584 307574 119640
rect 307630 119584 310132 119640
rect 307569 119582 310132 119584
rect 307569 119579 307635 119582
rect 214097 119506 214163 119509
rect 214097 119504 217212 119506
rect 214097 119448 214102 119504
rect 214158 119448 217212 119504
rect 214097 119446 217212 119448
rect 214097 119443 214163 119446
rect 324497 119370 324563 119373
rect 321908 119368 324563 119370
rect 321908 119312 324502 119368
rect 324558 119312 324563 119368
rect 321908 119310 324563 119312
rect 324497 119307 324563 119310
rect 251817 119234 251883 119237
rect 248860 119232 251883 119234
rect 248860 119176 251822 119232
rect 251878 119176 251883 119232
rect 248860 119174 251883 119176
rect 251817 119171 251883 119174
rect 307661 119098 307727 119101
rect 307661 119096 310132 119098
rect 307661 119040 307666 119096
rect 307722 119040 310132 119096
rect 307661 119038 310132 119040
rect 307661 119035 307727 119038
rect 305729 118962 305795 118965
rect 307569 118962 307635 118965
rect 305729 118960 307635 118962
rect 305729 118904 305734 118960
rect 305790 118904 307574 118960
rect 307630 118904 307635 118960
rect 305729 118902 307635 118904
rect 305729 118899 305795 118902
rect 307569 118899 307635 118902
rect 213913 118826 213979 118829
rect 252461 118826 252527 118829
rect 213913 118824 217212 118826
rect 213913 118768 213918 118824
rect 213974 118768 217212 118824
rect 213913 118766 217212 118768
rect 248860 118824 252527 118826
rect 248860 118768 252466 118824
rect 252522 118768 252527 118824
rect 248860 118766 252527 118768
rect 213913 118763 213979 118766
rect 252461 118763 252527 118766
rect 307477 118690 307543 118693
rect 307477 118688 310132 118690
rect 307477 118632 307482 118688
rect 307538 118632 310132 118688
rect 307477 118630 310132 118632
rect 307477 118627 307543 118630
rect 324313 118554 324379 118557
rect 321908 118552 324379 118554
rect 321908 118496 324318 118552
rect 324374 118496 324379 118552
rect 321908 118494 324379 118496
rect 324313 118491 324379 118494
rect 252461 118282 252527 118285
rect 248860 118280 252527 118282
rect 248860 118224 252466 118280
rect 252522 118224 252527 118280
rect 248860 118222 252527 118224
rect 252461 118219 252527 118222
rect 304206 118220 304212 118284
rect 304276 118282 304282 118284
rect 304276 118222 310132 118282
rect 304276 118220 304282 118222
rect 213913 118146 213979 118149
rect 213913 118144 217212 118146
rect 213913 118088 213918 118144
rect 213974 118088 217212 118144
rect 213913 118086 217212 118088
rect 213913 118083 213979 118086
rect 251817 117874 251883 117877
rect 248860 117872 251883 117874
rect 248860 117816 251822 117872
rect 251878 117816 251883 117872
rect 248860 117814 251883 117816
rect 251817 117811 251883 117814
rect 307569 117874 307635 117877
rect 324405 117874 324471 117877
rect 307569 117872 310132 117874
rect 307569 117816 307574 117872
rect 307630 117816 310132 117872
rect 307569 117814 310132 117816
rect 321908 117872 324471 117874
rect 321908 117816 324410 117872
rect 324466 117816 324471 117872
rect 321908 117814 324471 117816
rect 307569 117811 307635 117814
rect 324405 117811 324471 117814
rect 213177 117466 213243 117469
rect 307661 117466 307727 117469
rect 213177 117464 217212 117466
rect 213177 117408 213182 117464
rect 213238 117408 217212 117464
rect 213177 117406 217212 117408
rect 307661 117464 310132 117466
rect 307661 117408 307666 117464
rect 307722 117408 310132 117464
rect 307661 117406 310132 117408
rect 213177 117403 213243 117406
rect 307661 117403 307727 117406
rect 251173 117330 251239 117333
rect 248860 117328 251239 117330
rect 248860 117272 251178 117328
rect 251234 117272 251239 117328
rect 248860 117270 251239 117272
rect 251173 117267 251239 117270
rect 307661 117058 307727 117061
rect 324313 117058 324379 117061
rect 307661 117056 310132 117058
rect 307661 117000 307666 117056
rect 307722 117000 310132 117056
rect 307661 116998 310132 117000
rect 321908 117056 324379 117058
rect 321908 117000 324318 117056
rect 324374 117000 324379 117056
rect 321908 116998 324379 117000
rect 307661 116995 307727 116998
rect 324313 116995 324379 116998
rect 252461 116922 252527 116925
rect 248860 116920 252527 116922
rect 248860 116864 252466 116920
rect 252522 116864 252527 116920
rect 248860 116862 252527 116864
rect 252461 116859 252527 116862
rect 214005 116786 214071 116789
rect 214005 116784 217212 116786
rect 214005 116728 214010 116784
rect 214066 116728 217212 116784
rect 214005 116726 217212 116728
rect 214005 116723 214071 116726
rect 306741 116650 306807 116653
rect 306741 116648 310132 116650
rect 306741 116592 306746 116648
rect 306802 116592 310132 116648
rect 306741 116590 310132 116592
rect 306741 116587 306807 116590
rect 251909 116378 251975 116381
rect 324405 116378 324471 116381
rect 248860 116376 251975 116378
rect 248860 116320 251914 116376
rect 251970 116320 251975 116376
rect 248860 116318 251975 116320
rect 321908 116376 324471 116378
rect 321908 116320 324410 116376
rect 324466 116320 324471 116376
rect 321908 116318 324471 116320
rect 251909 116315 251975 116318
rect 324405 116315 324471 116318
rect 307201 116242 307267 116245
rect 307201 116240 310132 116242
rect 307201 116184 307206 116240
rect 307262 116184 310132 116240
rect 307201 116182 310132 116184
rect 307201 116179 307267 116182
rect 213913 116106 213979 116109
rect 213913 116104 217212 116106
rect 213913 116048 213918 116104
rect 213974 116048 217212 116104
rect 213913 116046 217212 116048
rect 213913 116043 213979 116046
rect 252369 115970 252435 115973
rect 248860 115968 252435 115970
rect 248860 115912 252374 115968
rect 252430 115912 252435 115968
rect 248860 115910 252435 115912
rect 252369 115907 252435 115910
rect 306741 115698 306807 115701
rect 306741 115696 310132 115698
rect 306741 115640 306746 115696
rect 306802 115640 310132 115696
rect 306741 115638 310132 115640
rect 306741 115635 306807 115638
rect 324313 115562 324379 115565
rect 321908 115560 324379 115562
rect 321908 115504 324318 115560
rect 324374 115504 324379 115560
rect 321908 115502 324379 115504
rect 324313 115499 324379 115502
rect 214005 115426 214071 115429
rect 252461 115426 252527 115429
rect 214005 115424 217212 115426
rect 214005 115368 214010 115424
rect 214066 115368 217212 115424
rect 214005 115366 217212 115368
rect 248860 115424 252527 115426
rect 248860 115368 252466 115424
rect 252522 115368 252527 115424
rect 248860 115366 252527 115368
rect 214005 115363 214071 115366
rect 252461 115363 252527 115366
rect 297214 115228 297220 115292
rect 297284 115290 297290 115292
rect 297284 115230 310132 115290
rect 297284 115228 297290 115230
rect 252369 115018 252435 115021
rect 248860 115016 252435 115018
rect 248860 114960 252374 115016
rect 252430 114960 252435 115016
rect 248860 114958 252435 114960
rect 252369 114955 252435 114958
rect 213913 114882 213979 114885
rect 307661 114882 307727 114885
rect 213913 114880 217212 114882
rect 213913 114824 213918 114880
rect 213974 114824 217212 114880
rect 213913 114822 217212 114824
rect 307661 114880 310132 114882
rect 307661 114824 307666 114880
rect 307722 114824 310132 114880
rect 307661 114822 310132 114824
rect 213913 114819 213979 114822
rect 307661 114819 307727 114822
rect 321908 114686 325710 114746
rect 325650 114610 325710 114686
rect 338246 114610 338252 114612
rect 325650 114550 338252 114610
rect 338246 114548 338252 114550
rect 338316 114548 338322 114612
rect 251633 114474 251699 114477
rect 248860 114472 251699 114474
rect 248860 114416 251638 114472
rect 251694 114416 251699 114472
rect 248860 114414 251699 114416
rect 251633 114411 251699 114414
rect 306741 114474 306807 114477
rect 306741 114472 310132 114474
rect 306741 114416 306746 114472
rect 306802 114416 310132 114472
rect 306741 114414 310132 114416
rect 306741 114411 306807 114414
rect 214005 114202 214071 114205
rect 214005 114200 217212 114202
rect 214005 114144 214010 114200
rect 214066 114144 217212 114200
rect 214005 114142 217212 114144
rect 214005 114139 214071 114142
rect 252461 114066 252527 114069
rect 248860 114064 252527 114066
rect 248860 114008 252466 114064
rect 252522 114008 252527 114064
rect 248860 114006 252527 114008
rect 252461 114003 252527 114006
rect 307150 114004 307156 114068
rect 307220 114066 307226 114068
rect 324313 114066 324379 114069
rect 307220 114006 310132 114066
rect 321908 114064 324379 114066
rect 321908 114008 324318 114064
rect 324374 114008 324379 114064
rect 321908 114006 324379 114008
rect 307220 114004 307226 114006
rect 324313 114003 324379 114006
rect 307569 113658 307635 113661
rect 307569 113656 310132 113658
rect 307569 113600 307574 113656
rect 307630 113600 310132 113656
rect 307569 113598 310132 113600
rect 307569 113595 307635 113598
rect 213913 113522 213979 113525
rect 252369 113522 252435 113525
rect 213913 113520 217212 113522
rect 213913 113464 213918 113520
rect 213974 113464 217212 113520
rect 213913 113462 217212 113464
rect 248860 113520 252435 113522
rect 248860 113464 252374 113520
rect 252430 113464 252435 113520
rect 248860 113462 252435 113464
rect 213913 113459 213979 113462
rect 252369 113459 252435 113462
rect 307661 113250 307727 113253
rect 324405 113250 324471 113253
rect 307661 113248 310132 113250
rect 307661 113192 307666 113248
rect 307722 113192 310132 113248
rect 307661 113190 310132 113192
rect 321908 113248 324471 113250
rect 321908 113192 324410 113248
rect 324466 113192 324471 113248
rect 321908 113190 324471 113192
rect 307661 113187 307727 113190
rect 324405 113187 324471 113190
rect 252093 113114 252159 113117
rect 248860 113112 252159 113114
rect 248860 113056 252098 113112
rect 252154 113056 252159 113112
rect 248860 113054 252159 113056
rect 252093 113051 252159 113054
rect 214005 112842 214071 112845
rect 582649 112842 582715 112845
rect 583520 112842 584960 112932
rect 214005 112840 217212 112842
rect 214005 112784 214010 112840
rect 214066 112784 217212 112840
rect 214005 112782 217212 112784
rect 582649 112840 584960 112842
rect 582649 112784 582654 112840
rect 582710 112784 584960 112840
rect 582649 112782 584960 112784
rect 214005 112779 214071 112782
rect 582649 112779 582715 112782
rect 252001 112706 252067 112709
rect 248860 112704 252067 112706
rect 248860 112648 252006 112704
rect 252062 112648 252067 112704
rect 248860 112646 252067 112648
rect 252001 112643 252067 112646
rect 305494 112644 305500 112708
rect 305564 112706 305570 112708
rect 305564 112646 310132 112706
rect 583520 112692 584960 112782
rect 305564 112644 305570 112646
rect 324313 112434 324379 112437
rect 321908 112432 324379 112434
rect 321908 112376 324318 112432
rect 324374 112376 324379 112432
rect 321908 112374 324379 112376
rect 324313 112371 324379 112374
rect 307569 112298 307635 112301
rect 307569 112296 310132 112298
rect 307569 112240 307574 112296
rect 307630 112240 310132 112296
rect 307569 112238 310132 112240
rect 307569 112235 307635 112238
rect 213913 112162 213979 112165
rect 252461 112162 252527 112165
rect 213913 112160 217212 112162
rect 213913 112104 213918 112160
rect 213974 112104 217212 112160
rect 213913 112102 217212 112104
rect 248860 112160 252527 112162
rect 248860 112104 252466 112160
rect 252522 112104 252527 112160
rect 248860 112102 252527 112104
rect 213913 112099 213979 112102
rect 252461 112099 252527 112102
rect 307661 111890 307727 111893
rect 307661 111888 310132 111890
rect 307661 111832 307666 111888
rect 307722 111832 310132 111888
rect 307661 111830 310132 111832
rect 307661 111827 307727 111830
rect 167913 111754 167979 111757
rect 252277 111754 252343 111757
rect 324313 111754 324379 111757
rect 164694 111752 167979 111754
rect 164694 111696 167918 111752
rect 167974 111696 167979 111752
rect 164694 111694 167979 111696
rect 248860 111752 252343 111754
rect 248860 111696 252282 111752
rect 252338 111696 252343 111752
rect 248860 111694 252343 111696
rect 321908 111752 324379 111754
rect 321908 111696 324318 111752
rect 324374 111696 324379 111752
rect 321908 111694 324379 111696
rect -960 110666 480 110756
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 167913 111691 167979 111694
rect 252277 111691 252343 111694
rect 324313 111691 324379 111694
rect 214005 111482 214071 111485
rect 307477 111482 307543 111485
rect 214005 111480 217212 111482
rect 214005 111424 214010 111480
rect 214066 111424 217212 111480
rect 214005 111422 217212 111424
rect 307477 111480 310132 111482
rect 307477 111424 307482 111480
rect 307538 111424 310132 111480
rect 307477 111422 310132 111424
rect 214005 111419 214071 111422
rect 307477 111419 307543 111422
rect 252461 111210 252527 111213
rect 248860 111208 252527 111210
rect 248860 111152 252466 111208
rect 252522 111152 252527 111208
rect 248860 111150 252527 111152
rect 252461 111147 252527 111150
rect 307569 111074 307635 111077
rect 307569 111072 310132 111074
rect 307569 111016 307574 111072
rect 307630 111016 310132 111072
rect 307569 111014 310132 111016
rect 307569 111011 307635 111014
rect 213913 110802 213979 110805
rect 251541 110802 251607 110805
rect 213913 110800 217212 110802
rect 213913 110744 213918 110800
rect 213974 110744 217212 110800
rect 213913 110742 217212 110744
rect 248860 110800 251607 110802
rect 248860 110744 251546 110800
rect 251602 110744 251607 110800
rect 248860 110742 251607 110744
rect 213913 110739 213979 110742
rect 251541 110739 251607 110742
rect 307661 110666 307727 110669
rect 307661 110664 310132 110666
rect 307661 110608 307666 110664
rect 307722 110608 310132 110664
rect 307661 110606 310132 110608
rect 307661 110603 307727 110606
rect 321878 110530 321938 110908
rect 336774 110530 336780 110532
rect 321878 110470 336780 110530
rect 336774 110468 336780 110470
rect 336844 110468 336850 110532
rect 213913 110258 213979 110261
rect 252461 110258 252527 110261
rect 213913 110256 217212 110258
rect 213913 110200 213918 110256
rect 213974 110200 217212 110256
rect 213913 110198 217212 110200
rect 248860 110256 252527 110258
rect 248860 110200 252466 110256
rect 252522 110200 252527 110256
rect 248860 110198 252527 110200
rect 213913 110195 213979 110198
rect 252461 110195 252527 110198
rect 307477 110258 307543 110261
rect 307477 110256 310132 110258
rect 307477 110200 307482 110256
rect 307538 110200 310132 110256
rect 307477 110198 310132 110200
rect 307477 110195 307543 110198
rect 168189 110122 168255 110125
rect 164694 110120 168255 110122
rect 164694 110064 168194 110120
rect 168250 110064 168255 110120
rect 164694 110062 168255 110064
rect 168189 110059 168255 110062
rect 252369 109850 252435 109853
rect 248860 109848 252435 109850
rect 248860 109792 252374 109848
rect 252430 109792 252435 109848
rect 248860 109790 252435 109792
rect 252369 109787 252435 109790
rect 307569 109850 307635 109853
rect 307569 109848 310132 109850
rect 307569 109792 307574 109848
rect 307630 109792 310132 109848
rect 307569 109790 310132 109792
rect 307569 109787 307635 109790
rect 321878 109578 321938 110092
rect 332726 109578 332732 109580
rect 167678 109108 167684 109172
rect 167748 109170 167754 109172
rect 217182 109170 217242 109548
rect 321878 109518 332732 109578
rect 332726 109516 332732 109518
rect 332796 109516 332802 109580
rect 251909 109306 251975 109309
rect 248860 109304 251975 109306
rect 248860 109248 251914 109304
rect 251970 109248 251975 109304
rect 248860 109246 251975 109248
rect 251909 109243 251975 109246
rect 307661 109306 307727 109309
rect 307661 109304 310132 109306
rect 307661 109248 307666 109304
rect 307722 109248 310132 109304
rect 307661 109246 310132 109248
rect 307661 109243 307727 109246
rect 167748 109110 217242 109170
rect 321878 109170 321938 109412
rect 335670 109170 335676 109172
rect 321878 109110 335676 109170
rect 167748 109108 167754 109110
rect 335670 109108 335676 109110
rect 335740 109108 335746 109172
rect 214005 108898 214071 108901
rect 252461 108898 252527 108901
rect 214005 108896 217212 108898
rect 214005 108840 214010 108896
rect 214066 108840 217212 108896
rect 214005 108838 217212 108840
rect 248860 108896 252527 108898
rect 248860 108840 252466 108896
rect 252522 108840 252527 108896
rect 248860 108838 252527 108840
rect 214005 108835 214071 108838
rect 252461 108835 252527 108838
rect 306741 108898 306807 108901
rect 306741 108896 310132 108898
rect 306741 108840 306746 108896
rect 306802 108840 310132 108896
rect 306741 108838 310132 108840
rect 306741 108835 306807 108838
rect 167729 108762 167795 108765
rect 164694 108760 167795 108762
rect 164694 108704 167734 108760
rect 167790 108704 167795 108760
rect 164694 108702 167795 108704
rect 167729 108699 167795 108702
rect 324405 108626 324471 108629
rect 321908 108624 324471 108626
rect 321908 108568 324410 108624
rect 324466 108568 324471 108624
rect 321908 108566 324471 108568
rect 324405 108563 324471 108566
rect 306005 108490 306071 108493
rect 306005 108488 310132 108490
rect 306005 108432 306010 108488
rect 306066 108432 310132 108488
rect 306005 108430 310132 108432
rect 306005 108427 306071 108430
rect 251725 108354 251791 108357
rect 248860 108352 251791 108354
rect 248860 108296 251730 108352
rect 251786 108296 251791 108352
rect 248860 108294 251791 108296
rect 251725 108291 251791 108294
rect 213913 108218 213979 108221
rect 213913 108216 217212 108218
rect 213913 108160 213918 108216
rect 213974 108160 217212 108216
rect 213913 108158 217212 108160
rect 213913 108155 213979 108158
rect 307569 108082 307635 108085
rect 307569 108080 310132 108082
rect 307569 108024 307574 108080
rect 307630 108024 310132 108080
rect 307569 108022 310132 108024
rect 307569 108019 307635 108022
rect 251357 107946 251423 107949
rect 248860 107944 251423 107946
rect 248860 107888 251362 107944
rect 251418 107888 251423 107944
rect 248860 107886 251423 107888
rect 251357 107883 251423 107886
rect 324313 107810 324379 107813
rect 321908 107808 324379 107810
rect 321908 107752 324318 107808
rect 324374 107752 324379 107808
rect 321908 107750 324379 107752
rect 324313 107747 324379 107750
rect 307661 107674 307727 107677
rect 307661 107672 310132 107674
rect 307661 107616 307666 107672
rect 307722 107616 310132 107672
rect 307661 107614 310132 107616
rect 307661 107611 307727 107614
rect 213913 107538 213979 107541
rect 251265 107538 251331 107541
rect 213913 107536 217212 107538
rect 213913 107480 213918 107536
rect 213974 107480 217212 107536
rect 213913 107478 217212 107480
rect 248860 107536 251331 107538
rect 248860 107480 251270 107536
rect 251326 107480 251331 107536
rect 248860 107478 251331 107480
rect 213913 107475 213979 107478
rect 251265 107475 251331 107478
rect 307477 107266 307543 107269
rect 307477 107264 310132 107266
rect 307477 107208 307482 107264
rect 307538 107208 310132 107264
rect 307477 107206 310132 107208
rect 307477 107203 307543 107206
rect 252461 106994 252527 106997
rect 248860 106992 252527 106994
rect 248860 106936 252466 106992
rect 252522 106936 252527 106992
rect 248860 106934 252527 106936
rect 252461 106931 252527 106934
rect 214649 106858 214715 106861
rect 307569 106858 307635 106861
rect 214649 106856 217212 106858
rect 214649 106800 214654 106856
rect 214710 106800 217212 106856
rect 214649 106798 217212 106800
rect 307569 106856 310132 106858
rect 307569 106800 307574 106856
rect 307630 106800 310132 106856
rect 307569 106798 310132 106800
rect 214649 106795 214715 106798
rect 307569 106795 307635 106798
rect 251357 106586 251423 106589
rect 248860 106584 251423 106586
rect 248860 106528 251362 106584
rect 251418 106528 251423 106584
rect 248860 106526 251423 106528
rect 321878 106586 321938 107100
rect 323485 106586 323551 106589
rect 321878 106584 323551 106586
rect 321878 106528 323490 106584
rect 323546 106528 323551 106584
rect 321878 106526 323551 106528
rect 251357 106523 251423 106526
rect 323485 106523 323551 106526
rect 307661 106450 307727 106453
rect 328494 106450 328500 106452
rect 307661 106448 310132 106450
rect 307661 106392 307666 106448
rect 307722 106392 310132 106448
rect 307661 106390 310132 106392
rect 321878 106390 328500 106450
rect 307661 106387 307727 106390
rect 321878 106284 321938 106390
rect 328494 106388 328500 106390
rect 328564 106388 328570 106452
rect 323485 106314 323551 106317
rect 342294 106314 342300 106316
rect 323485 106312 342300 106314
rect 323485 106256 323490 106312
rect 323546 106256 342300 106312
rect 323485 106254 342300 106256
rect 323485 106251 323551 106254
rect 342294 106252 342300 106254
rect 342364 106252 342370 106316
rect 214005 106178 214071 106181
rect 214005 106176 217212 106178
rect 214005 106120 214010 106176
rect 214066 106120 217212 106176
rect 214005 106118 217212 106120
rect 214005 106115 214071 106118
rect 252001 106042 252067 106045
rect 321553 106042 321619 106045
rect 248860 106040 252067 106042
rect 248860 105984 252006 106040
rect 252062 105984 252067 106040
rect 248860 105982 252067 105984
rect 252001 105979 252067 105982
rect 321510 106040 321619 106042
rect 321510 105984 321558 106040
rect 321614 105984 321619 106040
rect 321510 105979 321619 105984
rect 306557 105906 306623 105909
rect 306557 105904 310132 105906
rect 306557 105848 306562 105904
rect 306618 105848 310132 105904
rect 306557 105846 310132 105848
rect 306557 105843 306623 105846
rect 213913 105634 213979 105637
rect 252277 105634 252343 105637
rect 213913 105632 217212 105634
rect 213913 105576 213918 105632
rect 213974 105576 217212 105632
rect 213913 105574 217212 105576
rect 248860 105632 252343 105634
rect 248860 105576 252282 105632
rect 252338 105576 252343 105632
rect 248860 105574 252343 105576
rect 213913 105571 213979 105574
rect 252277 105571 252343 105574
rect 305637 105498 305703 105501
rect 305637 105496 310132 105498
rect 305637 105440 305642 105496
rect 305698 105440 310132 105496
rect 321510 105468 321570 105979
rect 305637 105438 310132 105440
rect 305637 105435 305703 105438
rect 251766 105090 251772 105092
rect 248860 105030 251772 105090
rect 251766 105028 251772 105030
rect 251836 105028 251842 105092
rect 307661 105090 307727 105093
rect 307661 105088 310132 105090
rect 307661 105032 307666 105088
rect 307722 105032 310132 105088
rect 307661 105030 310132 105032
rect 307661 105027 307727 105030
rect 214414 104892 214420 104956
rect 214484 104954 214490 104956
rect 214484 104894 217212 104954
rect 214484 104892 214490 104894
rect 324262 104818 324268 104820
rect 321908 104758 324268 104818
rect 324262 104756 324268 104758
rect 324332 104756 324338 104820
rect 252001 104682 252067 104685
rect 248860 104680 252067 104682
rect 248860 104624 252006 104680
rect 252062 104624 252067 104680
rect 248860 104622 252067 104624
rect 252001 104619 252067 104622
rect 307569 104682 307635 104685
rect 307569 104680 310132 104682
rect 307569 104624 307574 104680
rect 307630 104624 310132 104680
rect 307569 104622 310132 104624
rect 307569 104619 307635 104622
rect 213913 104274 213979 104277
rect 305821 104274 305887 104277
rect 213913 104272 217212 104274
rect 213913 104216 213918 104272
rect 213974 104216 217212 104272
rect 213913 104214 217212 104216
rect 305821 104272 310132 104274
rect 305821 104216 305826 104272
rect 305882 104216 310132 104272
rect 305821 104214 310132 104216
rect 213913 104211 213979 104214
rect 305821 104211 305887 104214
rect 252461 104138 252527 104141
rect 248860 104136 252527 104138
rect 248860 104080 252466 104136
rect 252522 104080 252527 104136
rect 248860 104078 252527 104080
rect 252461 104075 252527 104078
rect 327022 104002 327028 104004
rect 321908 103942 327028 104002
rect 327022 103940 327028 103942
rect 327092 103940 327098 104004
rect 307661 103866 307727 103869
rect 307661 103864 310132 103866
rect 307661 103808 307666 103864
rect 307722 103808 310132 103864
rect 307661 103806 310132 103808
rect 307661 103803 307727 103806
rect 251173 103730 251239 103733
rect 248860 103728 251239 103730
rect 248860 103672 251178 103728
rect 251234 103672 251239 103728
rect 248860 103670 251239 103672
rect 251173 103667 251239 103670
rect 169150 103532 169156 103596
rect 169220 103594 169226 103596
rect 169220 103534 217212 103594
rect 169220 103532 169226 103534
rect 306741 103458 306807 103461
rect 306741 103456 310132 103458
rect 306741 103400 306746 103456
rect 306802 103400 310132 103456
rect 306741 103398 310132 103400
rect 306741 103395 306807 103398
rect 252461 103186 252527 103189
rect 324313 103186 324379 103189
rect 248860 103184 252527 103186
rect 248860 103128 252466 103184
rect 252522 103128 252527 103184
rect 248860 103126 252527 103128
rect 321908 103184 324379 103186
rect 321908 103128 324318 103184
rect 324374 103128 324379 103184
rect 321908 103126 324379 103128
rect 252461 103123 252527 103126
rect 324313 103123 324379 103126
rect 307477 103050 307543 103053
rect 307477 103048 310132 103050
rect 307477 102992 307482 103048
rect 307538 102992 310132 103048
rect 307477 102990 310132 102992
rect 307477 102987 307543 102990
rect 216029 102914 216095 102917
rect 216029 102912 217212 102914
rect 216029 102856 216034 102912
rect 216090 102856 217212 102912
rect 216029 102854 217212 102856
rect 216029 102851 216095 102854
rect 251173 102778 251239 102781
rect 248860 102776 251239 102778
rect 248860 102720 251178 102776
rect 251234 102720 251239 102776
rect 248860 102718 251239 102720
rect 251173 102715 251239 102718
rect 306925 102506 306991 102509
rect 306925 102504 310132 102506
rect 306925 102448 306930 102504
rect 306986 102448 310132 102504
rect 306925 102446 310132 102448
rect 321908 102446 325710 102506
rect 306925 102443 306991 102446
rect 66069 102370 66135 102373
rect 68142 102370 68816 102376
rect 66069 102368 68816 102370
rect 66069 102312 66074 102368
rect 66130 102316 68816 102368
rect 66130 102312 68202 102316
rect 66069 102310 68202 102312
rect 66069 102307 66135 102310
rect 325650 102370 325710 102446
rect 334014 102370 334020 102372
rect 325650 102310 334020 102370
rect 334014 102308 334020 102310
rect 334084 102308 334090 102372
rect 213913 102234 213979 102237
rect 251541 102234 251607 102237
rect 213913 102232 217212 102234
rect 213913 102176 213918 102232
rect 213974 102176 217212 102232
rect 213913 102174 217212 102176
rect 248860 102232 251607 102234
rect 248860 102176 251546 102232
rect 251602 102176 251607 102232
rect 248860 102174 251607 102176
rect 213913 102171 213979 102174
rect 251541 102171 251607 102174
rect 307569 102098 307635 102101
rect 307569 102096 310132 102098
rect 307569 102040 307574 102096
rect 307630 102040 310132 102096
rect 307569 102038 310132 102040
rect 307569 102035 307635 102038
rect 252461 101826 252527 101829
rect 248860 101824 252527 101826
rect 248860 101768 252466 101824
rect 252522 101768 252527 101824
rect 248860 101766 252527 101768
rect 252461 101763 252527 101766
rect 307477 101690 307543 101693
rect 307477 101688 310132 101690
rect 307477 101632 307482 101688
rect 307538 101632 310132 101688
rect 307477 101630 310132 101632
rect 307477 101627 307543 101630
rect 214005 101554 214071 101557
rect 214005 101552 217212 101554
rect 214005 101496 214010 101552
rect 214066 101496 217212 101552
rect 214005 101494 217212 101496
rect 214005 101491 214071 101494
rect 252369 101418 252435 101421
rect 248860 101416 252435 101418
rect 248860 101360 252374 101416
rect 252430 101360 252435 101416
rect 248860 101358 252435 101360
rect 252369 101355 252435 101358
rect 305678 101220 305684 101284
rect 305748 101282 305754 101284
rect 305748 101222 310132 101282
rect 305748 101220 305754 101222
rect 213913 101010 213979 101013
rect 321878 101010 321938 101660
rect 332542 101010 332548 101012
rect 213913 101008 217212 101010
rect 213913 100952 213918 101008
rect 213974 100952 217212 101008
rect 213913 100950 217212 100952
rect 321878 100950 332548 101010
rect 213913 100947 213979 100950
rect 332542 100948 332548 100950
rect 332612 100948 332618 101012
rect 252093 100874 252159 100877
rect 248860 100872 252159 100874
rect 248860 100816 252098 100872
rect 252154 100816 252159 100872
rect 248860 100814 252159 100816
rect 252093 100811 252159 100814
rect 307661 100874 307727 100877
rect 324589 100874 324655 100877
rect 307661 100872 310132 100874
rect 307661 100816 307666 100872
rect 307722 100816 310132 100872
rect 307661 100814 310132 100816
rect 321908 100872 324655 100874
rect 321908 100816 324594 100872
rect 324650 100816 324655 100872
rect 321908 100814 324655 100816
rect 307661 100811 307727 100814
rect 324589 100811 324655 100814
rect 67265 100738 67331 100741
rect 68142 100738 68816 100744
rect 67265 100736 68816 100738
rect 67265 100680 67270 100736
rect 67326 100684 68816 100736
rect 67326 100680 68202 100684
rect 67265 100678 68202 100680
rect 67265 100675 67331 100678
rect -960 97610 480 97700
rect 2773 97610 2839 97613
rect -960 97608 2839 97610
rect -960 97552 2778 97608
rect 2834 97552 2839 97608
rect -960 97550 2839 97552
rect -960 97460 480 97550
rect 2773 97547 2839 97550
rect 252461 100466 252527 100469
rect 248860 100464 252527 100466
rect 248860 100408 252466 100464
rect 252522 100408 252527 100464
rect 248860 100406 252527 100408
rect 252461 100403 252527 100406
rect 307477 100466 307543 100469
rect 307477 100464 310132 100466
rect 307477 100408 307482 100464
rect 307538 100408 310132 100464
rect 307477 100406 310132 100408
rect 307477 100403 307543 100406
rect 214005 100330 214071 100333
rect 214005 100328 217212 100330
rect 214005 100272 214010 100328
rect 214066 100272 217212 100328
rect 214005 100270 217212 100272
rect 214005 100267 214071 100270
rect 324497 100194 324563 100197
rect 321908 100192 324563 100194
rect 321908 100136 324502 100192
rect 324558 100136 324563 100192
rect 321908 100134 324563 100136
rect 324497 100131 324563 100134
rect 307661 100058 307727 100061
rect 307661 100056 310132 100058
rect 307661 100000 307666 100056
rect 307722 100000 310132 100056
rect 307661 99998 310132 100000
rect 307661 99995 307727 99998
rect 251173 99922 251239 99925
rect 248860 99920 251239 99922
rect 248860 99864 251178 99920
rect 251234 99864 251239 99920
rect 248860 99862 251239 99864
rect 251173 99859 251239 99862
rect 213913 99650 213979 99653
rect 213913 99648 217212 99650
rect 213913 99592 213918 99648
rect 213974 99592 217212 99648
rect 213913 99590 217212 99592
rect 213913 99587 213979 99590
rect 299974 99588 299980 99652
rect 300044 99650 300050 99652
rect 300044 99590 310132 99650
rect 300044 99588 300050 99590
rect 252093 99514 252159 99517
rect 248860 99512 252159 99514
rect 248860 99456 252098 99512
rect 252154 99456 252159 99512
rect 248860 99454 252159 99456
rect 252093 99451 252159 99454
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect 307477 99106 307543 99109
rect 307477 99104 310132 99106
rect 307477 99048 307482 99104
rect 307538 99048 310132 99104
rect 307477 99046 310132 99048
rect 307477 99043 307543 99046
rect 213913 98970 213979 98973
rect 252277 98970 252343 98973
rect 213913 98968 217212 98970
rect 213913 98912 213918 98968
rect 213974 98912 217212 98968
rect 213913 98910 217212 98912
rect 248860 98968 252343 98970
rect 248860 98912 252282 98968
rect 252338 98912 252343 98968
rect 248860 98910 252343 98912
rect 213913 98907 213979 98910
rect 252277 98907 252343 98910
rect 307661 98698 307727 98701
rect 321878 98698 321938 99348
rect 331254 98698 331260 98700
rect 307661 98696 310132 98698
rect 307661 98640 307666 98696
rect 307722 98640 310132 98696
rect 307661 98638 310132 98640
rect 321878 98638 331260 98698
rect 307661 98635 307727 98638
rect 331254 98636 331260 98638
rect 331324 98636 331330 98700
rect 251173 98562 251239 98565
rect 248860 98560 251239 98562
rect 248860 98504 251178 98560
rect 251234 98504 251239 98560
rect 248860 98502 251239 98504
rect 251173 98499 251239 98502
rect 214833 98290 214899 98293
rect 307569 98290 307635 98293
rect 214833 98288 217212 98290
rect 214833 98232 214838 98288
rect 214894 98232 217212 98288
rect 214833 98230 217212 98232
rect 307569 98288 310132 98290
rect 307569 98232 307574 98288
rect 307630 98232 310132 98288
rect 307569 98230 310132 98232
rect 214833 98227 214899 98230
rect 307569 98227 307635 98230
rect 321694 98157 321754 98532
rect 321694 98152 321803 98157
rect 321694 98096 321742 98152
rect 321798 98096 321803 98152
rect 321694 98094 321803 98096
rect 321737 98091 321803 98094
rect 252185 98018 252251 98021
rect 248860 98016 252251 98018
rect 248860 97960 252190 98016
rect 252246 97960 252251 98016
rect 248860 97958 252251 97960
rect 252185 97955 252251 97958
rect 306741 97882 306807 97885
rect 306741 97880 310132 97882
rect 306741 97824 306746 97880
rect 306802 97824 310132 97880
rect 306741 97822 310132 97824
rect 306741 97819 306807 97822
rect 213913 97610 213979 97613
rect 252461 97610 252527 97613
rect 213913 97608 217212 97610
rect 213913 97552 213918 97608
rect 213974 97552 217212 97608
rect 213913 97550 217212 97552
rect 248860 97608 252527 97610
rect 248860 97552 252466 97608
rect 252522 97552 252527 97608
rect 248860 97550 252527 97552
rect 213913 97547 213979 97550
rect 252461 97547 252527 97550
rect 307477 97474 307543 97477
rect 307477 97472 310132 97474
rect 307477 97416 307482 97472
rect 307538 97416 310132 97472
rect 307477 97414 310132 97416
rect 307477 97411 307543 97414
rect 321510 97341 321570 97852
rect 321510 97336 321619 97341
rect 321510 97280 321558 97336
rect 321614 97280 321619 97336
rect 321510 97278 321619 97280
rect 321553 97275 321619 97278
rect 251173 97066 251239 97069
rect 260046 97066 260052 97068
rect 248860 97064 260052 97066
rect 248860 97008 251178 97064
rect 251234 97008 260052 97064
rect 248860 97006 260052 97008
rect 251173 97003 251239 97006
rect 260046 97004 260052 97006
rect 260116 97004 260122 97068
rect 307017 97066 307083 97069
rect 307017 97064 310132 97066
rect 307017 97008 307022 97064
rect 307078 97008 310132 97064
rect 307017 97006 310132 97008
rect 307017 97003 307083 97006
rect 214741 96930 214807 96933
rect 214741 96928 217212 96930
rect 214741 96872 214746 96928
rect 214802 96872 217212 96928
rect 214741 96870 217212 96872
rect 214741 96867 214807 96870
rect 321694 96661 321754 97036
rect 249149 96658 249215 96661
rect 249517 96658 249583 96661
rect 248860 96656 249583 96658
rect 248860 96600 249154 96656
rect 249210 96600 249522 96656
rect 249578 96600 249583 96656
rect 248860 96598 249583 96600
rect 249149 96595 249215 96598
rect 249517 96595 249583 96598
rect 302734 96596 302740 96660
rect 302804 96658 302810 96660
rect 321461 96658 321527 96661
rect 302804 96598 310132 96658
rect 321461 96656 321570 96658
rect 321461 96600 321466 96656
rect 321522 96600 321570 96656
rect 302804 96596 302810 96598
rect 321461 96595 321570 96600
rect 321645 96656 321754 96661
rect 321645 96600 321650 96656
rect 321706 96600 321754 96656
rect 321645 96598 321754 96600
rect 321645 96595 321711 96598
rect 214557 96386 214623 96389
rect 214557 96384 217212 96386
rect 214557 96328 214562 96384
rect 214618 96328 217212 96384
rect 321510 96356 321570 96595
rect 214557 96326 217212 96328
rect 214557 96323 214623 96326
rect 307661 96250 307727 96253
rect 307661 96248 310132 96250
rect 248462 95709 248522 96220
rect 307661 96192 307666 96248
rect 307722 96192 310132 96248
rect 307661 96190 310132 96192
rect 307661 96187 307727 96190
rect 308489 95978 308555 95981
rect 324262 95978 324268 95980
rect 308489 95976 324268 95978
rect 308489 95920 308494 95976
rect 308550 95920 324268 95976
rect 308489 95918 324268 95920
rect 308489 95915 308555 95918
rect 324262 95916 324268 95918
rect 324332 95916 324338 95980
rect 248413 95704 248522 95709
rect 248413 95648 248418 95704
rect 248474 95648 248522 95704
rect 248413 95646 248522 95648
rect 248413 95643 248479 95646
rect 180057 95162 180123 95165
rect 321645 95162 321711 95165
rect 180057 95160 321711 95162
rect 180057 95104 180062 95160
rect 180118 95104 321650 95160
rect 321706 95104 321711 95160
rect 180057 95102 321711 95104
rect 180057 95099 180123 95102
rect 321645 95099 321711 95102
rect 64689 94890 64755 94893
rect 209129 94890 209195 94893
rect 64689 94888 209195 94890
rect 64689 94832 64694 94888
rect 64750 94832 209134 94888
rect 209190 94832 209195 94888
rect 64689 94830 209195 94832
rect 64689 94827 64755 94830
rect 209129 94827 209195 94830
rect 105445 94756 105511 94757
rect 117957 94756 118023 94757
rect 105384 94692 105390 94756
rect 105454 94754 105511 94756
rect 105454 94752 105546 94754
rect 105506 94696 105546 94752
rect 105454 94694 105546 94696
rect 105454 94692 105511 94694
rect 106222 94692 106228 94756
rect 106292 94754 106298 94756
rect 106608 94754 106614 94756
rect 106292 94694 106614 94754
rect 106292 94692 106298 94694
rect 106608 94692 106614 94694
rect 106678 94692 106684 94756
rect 117896 94692 117902 94756
rect 117966 94754 118023 94756
rect 119521 94756 119587 94757
rect 129365 94756 129431 94757
rect 119521 94754 119534 94756
rect 117966 94752 118058 94754
rect 118018 94696 118058 94752
rect 117966 94694 118058 94696
rect 119442 94752 119534 94754
rect 119442 94696 119526 94752
rect 119442 94694 119534 94696
rect 117966 94692 118023 94694
rect 105445 94691 105511 94692
rect 117957 94691 118023 94692
rect 119521 94692 119534 94694
rect 119598 94692 119604 94756
rect 129320 94692 129326 94756
rect 129390 94754 129431 94756
rect 134333 94756 134399 94757
rect 134333 94754 134358 94756
rect 129390 94752 129482 94754
rect 129426 94696 129482 94752
rect 129390 94694 129482 94696
rect 134266 94752 134358 94754
rect 134266 94696 134338 94752
rect 134266 94694 134358 94696
rect 129390 94692 129431 94694
rect 119521 94691 119587 94692
rect 129365 94691 129431 94692
rect 134333 94692 134358 94694
rect 134422 94692 134428 94756
rect 151302 94692 151308 94756
rect 151372 94754 151378 94756
rect 151624 94754 151630 94756
rect 151372 94694 151630 94754
rect 151372 94692 151378 94694
rect 151624 94692 151630 94694
rect 151694 94692 151700 94756
rect 134333 94691 134399 94692
rect 67633 93802 67699 93805
rect 214414 93802 214420 93804
rect 67633 93800 214420 93802
rect 67633 93744 67638 93800
rect 67694 93744 214420 93800
rect 67633 93742 214420 93744
rect 67633 93739 67699 93742
rect 214414 93740 214420 93742
rect 214484 93740 214490 93804
rect 130745 93668 130811 93669
rect 151721 93668 151787 93669
rect 130694 93666 130700 93668
rect 130654 93606 130700 93666
rect 130764 93664 130811 93668
rect 151670 93666 151676 93668
rect 130806 93608 130811 93664
rect 130694 93604 130700 93606
rect 130764 93604 130811 93608
rect 151630 93606 151676 93666
rect 151740 93664 151787 93668
rect 151782 93608 151787 93664
rect 151670 93604 151676 93606
rect 151740 93604 151787 93608
rect 130745 93603 130811 93604
rect 151721 93603 151787 93604
rect 110689 93532 110755 93533
rect 115841 93532 115907 93533
rect 110638 93530 110644 93532
rect 110598 93470 110644 93530
rect 110708 93528 110755 93532
rect 115790 93530 115796 93532
rect 110750 93472 110755 93528
rect 110638 93468 110644 93470
rect 110708 93468 110755 93472
rect 115750 93470 115796 93530
rect 115860 93528 115907 93532
rect 115902 93472 115907 93528
rect 115790 93468 115796 93470
rect 115860 93468 115907 93472
rect 110689 93467 110755 93468
rect 115841 93467 115907 93468
rect 110321 93260 110387 93261
rect 128169 93260 128235 93261
rect 110270 93258 110276 93260
rect 110230 93198 110276 93258
rect 110340 93256 110387 93260
rect 128118 93258 128124 93260
rect 110382 93200 110387 93256
rect 110270 93196 110276 93198
rect 110340 93196 110387 93200
rect 128078 93198 128124 93258
rect 128188 93256 128235 93260
rect 128230 93200 128235 93256
rect 128118 93196 128124 93198
rect 128188 93196 128235 93200
rect 110321 93195 110387 93196
rect 128169 93195 128235 93196
rect 85665 92444 85731 92445
rect 85614 92442 85620 92444
rect 85574 92382 85620 92442
rect 85684 92440 85731 92444
rect 85726 92384 85731 92440
rect 85614 92380 85620 92382
rect 85684 92380 85731 92384
rect 91318 92380 91324 92444
rect 91388 92442 91394 92444
rect 91645 92442 91711 92445
rect 107745 92444 107811 92445
rect 114185 92444 114251 92445
rect 115473 92444 115539 92445
rect 116761 92444 116827 92445
rect 119705 92444 119771 92445
rect 107694 92442 107700 92444
rect 91388 92440 91711 92442
rect 91388 92384 91650 92440
rect 91706 92384 91711 92440
rect 91388 92382 91711 92384
rect 107654 92382 107700 92442
rect 107764 92440 107811 92444
rect 114134 92442 114140 92444
rect 107806 92384 107811 92440
rect 91388 92380 91394 92382
rect 85665 92379 85731 92380
rect 91645 92379 91711 92382
rect 107694 92380 107700 92382
rect 107764 92380 107811 92384
rect 114094 92382 114140 92442
rect 114204 92440 114251 92444
rect 115422 92442 115428 92444
rect 114246 92384 114251 92440
rect 114134 92380 114140 92382
rect 114204 92380 114251 92384
rect 115382 92382 115428 92442
rect 115492 92440 115539 92444
rect 116710 92442 116716 92444
rect 115534 92384 115539 92440
rect 115422 92380 115428 92382
rect 115492 92380 115539 92384
rect 116670 92382 116716 92442
rect 116780 92440 116827 92444
rect 119654 92442 119660 92444
rect 116822 92384 116827 92440
rect 116710 92380 116716 92382
rect 116780 92380 116827 92384
rect 119614 92382 119660 92442
rect 119724 92440 119771 92444
rect 119766 92384 119771 92440
rect 119654 92380 119660 92382
rect 119724 92380 119771 92384
rect 122046 92380 122052 92444
rect 122116 92442 122122 92444
rect 122465 92442 122531 92445
rect 125777 92444 125843 92445
rect 151537 92444 151603 92445
rect 152089 92444 152155 92445
rect 125726 92442 125732 92444
rect 122116 92440 122531 92442
rect 122116 92384 122470 92440
rect 122526 92384 122531 92440
rect 122116 92382 122531 92384
rect 125686 92382 125732 92442
rect 125796 92440 125843 92444
rect 151486 92442 151492 92444
rect 125838 92384 125843 92440
rect 122116 92380 122122 92382
rect 107745 92379 107811 92380
rect 114185 92379 114251 92380
rect 115473 92379 115539 92380
rect 116761 92379 116827 92380
rect 119705 92379 119771 92380
rect 122465 92379 122531 92382
rect 125726 92380 125732 92382
rect 125796 92380 125843 92384
rect 151446 92382 151492 92442
rect 151556 92440 151603 92444
rect 152038 92442 152044 92444
rect 151598 92384 151603 92440
rect 151486 92380 151492 92382
rect 151556 92380 151603 92384
rect 151998 92382 152044 92442
rect 152108 92440 152155 92444
rect 152150 92384 152155 92440
rect 152038 92380 152044 92382
rect 152108 92380 152155 92384
rect 125777 92379 125843 92380
rect 151537 92379 151603 92380
rect 152089 92379 152155 92380
rect 106038 92244 106044 92308
rect 106108 92306 106114 92308
rect 180149 92306 180215 92309
rect 106108 92304 180215 92306
rect 106108 92248 180154 92304
rect 180210 92248 180215 92304
rect 106108 92246 180215 92248
rect 106108 92244 106114 92246
rect 180149 92243 180215 92246
rect 125358 92108 125364 92172
rect 125428 92170 125434 92172
rect 125501 92170 125567 92173
rect 125428 92168 125567 92170
rect 125428 92112 125506 92168
rect 125562 92112 125567 92168
rect 125428 92110 125567 92112
rect 125428 92108 125434 92110
rect 125501 92107 125567 92110
rect 151302 92108 151308 92172
rect 151372 92170 151378 92172
rect 151445 92170 151511 92173
rect 151372 92168 151511 92170
rect 151372 92112 151450 92168
rect 151506 92112 151511 92168
rect 151372 92110 151511 92112
rect 151372 92108 151378 92110
rect 151445 92107 151511 92110
rect 88926 91700 88932 91764
rect 88996 91762 89002 91764
rect 89345 91762 89411 91765
rect 88996 91760 89411 91762
rect 88996 91704 89350 91760
rect 89406 91704 89411 91760
rect 88996 91702 89411 91704
rect 88996 91700 89002 91702
rect 89345 91699 89411 91702
rect 90214 91700 90220 91764
rect 90284 91762 90290 91764
rect 90541 91762 90607 91765
rect 90284 91760 90607 91762
rect 90284 91704 90546 91760
rect 90602 91704 90607 91760
rect 90284 91702 90607 91704
rect 90284 91700 90290 91702
rect 90541 91699 90607 91702
rect 99598 91700 99604 91764
rect 99668 91762 99674 91764
rect 99741 91762 99807 91765
rect 117129 91764 117195 91765
rect 117078 91762 117084 91764
rect 99668 91760 99807 91762
rect 99668 91704 99746 91760
rect 99802 91704 99807 91760
rect 99668 91702 99807 91704
rect 117038 91702 117084 91762
rect 117148 91760 117195 91764
rect 117190 91704 117195 91760
rect 99668 91700 99674 91702
rect 99741 91699 99807 91702
rect 117078 91700 117084 91702
rect 117148 91700 117195 91704
rect 117129 91699 117195 91700
rect 102910 91564 102916 91628
rect 102980 91626 102986 91628
rect 103145 91626 103211 91629
rect 102980 91624 103211 91626
rect 102980 91568 103150 91624
rect 103206 91568 103211 91624
rect 102980 91566 103211 91568
rect 102980 91564 102986 91566
rect 103145 91563 103211 91566
rect 108062 91564 108068 91628
rect 108132 91626 108138 91628
rect 211889 91626 211955 91629
rect 108132 91624 211955 91626
rect 108132 91568 211894 91624
rect 211950 91568 211955 91624
rect 108132 91566 211955 91568
rect 108132 91564 108138 91566
rect 211889 91563 211955 91566
rect 98126 91428 98132 91492
rect 98196 91490 98202 91492
rect 99281 91490 99347 91493
rect 98196 91488 99347 91490
rect 98196 91432 99286 91488
rect 99342 91432 99347 91488
rect 98196 91430 99347 91432
rect 98196 91428 98202 91430
rect 99281 91427 99347 91430
rect 101806 91428 101812 91492
rect 101876 91490 101882 91492
rect 102041 91490 102107 91493
rect 122833 91492 122899 91493
rect 101876 91488 102107 91490
rect 101876 91432 102046 91488
rect 102102 91432 102107 91488
rect 101876 91430 102107 91432
rect 101876 91428 101882 91430
rect 102041 91427 102107 91430
rect 122782 91428 122788 91492
rect 122852 91490 122899 91492
rect 122852 91488 122944 91490
rect 122894 91432 122944 91488
rect 122852 91430 122944 91432
rect 122852 91428 122899 91430
rect 135662 91428 135668 91492
rect 135732 91490 135738 91492
rect 136449 91490 136515 91493
rect 135732 91488 136515 91490
rect 135732 91432 136454 91488
rect 136510 91432 136515 91488
rect 135732 91430 136515 91432
rect 135732 91428 135738 91430
rect 122833 91427 122899 91428
rect 136449 91427 136515 91430
rect 93894 91292 93900 91356
rect 93964 91354 93970 91356
rect 95049 91354 95115 91357
rect 93964 91352 95115 91354
rect 93964 91296 95054 91352
rect 95110 91296 95115 91352
rect 93964 91294 95115 91296
rect 93964 91292 93970 91294
rect 95049 91291 95115 91294
rect 97022 91292 97028 91356
rect 97092 91354 97098 91356
rect 97809 91354 97875 91357
rect 97092 91352 97875 91354
rect 97092 91296 97814 91352
rect 97870 91296 97875 91352
rect 97092 91294 97875 91296
rect 97092 91292 97098 91294
rect 97809 91291 97875 91294
rect 98494 91292 98500 91356
rect 98564 91354 98570 91356
rect 99097 91354 99163 91357
rect 98564 91352 99163 91354
rect 98564 91296 99102 91352
rect 99158 91296 99163 91352
rect 98564 91294 99163 91296
rect 98564 91292 98570 91294
rect 99097 91291 99163 91294
rect 101622 91292 101628 91356
rect 101692 91354 101698 91356
rect 101857 91354 101923 91357
rect 101692 91352 101923 91354
rect 101692 91296 101862 91352
rect 101918 91296 101923 91352
rect 101692 91294 101923 91296
rect 101692 91292 101698 91294
rect 101857 91291 101923 91294
rect 106222 91292 106228 91356
rect 106292 91354 106298 91356
rect 107561 91354 107627 91357
rect 106292 91352 107627 91354
rect 106292 91296 107566 91352
rect 107622 91296 107627 91352
rect 106292 91294 107627 91296
rect 106292 91292 106298 91294
rect 107561 91291 107627 91294
rect 120206 91292 120212 91356
rect 120276 91354 120282 91356
rect 121269 91354 121335 91357
rect 120276 91352 121335 91354
rect 120276 91296 121274 91352
rect 121330 91296 121335 91352
rect 120276 91294 121335 91296
rect 120276 91292 120282 91294
rect 121269 91291 121335 91294
rect 74758 91156 74764 91220
rect 74828 91218 74834 91220
rect 75361 91218 75427 91221
rect 74828 91216 75427 91218
rect 74828 91160 75366 91216
rect 75422 91160 75427 91216
rect 74828 91158 75427 91160
rect 74828 91156 74834 91158
rect 75361 91155 75427 91158
rect 84326 91156 84332 91220
rect 84396 91218 84402 91220
rect 85481 91218 85547 91221
rect 84396 91216 85547 91218
rect 84396 91160 85486 91216
rect 85542 91160 85547 91216
rect 84396 91158 85547 91160
rect 84396 91156 84402 91158
rect 85481 91155 85547 91158
rect 86718 91156 86724 91220
rect 86788 91218 86794 91220
rect 86861 91218 86927 91221
rect 88057 91220 88123 91221
rect 88006 91218 88012 91220
rect 86788 91216 86927 91218
rect 86788 91160 86866 91216
rect 86922 91160 86927 91216
rect 86788 91158 86927 91160
rect 87966 91158 88012 91218
rect 88076 91216 88123 91220
rect 88118 91160 88123 91216
rect 86788 91156 86794 91158
rect 86861 91155 86927 91158
rect 88006 91156 88012 91158
rect 88076 91156 88123 91160
rect 92606 91156 92612 91220
rect 92676 91218 92682 91220
rect 93761 91218 93827 91221
rect 92676 91216 93827 91218
rect 92676 91160 93766 91216
rect 93822 91160 93827 91216
rect 92676 91158 93827 91160
rect 92676 91156 92682 91158
rect 88057 91155 88123 91156
rect 93761 91155 93827 91158
rect 94998 91156 95004 91220
rect 95068 91218 95074 91220
rect 95141 91218 95207 91221
rect 95068 91216 95207 91218
rect 95068 91160 95146 91216
rect 95202 91160 95207 91216
rect 95068 91158 95207 91160
rect 95068 91156 95074 91158
rect 95141 91155 95207 91158
rect 96102 91156 96108 91220
rect 96172 91218 96178 91220
rect 96521 91218 96587 91221
rect 96172 91216 96587 91218
rect 96172 91160 96526 91216
rect 96582 91160 96587 91216
rect 96172 91158 96587 91160
rect 96172 91156 96178 91158
rect 96521 91155 96587 91158
rect 97206 91156 97212 91220
rect 97276 91218 97282 91220
rect 97901 91218 97967 91221
rect 99189 91220 99255 91221
rect 100569 91220 100635 91221
rect 99189 91218 99236 91220
rect 97276 91216 97967 91218
rect 97276 91160 97906 91216
rect 97962 91160 97967 91216
rect 97276 91158 97967 91160
rect 99144 91216 99236 91218
rect 99144 91160 99194 91216
rect 99144 91158 99236 91160
rect 97276 91156 97282 91158
rect 97901 91155 97967 91158
rect 99189 91156 99236 91158
rect 99300 91156 99306 91220
rect 100518 91218 100524 91220
rect 100478 91158 100524 91218
rect 100588 91216 100635 91220
rect 101949 91220 102015 91221
rect 101949 91218 101996 91220
rect 100630 91160 100635 91216
rect 100518 91156 100524 91158
rect 100588 91156 100635 91160
rect 101904 91216 101996 91218
rect 101904 91160 101954 91216
rect 101904 91158 101996 91160
rect 99189 91155 99255 91156
rect 100569 91155 100635 91156
rect 101949 91156 101996 91158
rect 102060 91156 102066 91220
rect 103278 91156 103284 91220
rect 103348 91218 103354 91220
rect 103421 91218 103487 91221
rect 103348 91216 103487 91218
rect 103348 91160 103426 91216
rect 103482 91160 103487 91216
rect 103348 91158 103487 91160
rect 103348 91156 103354 91158
rect 101949 91155 102015 91156
rect 103421 91155 103487 91158
rect 104198 91156 104204 91220
rect 104268 91218 104274 91220
rect 104341 91218 104407 91221
rect 104617 91220 104683 91221
rect 104566 91218 104572 91220
rect 104268 91216 104407 91218
rect 104268 91160 104346 91216
rect 104402 91160 104407 91216
rect 104268 91158 104407 91160
rect 104526 91158 104572 91218
rect 104636 91216 104683 91220
rect 104678 91160 104683 91216
rect 104268 91156 104274 91158
rect 104341 91155 104407 91158
rect 104566 91156 104572 91158
rect 104636 91156 104683 91160
rect 106590 91156 106596 91220
rect 106660 91218 106666 91220
rect 107469 91218 107535 91221
rect 109217 91220 109283 91221
rect 109166 91218 109172 91220
rect 106660 91216 107535 91218
rect 106660 91160 107474 91216
rect 107530 91160 107535 91216
rect 106660 91158 107535 91160
rect 109126 91158 109172 91218
rect 109236 91216 109283 91220
rect 109278 91160 109283 91216
rect 106660 91156 106666 91158
rect 104617 91155 104683 91156
rect 107469 91155 107535 91158
rect 109166 91156 109172 91158
rect 109236 91156 109283 91160
rect 109534 91156 109540 91220
rect 109604 91218 109610 91220
rect 109769 91218 109835 91221
rect 109604 91216 109835 91218
rect 109604 91160 109774 91216
rect 109830 91160 109835 91216
rect 109604 91158 109835 91160
rect 109604 91156 109610 91158
rect 109217 91155 109283 91156
rect 109769 91155 109835 91158
rect 111190 91156 111196 91220
rect 111260 91218 111266 91220
rect 111609 91218 111675 91221
rect 111977 91220 112043 91221
rect 112345 91220 112411 91221
rect 111926 91218 111932 91220
rect 111260 91216 111675 91218
rect 111260 91160 111614 91216
rect 111670 91160 111675 91216
rect 111260 91158 111675 91160
rect 111886 91158 111932 91218
rect 111996 91216 112043 91220
rect 112294 91218 112300 91220
rect 112038 91160 112043 91216
rect 111260 91156 111266 91158
rect 111609 91155 111675 91158
rect 111926 91156 111932 91158
rect 111996 91156 112043 91160
rect 112254 91158 112300 91218
rect 112364 91216 112411 91220
rect 112406 91160 112411 91216
rect 112294 91156 112300 91158
rect 112364 91156 112411 91160
rect 113766 91156 113772 91220
rect 113836 91218 113842 91220
rect 114461 91218 114527 91221
rect 113836 91216 114527 91218
rect 113836 91160 114466 91216
rect 114522 91160 114527 91216
rect 113836 91158 114527 91160
rect 113836 91156 113842 91158
rect 111977 91155 112043 91156
rect 112345 91155 112411 91156
rect 114461 91155 114527 91158
rect 115054 91156 115060 91220
rect 115124 91218 115130 91220
rect 115289 91218 115355 91221
rect 115124 91216 115355 91218
rect 115124 91160 115294 91216
rect 115350 91160 115355 91216
rect 115124 91158 115355 91160
rect 115124 91156 115130 91158
rect 115289 91155 115355 91158
rect 118182 91156 118188 91220
rect 118252 91218 118258 91220
rect 118601 91218 118667 91221
rect 118252 91216 118667 91218
rect 118252 91160 118606 91216
rect 118662 91160 118667 91216
rect 118252 91158 118667 91160
rect 118252 91156 118258 91158
rect 118601 91155 118667 91158
rect 120574 91156 120580 91220
rect 120644 91218 120650 91220
rect 121361 91218 121427 91221
rect 120644 91216 121427 91218
rect 120644 91160 121366 91216
rect 121422 91160 121427 91216
rect 120644 91158 121427 91160
rect 120644 91156 120650 91158
rect 121361 91155 121427 91158
rect 121678 91156 121684 91220
rect 121748 91218 121754 91220
rect 122741 91218 122807 91221
rect 121748 91216 122807 91218
rect 121748 91160 122746 91216
rect 122802 91160 122807 91216
rect 121748 91158 122807 91160
rect 121748 91156 121754 91158
rect 122741 91155 122807 91158
rect 122966 91156 122972 91220
rect 123036 91218 123042 91220
rect 123569 91218 123635 91221
rect 124121 91220 124187 91221
rect 124070 91218 124076 91220
rect 123036 91216 123635 91218
rect 123036 91160 123574 91216
rect 123630 91160 123635 91216
rect 123036 91158 123635 91160
rect 124030 91158 124076 91218
rect 124140 91216 124187 91220
rect 124182 91160 124187 91216
rect 123036 91156 123042 91158
rect 123569 91155 123635 91158
rect 124070 91156 124076 91158
rect 124140 91156 124187 91160
rect 124438 91156 124444 91220
rect 124508 91218 124514 91220
rect 125409 91218 125475 91221
rect 126513 91220 126579 91221
rect 126462 91218 126468 91220
rect 124508 91216 125475 91218
rect 124508 91160 125414 91216
rect 125470 91160 125475 91216
rect 124508 91158 125475 91160
rect 126422 91158 126468 91218
rect 126532 91216 126579 91220
rect 126574 91160 126579 91216
rect 124508 91156 124514 91158
rect 124121 91155 124187 91156
rect 125409 91155 125475 91158
rect 126462 91156 126468 91158
rect 126532 91156 126579 91160
rect 126646 91156 126652 91220
rect 126716 91218 126722 91220
rect 126881 91218 126947 91221
rect 132033 91220 132099 91221
rect 133137 91220 133203 91221
rect 131982 91218 131988 91220
rect 126716 91216 126947 91218
rect 126716 91160 126886 91216
rect 126942 91160 126947 91216
rect 126716 91158 126947 91160
rect 131942 91158 131988 91218
rect 132052 91216 132099 91220
rect 133086 91218 133092 91220
rect 132094 91160 132099 91216
rect 126716 91156 126722 91158
rect 126513 91155 126579 91156
rect 126881 91155 126947 91158
rect 131982 91156 131988 91158
rect 132052 91156 132099 91160
rect 133046 91158 133092 91218
rect 133156 91216 133203 91220
rect 133198 91160 133203 91216
rect 133086 91156 133092 91158
rect 133156 91156 133203 91160
rect 132033 91155 132099 91156
rect 133137 91155 133203 91156
rect 66161 91082 66227 91085
rect 169150 91082 169156 91084
rect 66161 91080 169156 91082
rect 66161 91024 66166 91080
rect 66222 91024 169156 91080
rect 66161 91022 169156 91024
rect 66161 91019 66227 91022
rect 169150 91020 169156 91022
rect 169220 91020 169226 91084
rect 113214 90884 113220 90948
rect 113284 90946 113290 90948
rect 170438 90946 170444 90948
rect 113284 90886 170444 90946
rect 113284 90884 113290 90886
rect 170438 90884 170444 90886
rect 170508 90884 170514 90948
rect 128169 89722 128235 89725
rect 174537 89722 174603 89725
rect 128169 89720 174603 89722
rect 128169 89664 128174 89720
rect 128230 89664 174542 89720
rect 174598 89664 174603 89720
rect 128169 89662 174603 89664
rect 128169 89659 128235 89662
rect 174537 89659 174603 89662
rect 104617 88226 104683 88229
rect 166390 88226 166396 88228
rect 104617 88224 166396 88226
rect 104617 88168 104622 88224
rect 104678 88168 166396 88224
rect 104617 88166 166396 88168
rect 104617 88163 104683 88166
rect 166390 88164 166396 88166
rect 166460 88164 166466 88228
rect 123569 86866 123635 86869
rect 167494 86866 167500 86868
rect 123569 86864 167500 86866
rect 123569 86808 123574 86864
rect 123630 86808 167500 86864
rect 123569 86806 167500 86808
rect 123569 86803 123635 86806
rect 167494 86804 167500 86806
rect 167564 86804 167570 86868
rect 582833 86186 582899 86189
rect 583520 86186 584960 86276
rect 582833 86184 584960 86186
rect 582833 86128 582838 86184
rect 582894 86128 584960 86184
rect 582833 86126 584960 86128
rect 582833 86123 582899 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 96521 84146 96587 84149
rect 167678 84146 167684 84148
rect 96521 84144 167684 84146
rect 96521 84088 96526 84144
rect 96582 84088 167684 84144
rect 96521 84086 167684 84088
rect 96521 84083 96587 84086
rect 167678 84084 167684 84086
rect 167748 84084 167754 84148
rect 121269 84010 121335 84013
rect 166206 84010 166212 84012
rect 121269 84008 166212 84010
rect 121269 83952 121274 84008
rect 121330 83952 166212 84008
rect 121269 83950 166212 83952
rect 121269 83947 121335 83950
rect 166206 83948 166212 83950
rect 166276 83948 166282 84012
rect 101949 82786 102015 82789
rect 171726 82786 171732 82788
rect 101949 82784 171732 82786
rect 101949 82728 101954 82784
rect 102010 82728 171732 82784
rect 101949 82726 171732 82728
rect 101949 82723 102015 82726
rect 171726 82724 171732 82726
rect 171796 82724 171802 82788
rect 107561 80066 107627 80069
rect 170254 80066 170260 80068
rect 107561 80064 170260 80066
rect 107561 80008 107566 80064
rect 107622 80008 170260 80064
rect 107561 80006 170260 80008
rect 107561 80003 107627 80006
rect 170254 80004 170260 80006
rect 170324 80004 170330 80068
rect 49693 75170 49759 75173
rect 301446 75170 301452 75172
rect 49693 75168 301452 75170
rect 49693 75112 49698 75168
rect 49754 75112 301452 75168
rect 49693 75110 301452 75112
rect 49693 75107 49759 75110
rect 301446 75108 301452 75110
rect 301516 75108 301522 75172
rect 580206 72932 580212 72996
rect 580276 72994 580282 72996
rect 583520 72994 584960 73084
rect 580276 72934 584960 72994
rect 580276 72932 580282 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect -960 71574 674 71634
rect -960 71498 480 71574
rect 614 71498 674 71574
rect -960 71484 674 71498
rect 246 71438 674 71484
rect 246 70954 306 71438
rect 246 70894 6930 70954
rect 6870 70410 6930 70894
rect 62614 70410 62620 70412
rect 6870 70350 62620 70410
rect 62614 70348 62620 70350
rect 62684 70348 62690 70412
rect 34513 69594 34579 69597
rect 297214 69594 297220 69596
rect 34513 69592 297220 69594
rect 34513 69536 34518 69592
rect 34574 69536 297220 69592
rect 34513 69534 297220 69536
rect 34513 69531 34579 69534
rect 297214 69532 297220 69534
rect 297284 69532 297290 69596
rect 28993 65514 29059 65517
rect 305678 65514 305684 65516
rect 28993 65512 305684 65514
rect 28993 65456 28998 65512
rect 29054 65456 305684 65512
rect 28993 65454 305684 65456
rect 28993 65451 29059 65454
rect 305678 65452 305684 65454
rect 305748 65452 305754 65516
rect 59353 64154 59419 64157
rect 304206 64154 304212 64156
rect 59353 64152 304212 64154
rect 59353 64096 59358 64152
rect 59414 64096 304212 64152
rect 59353 64094 304212 64096
rect 59353 64091 59419 64094
rect 304206 64092 304212 64094
rect 304276 64092 304282 64156
rect 2773 61434 2839 61437
rect 302734 61434 302740 61436
rect 2773 61432 302740 61434
rect 2773 61376 2778 61432
rect 2834 61376 302740 61432
rect 2773 61374 302740 61376
rect 2773 61371 2839 61374
rect 302734 61372 302740 61374
rect 302804 61372 302810 61436
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 8293 57218 8359 57221
rect 305494 57218 305500 57220
rect 8293 57216 305500 57218
rect 8293 57160 8298 57216
rect 8354 57160 305500 57216
rect 8293 57158 305500 57160
rect 8293 57155 8359 57158
rect 305494 57156 305500 57158
rect 305564 57156 305570 57220
rect 582465 46338 582531 46341
rect 583520 46338 584960 46428
rect 582465 46336 584960 46338
rect 582465 46280 582470 46336
rect 582526 46280 584960 46336
rect 582465 46278 584960 46280
rect 582465 46275 582531 46278
rect 22093 46202 22159 46205
rect 307150 46202 307156 46204
rect 22093 46200 307156 46202
rect 22093 46144 22098 46200
rect 22154 46144 307156 46200
rect 22093 46142 307156 46144
rect 22093 46139 22159 46142
rect 307150 46140 307156 46142
rect 307220 46140 307226 46204
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 112437 43482 112503 43485
rect 306966 43482 306972 43484
rect 112437 43480 306972 43482
rect 112437 43424 112442 43480
rect 112498 43424 306972 43480
rect 112437 43422 306972 43424
rect 112437 43419 112503 43422
rect 306966 43420 306972 43422
rect 307036 43420 307042 43484
rect 582741 33146 582807 33149
rect 583520 33146 584960 33236
rect 582741 33144 584960 33146
rect 582741 33088 582746 33144
rect 582802 33088 584960 33144
rect 582741 33086 584960 33088
rect 582741 33083 582807 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3233 32466 3299 32469
rect -960 32464 3299 32466
rect -960 32408 3238 32464
rect 3294 32408 3299 32464
rect -960 32406 3299 32408
rect -960 32316 480 32406
rect 3233 32403 3299 32406
rect 11053 22674 11119 22677
rect 299974 22674 299980 22676
rect 11053 22672 299980 22674
rect 11053 22616 11058 22672
rect 11114 22616 299980 22672
rect 11053 22614 299980 22616
rect 11053 22611 11119 22614
rect 299974 22612 299980 22614
rect 300044 22612 300050 22676
rect 582557 19818 582623 19821
rect 583520 19818 584960 19908
rect 582557 19816 584960 19818
rect 582557 19760 582562 19816
rect 582618 19760 584960 19816
rect 582557 19758 584960 19760
rect 582557 19755 582623 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3509 19410 3575 19413
rect -960 19408 3575 19410
rect -960 19352 3514 19408
rect 3570 19352 3575 19408
rect -960 19350 3575 19352
rect -960 19260 480 19350
rect 3509 19347 3575 19350
rect 582373 6626 582439 6629
rect 583520 6626 584960 6716
rect 582373 6624 584960 6626
rect -960 6490 480 6580
rect 582373 6568 582378 6624
rect 582434 6568 584960 6624
rect 582373 6566 584960 6568
rect 582373 6563 582439 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 125869 3362 125935 3365
rect 173934 3362 173940 3364
rect 125869 3360 173940 3362
rect 125869 3304 125874 3360
rect 125930 3304 173940 3360
rect 125869 3302 173940 3304
rect 125869 3299 125935 3302
rect 173934 3300 173940 3302
rect 174004 3300 174010 3364
<< obsm3 >>
rect 68800 171594 164756 174600
rect 68800 171534 164694 171594
rect 68800 129304 164756 171534
rect 68816 129244 164756 129304
rect 68800 128080 164756 129244
rect 68816 128020 164756 128080
rect 68800 126312 164756 128020
rect 68816 126252 164756 126312
rect 68800 125224 164756 126252
rect 68816 125164 164756 125224
rect 68800 123592 164756 125164
rect 68816 123532 164756 123592
rect 68800 122640 164756 123532
rect 68816 122580 164756 122640
rect 68800 120872 164756 122580
rect 68816 120812 164756 120872
rect 68800 111754 164756 120812
rect 68800 111694 164694 111754
rect 68800 110122 164756 111694
rect 68800 110062 164694 110122
rect 68800 108762 164756 110062
rect 68800 108702 164694 108762
rect 68800 102376 164756 108702
rect 68816 102316 164756 102376
rect 68800 100744 164756 102316
rect 68816 100684 164756 100744
rect 68800 95100 164756 100684
<< via3 >>
rect 120580 643180 120644 643244
rect 331260 302228 331324 302292
rect 265020 299508 265084 299572
rect 252508 296788 252572 296852
rect 256740 295428 256804 295492
rect 340828 295292 340892 295356
rect 119660 294068 119724 294132
rect 62620 292572 62684 292636
rect 335676 291892 335740 291956
rect 346164 291212 346228 291276
rect 64644 284412 64708 284476
rect 120028 279652 120092 279716
rect 173940 271900 174004 271964
rect 120028 264148 120092 264212
rect 337332 259524 337396 259588
rect 64460 254084 64524 254148
rect 63356 251364 63420 251428
rect 580212 246196 580276 246260
rect 66116 245652 66180 245716
rect 260972 243476 261036 243540
rect 120580 238580 120644 238644
rect 119660 238444 119724 238508
rect 63356 236540 63420 236604
rect 332548 232460 332612 232524
rect 64460 231100 64524 231164
rect 329788 224164 329852 224228
rect 328500 221444 328564 221508
rect 248644 214508 248708 214572
rect 263732 208932 263796 208996
rect 265204 207572 265268 207636
rect 335676 206212 335740 206276
rect 327028 204852 327092 204916
rect 338252 197916 338316 197980
rect 342300 196556 342364 196620
rect 263548 193836 263612 193900
rect 64644 191796 64708 191860
rect 327212 189620 327276 189684
rect 259500 188260 259564 188324
rect 320220 186900 320284 186964
rect 256924 184316 256988 184380
rect 262260 184180 262324 184244
rect 66116 182820 66180 182884
rect 334020 181324 334084 181388
rect 257844 180100 257908 180164
rect 255268 179964 255332 180028
rect 167500 179420 167564 179484
rect 332732 178740 332796 178804
rect 336780 178604 336844 178668
rect 99420 177516 99484 177580
rect 106044 177516 106108 177580
rect 106964 177516 107028 177580
rect 110644 177576 110708 177580
rect 110644 177520 110694 177576
rect 110694 177520 110708 177576
rect 110644 177516 110708 177520
rect 112116 177576 112180 177580
rect 112116 177520 112166 177576
rect 112166 177520 112180 177576
rect 112116 177516 112180 177520
rect 114140 177516 114204 177580
rect 116900 177516 116964 177580
rect 118372 177516 118436 177580
rect 122972 177516 123036 177580
rect 124444 177516 124508 177580
rect 125732 177516 125796 177580
rect 249380 177516 249444 177580
rect 331444 177244 331508 177308
rect 120764 177108 120828 177172
rect 133092 177168 133156 177172
rect 133092 177112 133142 177168
rect 133142 177112 133156 177168
rect 133092 177108 133156 177112
rect 103284 176972 103348 177036
rect 167684 176972 167748 177036
rect 97028 176836 97092 176900
rect 104572 176836 104636 176900
rect 166212 176836 166276 176900
rect 98316 176700 98380 176764
rect 101996 176760 102060 176764
rect 101996 176704 102046 176760
rect 102046 176704 102060 176760
rect 101996 176700 102060 176704
rect 108068 176760 108132 176764
rect 108068 176704 108118 176760
rect 108118 176704 108132 176760
rect 108068 176700 108132 176704
rect 109540 176700 109604 176764
rect 115796 176760 115860 176764
rect 115796 176704 115846 176760
rect 115846 176704 115860 176760
rect 115796 176700 115860 176704
rect 127020 176760 127084 176764
rect 127020 176704 127070 176760
rect 127070 176704 127084 176760
rect 127020 176700 127084 176704
rect 129412 176760 129476 176764
rect 129412 176704 129462 176760
rect 129462 176704 129476 176760
rect 129412 176700 129476 176704
rect 131988 176760 132052 176764
rect 131988 176704 132038 176760
rect 132038 176704 132052 176760
rect 131988 176700 132052 176704
rect 134380 176700 134444 176764
rect 135668 176760 135732 176764
rect 135668 176704 135718 176760
rect 135718 176704 135732 176760
rect 135668 176700 135732 176704
rect 148180 176760 148244 176764
rect 148180 176704 148230 176760
rect 148230 176704 148244 176760
rect 148180 176700 148244 176704
rect 260052 176700 260116 176764
rect 321324 176700 321388 176764
rect 128124 176428 128188 176492
rect 249748 176020 249812 176084
rect 321508 176156 321572 176220
rect 306972 175612 307036 175676
rect 113220 175476 113284 175540
rect 130700 175536 130764 175540
rect 130700 175480 130750 175536
rect 130750 175480 130764 175536
rect 100708 175400 100772 175404
rect 100708 175344 100758 175400
rect 100758 175344 100772 175400
rect 100708 175340 100772 175344
rect 121868 175400 121932 175404
rect 121868 175344 121918 175400
rect 121918 175344 121932 175400
rect 121868 175340 121932 175344
rect 130700 175476 130764 175480
rect 158852 175536 158916 175540
rect 158852 175480 158902 175536
rect 158902 175480 158916 175536
rect 158852 175476 158916 175480
rect 166396 175340 166460 175404
rect 119398 174992 119462 174996
rect 119398 174936 119434 174992
rect 119434 174936 119462 174992
rect 119398 174932 119462 174936
rect 321508 174388 321572 174452
rect 249380 174252 249444 174316
rect 249748 173708 249812 173772
rect 321324 170988 321388 171052
rect 321324 170308 321388 170372
rect 337332 165684 337396 165748
rect 166396 163100 166460 163164
rect 263732 163372 263796 163436
rect 265204 162012 265268 162076
rect 166212 158884 166276 158948
rect 167684 157388 167748 157452
rect 259500 156300 259564 156364
rect 251956 155212 252020 155276
rect 167500 154532 167564 154596
rect 257844 152900 257908 152964
rect 252508 152628 252572 152692
rect 256924 150180 256988 150244
rect 306972 144060 307036 144124
rect 307708 143788 307772 143852
rect 307708 142700 307772 142764
rect 331444 142700 331508 142764
rect 265020 142428 265084 142492
rect 306420 142428 306484 142492
rect 260972 142292 261036 142356
rect 335676 142156 335740 142220
rect 262260 141748 262324 141812
rect 306420 141340 306484 141404
rect 167500 140796 167564 140860
rect 307708 140796 307772 140860
rect 255268 140388 255332 140452
rect 166212 139436 166276 139500
rect 249196 139436 249260 139500
rect 251772 138620 251836 138684
rect 263548 138076 263612 138140
rect 346164 138076 346228 138140
rect 256740 137532 256804 137596
rect 170444 135492 170508 135556
rect 340828 134132 340892 134196
rect 251956 133724 252020 133788
rect 307708 133044 307772 133108
rect 170260 132500 170324 132564
rect 306972 132636 307036 132700
rect 166396 131140 166460 131204
rect 301452 130596 301516 130660
rect 171732 129780 171796 129844
rect 327212 129372 327276 129436
rect 329788 127060 329852 127124
rect 304212 118220 304276 118284
rect 297220 115228 297284 115292
rect 338252 114548 338316 114612
rect 307156 114004 307220 114068
rect 305500 112644 305564 112708
rect 336780 110468 336844 110532
rect 167684 109108 167748 109172
rect 332732 109516 332796 109580
rect 335676 109108 335740 109172
rect 328500 106388 328564 106452
rect 342300 106252 342364 106316
rect 251772 105028 251836 105092
rect 214420 104892 214484 104956
rect 324268 104756 324332 104820
rect 327028 103940 327092 104004
rect 169156 103532 169220 103596
rect 334020 102308 334084 102372
rect 305684 101220 305748 101284
rect 332548 100948 332612 101012
rect 299980 99588 300044 99652
rect 331260 98636 331324 98700
rect 260052 97004 260116 97068
rect 302740 96596 302804 96660
rect 324268 95916 324332 95980
rect 105390 94752 105454 94756
rect 105390 94696 105450 94752
rect 105450 94696 105454 94752
rect 105390 94692 105454 94696
rect 106228 94692 106292 94756
rect 106614 94692 106678 94756
rect 117902 94752 117966 94756
rect 117902 94696 117962 94752
rect 117962 94696 117966 94752
rect 117902 94692 117966 94696
rect 119534 94752 119598 94756
rect 119534 94696 119582 94752
rect 119582 94696 119598 94752
rect 119534 94692 119598 94696
rect 129326 94752 129390 94756
rect 129326 94696 129370 94752
rect 129370 94696 129390 94752
rect 129326 94692 129390 94696
rect 134358 94752 134422 94756
rect 134358 94696 134394 94752
rect 134394 94696 134422 94752
rect 134358 94692 134422 94696
rect 151308 94692 151372 94756
rect 151630 94692 151694 94756
rect 214420 93740 214484 93804
rect 130700 93664 130764 93668
rect 130700 93608 130750 93664
rect 130750 93608 130764 93664
rect 130700 93604 130764 93608
rect 151676 93664 151740 93668
rect 151676 93608 151726 93664
rect 151726 93608 151740 93664
rect 151676 93604 151740 93608
rect 110644 93528 110708 93532
rect 110644 93472 110694 93528
rect 110694 93472 110708 93528
rect 110644 93468 110708 93472
rect 115796 93528 115860 93532
rect 115796 93472 115846 93528
rect 115846 93472 115860 93528
rect 115796 93468 115860 93472
rect 110276 93256 110340 93260
rect 110276 93200 110326 93256
rect 110326 93200 110340 93256
rect 110276 93196 110340 93200
rect 128124 93256 128188 93260
rect 128124 93200 128174 93256
rect 128174 93200 128188 93256
rect 128124 93196 128188 93200
rect 85620 92440 85684 92444
rect 85620 92384 85670 92440
rect 85670 92384 85684 92440
rect 85620 92380 85684 92384
rect 91324 92380 91388 92444
rect 107700 92440 107764 92444
rect 107700 92384 107750 92440
rect 107750 92384 107764 92440
rect 107700 92380 107764 92384
rect 114140 92440 114204 92444
rect 114140 92384 114190 92440
rect 114190 92384 114204 92440
rect 114140 92380 114204 92384
rect 115428 92440 115492 92444
rect 115428 92384 115478 92440
rect 115478 92384 115492 92440
rect 115428 92380 115492 92384
rect 116716 92440 116780 92444
rect 116716 92384 116766 92440
rect 116766 92384 116780 92440
rect 116716 92380 116780 92384
rect 119660 92440 119724 92444
rect 119660 92384 119710 92440
rect 119710 92384 119724 92440
rect 119660 92380 119724 92384
rect 122052 92380 122116 92444
rect 125732 92440 125796 92444
rect 125732 92384 125782 92440
rect 125782 92384 125796 92440
rect 125732 92380 125796 92384
rect 151492 92440 151556 92444
rect 151492 92384 151542 92440
rect 151542 92384 151556 92440
rect 151492 92380 151556 92384
rect 152044 92440 152108 92444
rect 152044 92384 152094 92440
rect 152094 92384 152108 92440
rect 152044 92380 152108 92384
rect 106044 92244 106108 92308
rect 125364 92108 125428 92172
rect 151308 92108 151372 92172
rect 88932 91700 88996 91764
rect 90220 91700 90284 91764
rect 99604 91700 99668 91764
rect 117084 91760 117148 91764
rect 117084 91704 117134 91760
rect 117134 91704 117148 91760
rect 117084 91700 117148 91704
rect 102916 91564 102980 91628
rect 108068 91564 108132 91628
rect 98132 91428 98196 91492
rect 101812 91428 101876 91492
rect 122788 91488 122852 91492
rect 122788 91432 122838 91488
rect 122838 91432 122852 91488
rect 122788 91428 122852 91432
rect 135668 91428 135732 91492
rect 93900 91292 93964 91356
rect 97028 91292 97092 91356
rect 98500 91292 98564 91356
rect 101628 91292 101692 91356
rect 106228 91292 106292 91356
rect 120212 91292 120276 91356
rect 74764 91156 74828 91220
rect 84332 91156 84396 91220
rect 86724 91156 86788 91220
rect 88012 91216 88076 91220
rect 88012 91160 88062 91216
rect 88062 91160 88076 91216
rect 88012 91156 88076 91160
rect 92612 91156 92676 91220
rect 95004 91156 95068 91220
rect 96108 91156 96172 91220
rect 97212 91156 97276 91220
rect 99236 91216 99300 91220
rect 99236 91160 99250 91216
rect 99250 91160 99300 91216
rect 99236 91156 99300 91160
rect 100524 91216 100588 91220
rect 100524 91160 100574 91216
rect 100574 91160 100588 91216
rect 100524 91156 100588 91160
rect 101996 91216 102060 91220
rect 101996 91160 102010 91216
rect 102010 91160 102060 91216
rect 101996 91156 102060 91160
rect 103284 91156 103348 91220
rect 104204 91156 104268 91220
rect 104572 91216 104636 91220
rect 104572 91160 104622 91216
rect 104622 91160 104636 91216
rect 104572 91156 104636 91160
rect 106596 91156 106660 91220
rect 109172 91216 109236 91220
rect 109172 91160 109222 91216
rect 109222 91160 109236 91216
rect 109172 91156 109236 91160
rect 109540 91156 109604 91220
rect 111196 91156 111260 91220
rect 111932 91216 111996 91220
rect 111932 91160 111982 91216
rect 111982 91160 111996 91216
rect 111932 91156 111996 91160
rect 112300 91216 112364 91220
rect 112300 91160 112350 91216
rect 112350 91160 112364 91216
rect 112300 91156 112364 91160
rect 113772 91156 113836 91220
rect 115060 91156 115124 91220
rect 118188 91156 118252 91220
rect 120580 91156 120644 91220
rect 121684 91156 121748 91220
rect 122972 91156 123036 91220
rect 124076 91216 124140 91220
rect 124076 91160 124126 91216
rect 124126 91160 124140 91216
rect 124076 91156 124140 91160
rect 124444 91156 124508 91220
rect 126468 91216 126532 91220
rect 126468 91160 126518 91216
rect 126518 91160 126532 91216
rect 126468 91156 126532 91160
rect 126652 91156 126716 91220
rect 131988 91216 132052 91220
rect 131988 91160 132038 91216
rect 132038 91160 132052 91216
rect 131988 91156 132052 91160
rect 133092 91216 133156 91220
rect 133092 91160 133142 91216
rect 133142 91160 133156 91216
rect 133092 91156 133156 91160
rect 169156 91020 169220 91084
rect 113220 90884 113284 90948
rect 170444 90884 170508 90948
rect 166396 88164 166460 88228
rect 167500 86804 167564 86868
rect 167684 84084 167748 84148
rect 166212 83948 166276 84012
rect 171732 82724 171796 82788
rect 170260 80004 170324 80068
rect 301452 75108 301516 75172
rect 580212 72932 580276 72996
rect 62620 70348 62684 70412
rect 297220 69532 297284 69596
rect 305684 65452 305748 65516
rect 304212 64092 304276 64156
rect 302740 61372 302804 61436
rect 305500 57156 305564 57220
rect 307156 46140 307220 46204
rect 306972 43420 307036 43484
rect 299980 22612 300044 22676
rect 173940 3300 174004 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 62619 292636 62685 292637
rect 62619 292572 62620 292636
rect 62684 292572 62685 292636
rect 62619 292571 62685 292572
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 60294 205954 60914 241398
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 62622 70413 62682 292571
rect 64643 284476 64709 284477
rect 64643 284412 64644 284476
rect 64708 284412 64709 284476
rect 64643 284411 64709 284412
rect 64459 254148 64525 254149
rect 64459 254084 64460 254148
rect 64524 254084 64525 254148
rect 64459 254083 64525 254084
rect 63355 251428 63421 251429
rect 63355 251364 63356 251428
rect 63420 251364 63421 251428
rect 63355 251363 63421 251364
rect 63358 236605 63418 251363
rect 63355 236604 63421 236605
rect 63355 236540 63356 236604
rect 63420 236540 63421 236604
rect 63355 236539 63421 236540
rect 64462 231165 64522 254083
rect 64459 231164 64525 231165
rect 64459 231100 64460 231164
rect 64524 231100 64525 231164
rect 64459 231099 64525 231100
rect 64646 191861 64706 284411
rect 64794 282454 65414 317898
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 294000 69914 322398
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 294000 74414 326898
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 294000 78914 295398
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 294000 83414 299898
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 294000 87914 304398
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 294000 92414 308898
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 294000 96914 313398
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 294000 101414 317898
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 294000 105914 322398
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 294000 110414 326898
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 294000 114914 295398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 120579 643244 120645 643245
rect 120579 643180 120580 643244
rect 120644 643180 120645 643244
rect 120579 643179 120645 643180
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 294000 119414 299898
rect 119659 294132 119725 294133
rect 119659 294068 119660 294132
rect 119724 294068 119725 294132
rect 119659 294067 119725 294068
rect 119662 287070 119722 294067
rect 119662 287010 120090 287070
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 120030 279717 120090 287010
rect 120027 279716 120093 279717
rect 120027 279652 120028 279716
rect 120092 279652 120093 279716
rect 120027 279651 120093 279652
rect 120027 264212 120093 264213
rect 120027 264148 120028 264212
rect 120092 264148 120093 264212
rect 120027 264147 120093 264148
rect 89568 259954 89888 259986
rect 89568 259718 89610 259954
rect 89846 259718 89888 259954
rect 89568 259634 89888 259718
rect 89568 259398 89610 259634
rect 89846 259398 89888 259634
rect 89568 259366 89888 259398
rect 120030 258090 120090 264147
rect 119662 258030 120090 258090
rect 74208 255454 74528 255486
rect 74208 255218 74250 255454
rect 74486 255218 74528 255454
rect 74208 255134 74528 255218
rect 74208 254898 74250 255134
rect 74486 254898 74528 255134
rect 74208 254866 74528 254898
rect 104928 255454 105248 255486
rect 104928 255218 104970 255454
rect 105206 255218 105248 255454
rect 104928 255134 105248 255218
rect 104928 254898 104970 255134
rect 105206 254898 105248 255134
rect 104928 254866 105248 254898
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 66115 245716 66181 245717
rect 66115 245652 66116 245716
rect 66180 245652 66181 245716
rect 66115 245651 66181 245652
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64643 191860 64709 191861
rect 64643 191796 64644 191860
rect 64708 191796 64709 191860
rect 64643 191795 64709 191796
rect 64794 174454 65414 209898
rect 66118 182885 66178 245651
rect 119662 238509 119722 258030
rect 120582 238645 120642 643179
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 120579 238644 120645 238645
rect 120579 238580 120580 238644
rect 120644 238580 120645 238644
rect 120579 238579 120645 238580
rect 119659 238508 119725 238509
rect 119659 238444 119660 238508
rect 119724 238444 119725 238508
rect 119659 238443 119725 238444
rect 69294 214954 69914 238000
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 66115 182884 66181 182885
rect 66115 182820 66116 182884
rect 66180 182820 66181 182884
rect 66115 182819 66181 182820
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 176600 69914 178398
rect 73794 219454 74414 238000
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 176600 74414 182898
rect 78294 223954 78914 238000
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 176600 78914 187398
rect 82794 228454 83414 238000
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 176600 83414 191898
rect 87294 232954 87914 238000
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 176600 87914 196398
rect 91794 237454 92414 238000
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 176600 92414 200898
rect 105294 214954 105914 238000
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 99419 177580 99485 177581
rect 99419 177516 99420 177580
rect 99484 177516 99485 177580
rect 99419 177515 99485 177516
rect 97027 176900 97093 176901
rect 97027 176836 97028 176900
rect 97092 176836 97093 176900
rect 97027 176835 97093 176836
rect 97030 175130 97090 176835
rect 98315 176764 98381 176765
rect 98315 176700 98316 176764
rect 98380 176700 98381 176764
rect 98315 176699 98381 176700
rect 96960 175070 97090 175130
rect 98318 175130 98378 176699
rect 99422 175130 99482 177515
rect 103283 177036 103349 177037
rect 103283 176972 103284 177036
rect 103348 176972 103349 177036
rect 103283 176971 103349 176972
rect 101995 176764 102061 176765
rect 101995 176700 101996 176764
rect 102060 176700 102061 176764
rect 101995 176699 102061 176700
rect 100707 175404 100773 175405
rect 100707 175340 100708 175404
rect 100772 175340 100773 175404
rect 100707 175339 100773 175340
rect 98318 175070 98380 175130
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 62619 70412 62685 70413
rect 62619 70348 62620 70412
rect 62684 70348 62685 70412
rect 62619 70347 62685 70348
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 66454 65414 101898
rect 96960 174494 97020 175070
rect 98320 174494 98380 175070
rect 99408 175070 99482 175130
rect 100710 175130 100770 175339
rect 101998 175130 102058 176699
rect 100710 175070 100828 175130
rect 99408 174494 99468 175070
rect 100768 174494 100828 175070
rect 101992 175070 102058 175130
rect 103286 175130 103346 176971
rect 104571 176900 104637 176901
rect 104571 176836 104572 176900
rect 104636 176836 104637 176900
rect 104571 176835 104637 176836
rect 104574 175130 104634 176835
rect 105294 176600 105914 178398
rect 109794 219454 110414 238000
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 106043 177580 106109 177581
rect 106043 177516 106044 177580
rect 106108 177516 106109 177580
rect 106043 177515 106109 177516
rect 106963 177580 107029 177581
rect 106963 177516 106964 177580
rect 107028 177516 107029 177580
rect 106963 177515 107029 177516
rect 106046 175130 106106 177515
rect 103286 175070 103412 175130
rect 104574 175070 104636 175130
rect 101992 174494 102052 175070
rect 103352 174494 103412 175070
rect 104576 174494 104636 175070
rect 105664 175070 106106 175130
rect 106966 175130 107026 177515
rect 108067 176764 108133 176765
rect 108067 176700 108068 176764
rect 108132 176700 108133 176764
rect 108067 176699 108133 176700
rect 109539 176764 109605 176765
rect 109539 176700 109540 176764
rect 109604 176700 109605 176764
rect 109539 176699 109605 176700
rect 108070 175130 108130 176699
rect 109542 175130 109602 176699
rect 109794 176600 110414 182898
rect 114294 223954 114914 238000
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 110643 177580 110709 177581
rect 110643 177516 110644 177580
rect 110708 177516 110709 177580
rect 110643 177515 110709 177516
rect 112115 177580 112181 177581
rect 112115 177516 112116 177580
rect 112180 177516 112181 177580
rect 112115 177515 112181 177516
rect 114139 177580 114205 177581
rect 114139 177516 114140 177580
rect 114204 177516 114205 177580
rect 114139 177515 114205 177516
rect 106966 175070 107084 175130
rect 108070 175070 108172 175130
rect 105664 174494 105724 175070
rect 107024 174494 107084 175070
rect 108112 174494 108172 175070
rect 109472 175070 109602 175130
rect 110646 175130 110706 177515
rect 112118 175130 112178 177515
rect 113219 175540 113285 175541
rect 113219 175476 113220 175540
rect 113284 175476 113285 175540
rect 113219 175475 113285 175476
rect 113222 175130 113282 175475
rect 110646 175070 110756 175130
rect 109472 174494 109532 175070
rect 110696 174494 110756 175070
rect 112056 175070 112178 175130
rect 113144 175070 113282 175130
rect 114142 175130 114202 177515
rect 114294 176600 114914 187398
rect 118794 228454 119414 238000
rect 118794 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 119414 228454
rect 118794 228134 119414 228218
rect 118794 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 119414 228134
rect 118794 192454 119414 227898
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 116899 177580 116965 177581
rect 116899 177516 116900 177580
rect 116964 177516 116965 177580
rect 116899 177515 116965 177516
rect 118371 177580 118437 177581
rect 118371 177516 118372 177580
rect 118436 177516 118437 177580
rect 118371 177515 118437 177516
rect 115795 176764 115861 176765
rect 115795 176700 115796 176764
rect 115860 176700 115861 176764
rect 115795 176699 115861 176700
rect 115798 175130 115858 176699
rect 114142 175070 114428 175130
rect 112056 174494 112116 175070
rect 113144 174494 113204 175070
rect 114368 174494 114428 175070
rect 115728 175070 115858 175130
rect 116902 175130 116962 177515
rect 118374 175130 118434 177515
rect 118794 176600 119414 191898
rect 123294 232954 123914 268398
rect 123294 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 123914 232954
rect 123294 232634 123914 232718
rect 123294 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 123914 232634
rect 123294 196954 123914 232398
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 122971 177580 123037 177581
rect 122971 177516 122972 177580
rect 123036 177516 123037 177580
rect 122971 177515 123037 177516
rect 120763 177172 120829 177173
rect 120763 177108 120764 177172
rect 120828 177108 120829 177172
rect 120763 177107 120829 177108
rect 120766 175130 120826 177107
rect 121867 175404 121933 175405
rect 121867 175340 121868 175404
rect 121932 175340 121933 175404
rect 121867 175339 121933 175340
rect 121870 175130 121930 175339
rect 116902 175070 117012 175130
rect 115728 174494 115788 175070
rect 116952 174494 117012 175070
rect 118312 175070 118434 175130
rect 120760 175070 120826 175130
rect 121848 175070 121930 175130
rect 122974 175130 123034 177515
rect 123294 176600 123914 196398
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 124443 177580 124509 177581
rect 124443 177516 124444 177580
rect 124508 177516 124509 177580
rect 124443 177515 124509 177516
rect 125731 177580 125797 177581
rect 125731 177516 125732 177580
rect 125796 177516 125797 177580
rect 125731 177515 125797 177516
rect 124446 175130 124506 177515
rect 125734 175130 125794 177515
rect 127019 176764 127085 176765
rect 127019 176700 127020 176764
rect 127084 176700 127085 176764
rect 127019 176699 127085 176700
rect 127022 175130 127082 176699
rect 127794 176600 128414 200898
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 241954 132914 277398
rect 132294 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 132914 241954
rect 132294 241634 132914 241718
rect 132294 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 132914 241634
rect 132294 205954 132914 241398
rect 132294 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 132914 205954
rect 132294 205634 132914 205718
rect 132294 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 132914 205634
rect 129411 176764 129477 176765
rect 129411 176700 129412 176764
rect 129476 176700 129477 176764
rect 129411 176699 129477 176700
rect 131987 176764 132053 176765
rect 131987 176700 131988 176764
rect 132052 176700 132053 176764
rect 131987 176699 132053 176700
rect 128123 176492 128189 176493
rect 128123 176428 128124 176492
rect 128188 176428 128189 176492
rect 128123 176427 128189 176428
rect 128126 175130 128186 176427
rect 122974 175070 123132 175130
rect 118312 174494 118372 175070
rect 119397 174996 119463 174997
rect 119397 174932 119398 174996
rect 119462 174932 119463 174996
rect 119397 174931 119463 174932
rect 119400 174494 119460 174931
rect 120760 174494 120820 175070
rect 121848 174494 121908 175070
rect 123072 174494 123132 175070
rect 124432 175070 124506 175130
rect 125656 175070 125794 175130
rect 127016 175070 127082 175130
rect 128104 175070 128186 175130
rect 129414 175130 129474 176699
rect 130699 175540 130765 175541
rect 130699 175476 130700 175540
rect 130764 175476 130765 175540
rect 130699 175475 130765 175476
rect 130702 175130 130762 175475
rect 129414 175070 129524 175130
rect 124432 174494 124492 175070
rect 125656 174494 125716 175070
rect 127016 174494 127076 175070
rect 128104 174494 128164 175070
rect 129464 174494 129524 175070
rect 130688 175070 130762 175130
rect 131990 175130 132050 176699
rect 132294 176600 132914 205398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 246454 137414 281898
rect 136794 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 137414 246454
rect 136794 246134 137414 246218
rect 136794 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 137414 246134
rect 136794 210454 137414 245898
rect 136794 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 137414 210454
rect 136794 210134 137414 210218
rect 136794 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 137414 210134
rect 133091 177172 133157 177173
rect 133091 177108 133092 177172
rect 133156 177108 133157 177172
rect 133091 177107 133157 177108
rect 133094 175130 133154 177107
rect 134379 176764 134445 176765
rect 134379 176700 134380 176764
rect 134444 176700 134445 176764
rect 134379 176699 134445 176700
rect 135667 176764 135733 176765
rect 135667 176700 135668 176764
rect 135732 176700 135733 176764
rect 135667 176699 135733 176700
rect 134382 175130 134442 176699
rect 131990 175070 132108 175130
rect 133094 175070 133196 175130
rect 130688 174494 130748 175070
rect 132048 174494 132108 175070
rect 133136 174494 133196 175070
rect 134360 175070 134442 175130
rect 135670 175130 135730 176699
rect 136794 176600 137414 209898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 214954 141914 250398
rect 141294 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 141914 214954
rect 141294 214634 141914 214718
rect 141294 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 141914 214634
rect 141294 178954 141914 214398
rect 141294 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 141914 178954
rect 141294 178634 141914 178718
rect 141294 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 141914 178634
rect 141294 176600 141914 178398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 176600 146414 182898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 223954 150914 259398
rect 150294 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 150914 223954
rect 150294 223634 150914 223718
rect 150294 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 150914 223634
rect 150294 187954 150914 223398
rect 150294 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 150914 187954
rect 150294 187634 150914 187718
rect 150294 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 150914 187634
rect 148179 176764 148245 176765
rect 148179 176700 148180 176764
rect 148244 176700 148245 176764
rect 148179 176699 148245 176700
rect 148182 175130 148242 176699
rect 150294 176600 150914 187398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 228454 155414 263898
rect 154794 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 155414 228454
rect 154794 228134 155414 228218
rect 154794 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 155414 228134
rect 154794 192454 155414 227898
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 154794 176600 155414 191898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 232954 159914 268398
rect 159294 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 159914 232954
rect 159294 232634 159914 232718
rect 159294 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 159914 232634
rect 159294 196954 159914 232398
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 159294 196634 159914 196718
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 159294 176600 159914 196398
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 176600 164414 200898
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 241954 168914 277398
rect 168294 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 168914 241954
rect 168294 241634 168914 241718
rect 168294 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 168914 241634
rect 168294 205954 168914 241398
rect 168294 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 168914 205954
rect 168294 205634 168914 205718
rect 168294 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 168914 205634
rect 167499 179484 167565 179485
rect 167499 179420 167500 179484
rect 167564 179420 167565 179484
rect 167499 179419 167565 179420
rect 166211 176900 166277 176901
rect 166211 176836 166212 176900
rect 166276 176836 166277 176900
rect 166211 176835 166277 176836
rect 158851 175540 158917 175541
rect 158851 175476 158852 175540
rect 158916 175476 158917 175540
rect 158851 175475 158917 175476
rect 158854 175130 158914 175475
rect 135670 175070 135780 175130
rect 148182 175070 148292 175130
rect 134360 174494 134420 175070
rect 135720 174494 135780 175070
rect 148232 174494 148292 175070
rect 158840 175070 158914 175130
rect 158840 174494 158900 175070
rect 166214 158949 166274 176835
rect 166395 175404 166461 175405
rect 166395 175340 166396 175404
rect 166460 175340 166461 175404
rect 166395 175339 166461 175340
rect 166398 163165 166458 175339
rect 166395 163164 166461 163165
rect 166395 163100 166396 163164
rect 166460 163100 166461 163164
rect 166395 163099 166461 163100
rect 166211 158948 166277 158949
rect 166211 158884 166212 158948
rect 166276 158884 166277 158948
rect 166211 158883 166277 158884
rect 167502 154597 167562 179419
rect 167683 177036 167749 177037
rect 167683 176972 167684 177036
rect 167748 176972 167749 177036
rect 167683 176971 167749 176972
rect 167686 157453 167746 176971
rect 168294 169954 168914 205398
rect 168294 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 168914 169954
rect 168294 169634 168914 169718
rect 168294 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 168914 169634
rect 167683 157452 167749 157453
rect 167683 157388 167684 157452
rect 167748 157388 167749 157452
rect 167683 157387 167749 157388
rect 167499 154596 167565 154597
rect 167499 154532 167500 154596
rect 167564 154532 167565 154596
rect 167499 154531 167565 154532
rect 69072 151954 69420 151986
rect 69072 151718 69128 151954
rect 69364 151718 69420 151954
rect 69072 151634 69420 151718
rect 69072 151398 69128 151634
rect 69364 151398 69420 151634
rect 69072 151366 69420 151398
rect 164136 151954 164484 151986
rect 164136 151718 164192 151954
rect 164428 151718 164484 151954
rect 164136 151634 164484 151718
rect 164136 151398 164192 151634
rect 164428 151398 164484 151634
rect 164136 151366 164484 151398
rect 69752 147454 70100 147486
rect 69752 147218 69808 147454
rect 70044 147218 70100 147454
rect 69752 147134 70100 147218
rect 69752 146898 69808 147134
rect 70044 146898 70100 147134
rect 69752 146866 70100 146898
rect 163456 147454 163804 147486
rect 163456 147218 163512 147454
rect 163748 147218 163804 147454
rect 163456 147134 163804 147218
rect 163456 146898 163512 147134
rect 163748 146898 163804 147134
rect 163456 146866 163804 146898
rect 167499 140860 167565 140861
rect 167499 140796 167500 140860
rect 167564 140796 167565 140860
rect 167499 140795 167565 140796
rect 166211 139500 166277 139501
rect 166211 139436 166212 139500
rect 166276 139436 166277 139500
rect 166211 139435 166277 139436
rect 69072 115954 69420 115986
rect 69072 115718 69128 115954
rect 69364 115718 69420 115954
rect 69072 115634 69420 115718
rect 69072 115398 69128 115634
rect 69364 115398 69420 115634
rect 69072 115366 69420 115398
rect 164136 115954 164484 115986
rect 164136 115718 164192 115954
rect 164428 115718 164484 115954
rect 164136 115634 164484 115718
rect 164136 115398 164192 115634
rect 164428 115398 164484 115634
rect 164136 115366 164484 115398
rect 69752 111454 70100 111486
rect 69752 111218 69808 111454
rect 70044 111218 70100 111454
rect 69752 111134 70100 111218
rect 69752 110898 69808 111134
rect 70044 110898 70100 111134
rect 69752 110866 70100 110898
rect 163456 111454 163804 111486
rect 163456 111218 163512 111454
rect 163748 111218 163804 111454
rect 163456 111134 163804 111218
rect 163456 110898 163512 111134
rect 163748 110898 163804 111134
rect 163456 110866 163804 110898
rect 74656 94890 74716 95200
rect 84312 94890 84372 95200
rect 85536 94890 85596 95200
rect 86624 94890 86684 95200
rect 87984 94890 88044 95200
rect 88936 94890 88996 95200
rect 74656 94830 74826 94890
rect 84312 94830 84394 94890
rect 85536 94830 85682 94890
rect 86624 94830 86786 94890
rect 87984 94830 88074 94890
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 70954 69914 93100
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 75454 74414 93100
rect 74766 91221 74826 94830
rect 74763 91220 74829 91221
rect 74763 91156 74764 91220
rect 74828 91156 74829 91220
rect 74763 91155 74829 91156
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 79954 78914 93100
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 84454 83414 93100
rect 84334 91221 84394 94830
rect 85622 92445 85682 94830
rect 85619 92444 85685 92445
rect 85619 92380 85620 92444
rect 85684 92380 85685 92444
rect 85619 92379 85685 92380
rect 86726 91221 86786 94830
rect 84331 91220 84397 91221
rect 84331 91156 84332 91220
rect 84396 91156 84397 91220
rect 84331 91155 84397 91156
rect 86723 91220 86789 91221
rect 86723 91156 86724 91220
rect 86788 91156 86789 91220
rect 86723 91155 86789 91156
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 88954 87914 93100
rect 88014 91221 88074 94830
rect 88934 94830 88996 94890
rect 90160 94890 90220 95200
rect 91384 94890 91444 95200
rect 90160 94830 90282 94890
rect 88934 91765 88994 94830
rect 90222 91765 90282 94830
rect 91326 94830 91444 94890
rect 92472 94890 92532 95200
rect 93832 94890 93892 95200
rect 94920 94890 94980 95200
rect 96008 94890 96068 95200
rect 96688 94890 96748 95200
rect 97096 94890 97156 95200
rect 98048 94890 98108 95200
rect 98456 94890 98516 95200
rect 99136 94890 99196 95200
rect 99544 94890 99604 95200
rect 100632 94890 100692 95200
rect 92472 94830 92674 94890
rect 93832 94830 93962 94890
rect 94920 94830 95066 94890
rect 96008 94830 96170 94890
rect 96688 94830 96906 94890
rect 97096 94830 97274 94890
rect 98048 94830 98194 94890
rect 98456 94830 98562 94890
rect 99136 94830 99298 94890
rect 99544 94830 99666 94890
rect 91326 92445 91386 94830
rect 91323 92444 91389 92445
rect 91323 92380 91324 92444
rect 91388 92380 91389 92444
rect 91323 92379 91389 92380
rect 88931 91764 88997 91765
rect 88931 91700 88932 91764
rect 88996 91700 88997 91764
rect 88931 91699 88997 91700
rect 90219 91764 90285 91765
rect 90219 91700 90220 91764
rect 90284 91700 90285 91764
rect 90219 91699 90285 91700
rect 88011 91220 88077 91221
rect 88011 91156 88012 91220
rect 88076 91156 88077 91220
rect 88011 91155 88077 91156
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 57454 92414 93100
rect 92614 91221 92674 94830
rect 93902 91357 93962 94830
rect 93899 91356 93965 91357
rect 93899 91292 93900 91356
rect 93964 91292 93965 91356
rect 93899 91291 93965 91292
rect 95006 91221 95066 94830
rect 96110 91221 96170 94830
rect 96846 93870 96906 94830
rect 96846 93810 97090 93870
rect 92611 91220 92677 91221
rect 92611 91156 92612 91220
rect 92676 91156 92677 91220
rect 92611 91155 92677 91156
rect 95003 91220 95069 91221
rect 95003 91156 95004 91220
rect 95068 91156 95069 91220
rect 95003 91155 95069 91156
rect 96107 91220 96173 91221
rect 96107 91156 96108 91220
rect 96172 91156 96173 91220
rect 96107 91155 96173 91156
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 61954 96914 93100
rect 97030 91357 97090 93810
rect 97027 91356 97093 91357
rect 97027 91292 97028 91356
rect 97092 91292 97093 91356
rect 97027 91291 97093 91292
rect 97214 91221 97274 94830
rect 98134 91493 98194 94830
rect 98131 91492 98197 91493
rect 98131 91428 98132 91492
rect 98196 91428 98197 91492
rect 98131 91427 98197 91428
rect 98502 91357 98562 94830
rect 98499 91356 98565 91357
rect 98499 91292 98500 91356
rect 98564 91292 98565 91356
rect 98499 91291 98565 91292
rect 99238 91221 99298 94830
rect 99606 91765 99666 94830
rect 100526 94830 100692 94890
rect 100768 94890 100828 95200
rect 101856 94890 101916 95200
rect 100768 94830 101690 94890
rect 99603 91764 99669 91765
rect 99603 91700 99604 91764
rect 99668 91700 99669 91764
rect 99603 91699 99669 91700
rect 100526 91221 100586 94830
rect 97211 91220 97277 91221
rect 97211 91156 97212 91220
rect 97276 91156 97277 91220
rect 97211 91155 97277 91156
rect 99235 91220 99301 91221
rect 99235 91156 99236 91220
rect 99300 91156 99301 91220
rect 99235 91155 99301 91156
rect 100523 91220 100589 91221
rect 100523 91156 100524 91220
rect 100588 91156 100589 91220
rect 100523 91155 100589 91156
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 66454 101414 93100
rect 101630 91357 101690 94830
rect 101814 94830 101916 94890
rect 101992 94890 102052 95200
rect 102944 94890 103004 95200
rect 101992 94830 102058 94890
rect 101814 91493 101874 94830
rect 101811 91492 101877 91493
rect 101811 91428 101812 91492
rect 101876 91428 101877 91492
rect 101811 91427 101877 91428
rect 101627 91356 101693 91357
rect 101627 91292 101628 91356
rect 101692 91292 101693 91356
rect 101627 91291 101693 91292
rect 101998 91221 102058 94830
rect 102918 94830 103004 94890
rect 103216 94890 103276 95200
rect 104304 94890 104364 95200
rect 103216 94830 103346 94890
rect 102918 91629 102978 94830
rect 102915 91628 102981 91629
rect 102915 91564 102916 91628
rect 102980 91564 102981 91628
rect 102915 91563 102981 91564
rect 103286 91221 103346 94830
rect 104206 94830 104364 94890
rect 104440 94890 104500 95200
rect 104440 94830 104634 94890
rect 104206 91221 104266 94830
rect 104574 91221 104634 94830
rect 105392 94757 105452 95200
rect 105664 94890 105724 95200
rect 105664 94830 106106 94890
rect 105389 94756 105455 94757
rect 105389 94692 105390 94756
rect 105454 94692 105455 94756
rect 105389 94691 105455 94692
rect 101995 91220 102061 91221
rect 101995 91156 101996 91220
rect 102060 91156 102061 91220
rect 101995 91155 102061 91156
rect 103283 91220 103349 91221
rect 103283 91156 103284 91220
rect 103348 91156 103349 91220
rect 103283 91155 103349 91156
rect 104203 91220 104269 91221
rect 104203 91156 104204 91220
rect 104268 91156 104269 91220
rect 104203 91155 104269 91156
rect 104571 91220 104637 91221
rect 104571 91156 104572 91220
rect 104636 91156 104637 91220
rect 104571 91155 104637 91156
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 70954 105914 93100
rect 106046 92309 106106 94830
rect 106227 94756 106293 94757
rect 106227 94692 106228 94756
rect 106292 94692 106293 94756
rect 106227 94691 106293 94692
rect 106043 92308 106109 92309
rect 106043 92244 106044 92308
rect 106108 92244 106109 92308
rect 106043 92243 106109 92244
rect 106230 91357 106290 94691
rect 106480 94210 106540 95200
rect 106616 94757 106676 95200
rect 107704 94890 107764 95200
rect 108112 94890 108172 95200
rect 107702 94830 107764 94890
rect 108070 94830 108172 94890
rect 109064 94890 109124 95200
rect 109472 94890 109532 95200
rect 110152 94890 110212 95200
rect 110696 94890 110756 95200
rect 111240 94890 111300 95200
rect 109064 94830 109234 94890
rect 109472 94830 109602 94890
rect 110152 94830 110338 94890
rect 106613 94756 106679 94757
rect 106613 94692 106614 94756
rect 106678 94692 106679 94756
rect 106613 94691 106679 94692
rect 106480 94150 106658 94210
rect 106227 91356 106293 91357
rect 106227 91292 106228 91356
rect 106292 91292 106293 91356
rect 106227 91291 106293 91292
rect 106598 91221 106658 94150
rect 107702 92445 107762 94830
rect 107699 92444 107765 92445
rect 107699 92380 107700 92444
rect 107764 92380 107765 92444
rect 107699 92379 107765 92380
rect 108070 91629 108130 94830
rect 108067 91628 108133 91629
rect 108067 91564 108068 91628
rect 108132 91564 108133 91628
rect 108067 91563 108133 91564
rect 109174 91221 109234 94830
rect 109542 91221 109602 94830
rect 110278 93261 110338 94830
rect 110646 94830 110756 94890
rect 111198 94830 111300 94890
rect 111920 94890 111980 95200
rect 112328 94890 112388 95200
rect 111920 94830 111994 94890
rect 110646 93533 110706 94830
rect 110643 93532 110709 93533
rect 110643 93468 110644 93532
rect 110708 93468 110709 93532
rect 110643 93467 110709 93468
rect 110275 93260 110341 93261
rect 110275 93196 110276 93260
rect 110340 93196 110341 93260
rect 110275 93195 110341 93196
rect 106595 91220 106661 91221
rect 106595 91156 106596 91220
rect 106660 91156 106661 91220
rect 106595 91155 106661 91156
rect 109171 91220 109237 91221
rect 109171 91156 109172 91220
rect 109236 91156 109237 91220
rect 109171 91155 109237 91156
rect 109539 91220 109605 91221
rect 109539 91156 109540 91220
rect 109604 91156 109605 91220
rect 109539 91155 109605 91156
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 75454 110414 93100
rect 111198 91221 111258 94830
rect 111934 91221 111994 94830
rect 112302 94830 112388 94890
rect 113144 94890 113204 95200
rect 113688 94890 113748 95200
rect 114368 94890 114428 95200
rect 113144 94830 113282 94890
rect 113688 94830 113834 94890
rect 112302 91221 112362 94830
rect 111195 91220 111261 91221
rect 111195 91156 111196 91220
rect 111260 91156 111261 91220
rect 111195 91155 111261 91156
rect 111931 91220 111997 91221
rect 111931 91156 111932 91220
rect 111996 91156 111997 91220
rect 111931 91155 111997 91156
rect 112299 91220 112365 91221
rect 112299 91156 112300 91220
rect 112364 91156 112365 91220
rect 112299 91155 112365 91156
rect 113222 90949 113282 94830
rect 113774 91221 113834 94830
rect 114142 94830 114428 94890
rect 114776 94890 114836 95200
rect 115456 94890 115516 95200
rect 115864 94890 115924 95200
rect 114776 94830 115122 94890
rect 114142 92445 114202 94830
rect 114139 92444 114205 92445
rect 114139 92380 114140 92444
rect 114204 92380 114205 92444
rect 114139 92379 114205 92380
rect 113771 91220 113837 91221
rect 113771 91156 113772 91220
rect 113836 91156 113837 91220
rect 113771 91155 113837 91156
rect 113219 90948 113285 90949
rect 113219 90884 113220 90948
rect 113284 90884 113285 90948
rect 113219 90883 113285 90884
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 79954 114914 93100
rect 115062 91221 115122 94830
rect 115430 94830 115516 94890
rect 115798 94830 115924 94890
rect 116680 94890 116740 95200
rect 117088 94890 117148 95200
rect 116680 94830 116778 94890
rect 115430 92445 115490 94830
rect 115798 93533 115858 94830
rect 115795 93532 115861 93533
rect 115795 93468 115796 93532
rect 115860 93468 115861 93532
rect 115795 93467 115861 93468
rect 116718 92445 116778 94830
rect 117086 94830 117148 94890
rect 115427 92444 115493 92445
rect 115427 92380 115428 92444
rect 115492 92380 115493 92444
rect 115427 92379 115493 92380
rect 116715 92444 116781 92445
rect 116715 92380 116716 92444
rect 116780 92380 116781 92444
rect 116715 92379 116781 92380
rect 117086 91765 117146 94830
rect 117904 94757 117964 95200
rect 118176 94890 118236 95200
rect 119400 94890 119460 95200
rect 118176 94830 118250 94890
rect 117901 94756 117967 94757
rect 117901 94692 117902 94756
rect 117966 94692 117967 94756
rect 117901 94691 117967 94692
rect 117083 91764 117149 91765
rect 117083 91700 117084 91764
rect 117148 91700 117149 91764
rect 117083 91699 117149 91700
rect 118190 91221 118250 94830
rect 119294 94830 119460 94890
rect 119294 93870 119354 94830
rect 119536 94757 119596 95200
rect 120216 94890 120276 95200
rect 120624 94890 120684 95200
rect 121712 94890 121772 95200
rect 120214 94830 120276 94890
rect 120582 94830 120684 94890
rect 121686 94830 121772 94890
rect 121984 94890 122044 95200
rect 121984 94830 122114 94890
rect 119533 94756 119599 94757
rect 119533 94692 119534 94756
rect 119598 94692 119599 94756
rect 119533 94691 119599 94692
rect 119294 93810 119722 93870
rect 115059 91220 115125 91221
rect 115059 91156 115060 91220
rect 115124 91156 115125 91220
rect 115059 91155 115125 91156
rect 118187 91220 118253 91221
rect 118187 91156 118188 91220
rect 118252 91156 118253 91220
rect 118187 91155 118253 91156
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114294 43954 114914 79398
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 84454 119414 93100
rect 119662 92445 119722 93810
rect 119659 92444 119725 92445
rect 119659 92380 119660 92444
rect 119724 92380 119725 92444
rect 119659 92379 119725 92380
rect 120214 91357 120274 94830
rect 120211 91356 120277 91357
rect 120211 91292 120212 91356
rect 120276 91292 120277 91356
rect 120211 91291 120277 91292
rect 120582 91221 120642 94830
rect 121686 91221 121746 94830
rect 122054 92445 122114 94830
rect 122800 93870 122860 95200
rect 123208 94890 123268 95200
rect 122606 93810 122860 93870
rect 122974 94830 123268 94890
rect 124024 94890 124084 95200
rect 124432 94890 124492 95200
rect 125384 94890 125444 95200
rect 124024 94830 124138 94890
rect 124432 94830 124506 94890
rect 122051 92444 122117 92445
rect 122051 92380 122052 92444
rect 122116 92380 122117 92444
rect 122051 92379 122117 92380
rect 122606 91490 122666 93810
rect 122787 91492 122853 91493
rect 122787 91490 122788 91492
rect 122606 91430 122788 91490
rect 122787 91428 122788 91430
rect 122852 91428 122853 91492
rect 122787 91427 122853 91428
rect 122974 91221 123034 94830
rect 120579 91220 120645 91221
rect 120579 91156 120580 91220
rect 120644 91156 120645 91220
rect 120579 91155 120645 91156
rect 121683 91220 121749 91221
rect 121683 91156 121684 91220
rect 121748 91156 121749 91220
rect 121683 91155 121749 91156
rect 122971 91220 123037 91221
rect 122971 91156 122972 91220
rect 123036 91156 123037 91220
rect 122971 91155 123037 91156
rect 118794 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 119414 84454
rect 118794 84134 119414 84218
rect 118794 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 119414 84134
rect 118794 48454 119414 83898
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 88954 123914 93100
rect 124078 91221 124138 94830
rect 124446 91221 124506 94830
rect 125366 94830 125444 94890
rect 125656 94890 125716 95200
rect 126472 94890 126532 95200
rect 125656 94830 125794 94890
rect 125366 92173 125426 94830
rect 125734 92445 125794 94830
rect 126470 94830 126532 94890
rect 126608 94890 126668 95200
rect 128104 94890 128164 95200
rect 126608 94830 126714 94890
rect 128104 94830 128186 94890
rect 125731 92444 125797 92445
rect 125731 92380 125732 92444
rect 125796 92380 125797 92444
rect 125731 92379 125797 92380
rect 125363 92172 125429 92173
rect 125363 92108 125364 92172
rect 125428 92108 125429 92172
rect 125363 92107 125429 92108
rect 126470 91221 126530 94830
rect 126654 91221 126714 94830
rect 128126 93261 128186 94830
rect 129328 94757 129388 95200
rect 130688 94890 130748 95200
rect 131912 94890 131972 95200
rect 133136 94890 133196 95200
rect 130688 94830 130762 94890
rect 131912 94830 132050 94890
rect 129325 94756 129391 94757
rect 129325 94692 129326 94756
rect 129390 94692 129391 94756
rect 129325 94691 129391 94692
rect 130702 93669 130762 94830
rect 130699 93668 130765 93669
rect 130699 93604 130700 93668
rect 130764 93604 130765 93668
rect 130699 93603 130765 93604
rect 128123 93260 128189 93261
rect 128123 93196 128124 93260
rect 128188 93196 128189 93260
rect 128123 93195 128189 93196
rect 124075 91220 124141 91221
rect 124075 91156 124076 91220
rect 124140 91156 124141 91220
rect 124075 91155 124141 91156
rect 124443 91220 124509 91221
rect 124443 91156 124444 91220
rect 124508 91156 124509 91220
rect 124443 91155 124509 91156
rect 126467 91220 126533 91221
rect 126467 91156 126468 91220
rect 126532 91156 126533 91220
rect 126467 91155 126533 91156
rect 126651 91220 126717 91221
rect 126651 91156 126652 91220
rect 126716 91156 126717 91220
rect 126651 91155 126717 91156
rect 123294 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 123914 88954
rect 123294 88634 123914 88718
rect 123294 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 123914 88634
rect 123294 52954 123914 88398
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 57454 128414 93100
rect 131990 91221 132050 94830
rect 133094 94830 133196 94890
rect 131987 91220 132053 91221
rect 131987 91156 131988 91220
rect 132052 91156 132053 91220
rect 131987 91155 132053 91156
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 61954 132914 93100
rect 133094 91221 133154 94830
rect 134360 94757 134420 95200
rect 135584 94890 135644 95200
rect 151496 94890 151556 95200
rect 135584 94830 135730 94890
rect 134357 94756 134423 94757
rect 134357 94692 134358 94756
rect 134422 94692 134423 94756
rect 134357 94691 134423 94692
rect 135670 91493 135730 94830
rect 151494 94830 151556 94890
rect 151307 94756 151373 94757
rect 151307 94692 151308 94756
rect 151372 94692 151373 94756
rect 151307 94691 151373 94692
rect 135667 91492 135733 91493
rect 135667 91428 135668 91492
rect 135732 91428 135733 91492
rect 135667 91427 135733 91428
rect 133091 91220 133157 91221
rect 133091 91156 133092 91220
rect 133156 91156 133157 91220
rect 133091 91155 133157 91156
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5146 132914 25398
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 66454 137414 93100
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6106 137414 29898
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 70954 141914 93100
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7066 141914 34398
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 75454 146414 93100
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 79954 150914 93100
rect 151310 92173 151370 94691
rect 151494 92445 151554 94830
rect 151632 94757 151692 95200
rect 151629 94756 151695 94757
rect 151629 94692 151630 94756
rect 151694 94692 151695 94756
rect 151629 94691 151695 94692
rect 151768 94210 151828 95200
rect 151904 94890 151964 95200
rect 151904 94830 152106 94890
rect 151678 94150 151828 94210
rect 151678 93669 151738 94150
rect 151675 93668 151741 93669
rect 151675 93604 151676 93668
rect 151740 93604 151741 93668
rect 151675 93603 151741 93604
rect 152046 92445 152106 94830
rect 151491 92444 151557 92445
rect 151491 92380 151492 92444
rect 151556 92380 151557 92444
rect 151491 92379 151557 92380
rect 152043 92444 152109 92445
rect 152043 92380 152044 92444
rect 152108 92380 152109 92444
rect 152043 92379 152109 92380
rect 151307 92172 151373 92173
rect 151307 92108 151308 92172
rect 151372 92108 151373 92172
rect 151307 92107 151373 92108
rect 150294 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 150914 79954
rect 150294 79634 150914 79718
rect 150294 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 150914 79634
rect 150294 43954 150914 79398
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 84454 155414 93100
rect 154794 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 155414 84454
rect 154794 84134 155414 84218
rect 154794 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 155414 84134
rect 154794 48454 155414 83898
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 88954 159914 93100
rect 159294 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 159914 88954
rect 159294 88634 159914 88718
rect 159294 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 159914 88634
rect 159294 52954 159914 88398
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 57454 164414 93100
rect 166214 84013 166274 139435
rect 166395 131204 166461 131205
rect 166395 131140 166396 131204
rect 166460 131140 166461 131204
rect 166395 131139 166461 131140
rect 166398 88229 166458 131139
rect 166395 88228 166461 88229
rect 166395 88164 166396 88228
rect 166460 88164 166461 88228
rect 166395 88163 166461 88164
rect 167502 86869 167562 140795
rect 168294 133954 168914 169398
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 246454 173414 281898
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 173939 271964 174005 271965
rect 173939 271900 173940 271964
rect 174004 271900 174005 271964
rect 173939 271899 174005 271900
rect 172794 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 173414 246454
rect 172794 246134 173414 246218
rect 172794 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 173414 246134
rect 172794 210454 173414 245898
rect 172794 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 173414 210454
rect 172794 210134 173414 210218
rect 172794 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 173414 210134
rect 172794 174454 173414 209898
rect 172794 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 173414 174454
rect 172794 174134 173414 174218
rect 172794 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 173414 174134
rect 172794 138454 173414 173898
rect 172794 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 173414 138454
rect 172794 138134 173414 138218
rect 172794 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 173414 138134
rect 170443 135556 170509 135557
rect 170443 135492 170444 135556
rect 170508 135492 170509 135556
rect 170443 135491 170509 135492
rect 168294 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 168914 133954
rect 168294 133634 168914 133718
rect 168294 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 168914 133634
rect 167683 109172 167749 109173
rect 167683 109108 167684 109172
rect 167748 109108 167749 109172
rect 167683 109107 167749 109108
rect 167499 86868 167565 86869
rect 167499 86804 167500 86868
rect 167564 86804 167565 86868
rect 167499 86803 167565 86804
rect 167686 84149 167746 109107
rect 168294 97954 168914 133398
rect 170259 132564 170325 132565
rect 170259 132500 170260 132564
rect 170324 132500 170325 132564
rect 170259 132499 170325 132500
rect 169155 103596 169221 103597
rect 169155 103532 169156 103596
rect 169220 103532 169221 103596
rect 169155 103531 169221 103532
rect 168294 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 168914 97954
rect 168294 97634 168914 97718
rect 168294 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 168914 97634
rect 167683 84148 167749 84149
rect 167683 84084 167684 84148
rect 167748 84084 167749 84148
rect 167683 84083 167749 84084
rect 166211 84012 166277 84013
rect 166211 83948 166212 84012
rect 166276 83948 166277 84012
rect 166211 83947 166277 83948
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 61954 168914 97398
rect 169158 91085 169218 103531
rect 169155 91084 169221 91085
rect 169155 91020 169156 91084
rect 169220 91020 169221 91084
rect 169155 91019 169221 91020
rect 170262 80069 170322 132499
rect 170446 90949 170506 135491
rect 171731 129844 171797 129845
rect 171731 129780 171732 129844
rect 171796 129780 171797 129844
rect 171731 129779 171797 129780
rect 170443 90948 170509 90949
rect 170443 90884 170444 90948
rect 170508 90884 170509 90948
rect 170443 90883 170509 90884
rect 171734 82789 171794 129779
rect 172794 102454 173414 137898
rect 172794 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 173414 102454
rect 172794 102134 173414 102218
rect 172794 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 173414 102134
rect 171731 82788 171797 82789
rect 171731 82724 171732 82788
rect 171796 82724 171797 82788
rect 171731 82723 171797 82724
rect 170259 80068 170325 80069
rect 170259 80004 170260 80068
rect 170324 80004 170325 80068
rect 170259 80003 170325 80004
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5146 168914 25398
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 66454 173414 101898
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6106 173414 29898
rect 173942 3365 174002 271899
rect 177294 250954 177914 286398
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 214954 177914 250398
rect 177294 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 177914 214954
rect 177294 214634 177914 214718
rect 177294 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 177914 214634
rect 177294 178954 177914 214398
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 106954 177914 142398
rect 177294 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 177914 106954
rect 177294 106634 177914 106718
rect 177294 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 177914 106634
rect 177294 70954 177914 106398
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 173939 3364 174005 3365
rect 173939 3300 173940 3364
rect 174004 3300 174005 3364
rect 173939 3299 174005 3300
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 259954 186914 295398
rect 186294 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 186914 259954
rect 186294 259634 186914 259718
rect 186294 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 186914 259634
rect 186294 223954 186914 259398
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 187954 186914 223398
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 115954 186914 151398
rect 186294 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 186914 115954
rect 186294 115634 186914 115718
rect 186294 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 186914 115634
rect 186294 79954 186914 115398
rect 186294 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 186914 79954
rect 186294 79634 186914 79718
rect 186294 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 186914 79634
rect 186294 43954 186914 79398
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 190794 264454 191414 299898
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 228454 191414 263898
rect 190794 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 191414 228454
rect 190794 228134 191414 228218
rect 190794 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 191414 228134
rect 190794 192454 191414 227898
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 120454 191414 155898
rect 190794 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 191414 120454
rect 190794 120134 191414 120218
rect 190794 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 191414 120134
rect 190794 84454 191414 119898
rect 190794 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 191414 84454
rect 190794 84134 191414 84218
rect 190794 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 191414 84134
rect 190794 48454 191414 83898
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 195294 232954 195914 268398
rect 195294 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 195914 232954
rect 195294 232634 195914 232718
rect 195294 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 195914 232634
rect 195294 196954 195914 232398
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 241954 204914 277398
rect 204294 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 204914 241954
rect 204294 241634 204914 241718
rect 204294 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 204914 241634
rect 204294 205954 204914 241398
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 246454 209414 281898
rect 208794 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 209414 246454
rect 208794 246134 209414 246218
rect 208794 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 209414 246134
rect 208794 210454 209414 245898
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 214954 213914 250398
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 178000 218414 182898
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 547954 222914 583398
rect 222294 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 222914 547954
rect 222294 547634 222914 547718
rect 222294 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 222914 547634
rect 222294 511954 222914 547398
rect 222294 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 222914 511954
rect 222294 511634 222914 511718
rect 222294 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 222914 511634
rect 222294 475954 222914 511398
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 223954 222914 259398
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 178000 222914 187398
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 552454 227414 587898
rect 226794 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 227414 552454
rect 226794 552134 227414 552218
rect 226794 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 227414 552134
rect 226794 516454 227414 551898
rect 226794 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 227414 516454
rect 226794 516134 227414 516218
rect 226794 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 227414 516134
rect 226794 480454 227414 515898
rect 226794 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 227414 480454
rect 226794 480134 227414 480218
rect 226794 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 227414 480134
rect 226794 444454 227414 479898
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 228454 227414 263898
rect 226794 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 227414 228454
rect 226794 228134 227414 228218
rect 226794 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 227414 228134
rect 226794 192454 227414 227898
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 178000 227414 191898
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 556954 231914 592398
rect 231294 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 231914 556954
rect 231294 556634 231914 556718
rect 231294 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 231914 556634
rect 231294 520954 231914 556398
rect 231294 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 231914 520954
rect 231294 520634 231914 520718
rect 231294 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 231914 520634
rect 231294 484954 231914 520398
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 231294 412954 231914 448398
rect 231294 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 231914 412954
rect 231294 412634 231914 412718
rect 231294 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 231914 412634
rect 231294 376954 231914 412398
rect 231294 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 231914 376954
rect 231294 376634 231914 376718
rect 231294 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 231914 376634
rect 231294 340954 231914 376398
rect 231294 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 231914 340954
rect 231294 340634 231914 340718
rect 231294 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 231914 340634
rect 231294 304954 231914 340398
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 232954 231914 268398
rect 231294 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 231914 232954
rect 231294 232634 231914 232718
rect 231294 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 231914 232634
rect 231294 196954 231914 232398
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 178000 231914 196398
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 178000 236414 200898
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 529954 240914 565398
rect 240294 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 240914 529954
rect 240294 529634 240914 529718
rect 240294 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 240914 529634
rect 240294 493954 240914 529398
rect 240294 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 240914 493954
rect 240294 493634 240914 493718
rect 240294 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 240914 493634
rect 240294 457954 240914 493398
rect 240294 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 240914 457954
rect 240294 457634 240914 457718
rect 240294 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 240914 457634
rect 240294 421954 240914 457398
rect 240294 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 240914 421954
rect 240294 421634 240914 421718
rect 240294 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 240914 421634
rect 240294 385954 240914 421398
rect 240294 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 240914 385954
rect 240294 385634 240914 385718
rect 240294 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 240914 385634
rect 240294 349954 240914 385398
rect 240294 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 240914 349954
rect 240294 349634 240914 349718
rect 240294 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 240914 349634
rect 240294 313954 240914 349398
rect 240294 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 240914 313954
rect 240294 313634 240914 313718
rect 240294 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 240914 313634
rect 240294 277954 240914 313398
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 240294 241954 240914 277398
rect 240294 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 240914 241954
rect 240294 241634 240914 241718
rect 240294 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 240914 241634
rect 240294 205954 240914 241398
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 240294 178000 240914 205398
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 534454 245414 569898
rect 244794 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 245414 534454
rect 244794 534134 245414 534218
rect 244794 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 245414 534134
rect 244794 498454 245414 533898
rect 244794 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 245414 498454
rect 244794 498134 245414 498218
rect 244794 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 245414 498134
rect 244794 462454 245414 497898
rect 244794 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 245414 462454
rect 244794 462134 245414 462218
rect 244794 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 245414 462134
rect 244794 426454 245414 461898
rect 244794 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 245414 426454
rect 244794 426134 245414 426218
rect 244794 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 245414 426134
rect 244794 390454 245414 425898
rect 244794 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 245414 390454
rect 244794 390134 245414 390218
rect 244794 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 245414 390134
rect 244794 354454 245414 389898
rect 244794 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 245414 354454
rect 244794 354134 245414 354218
rect 244794 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 245414 354134
rect 244794 318454 245414 353898
rect 244794 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 245414 318454
rect 244794 318134 245414 318218
rect 244794 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 245414 318134
rect 244794 282454 245414 317898
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 246454 245414 281898
rect 244794 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 245414 246454
rect 244794 246134 245414 246218
rect 244794 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 245414 246134
rect 244794 210454 245414 245898
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 538954 249914 574398
rect 249294 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 249914 538954
rect 249294 538634 249914 538718
rect 249294 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 249914 538634
rect 249294 502954 249914 538398
rect 249294 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 249914 502954
rect 249294 502634 249914 502718
rect 249294 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 249914 502634
rect 249294 466954 249914 502398
rect 249294 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 249914 466954
rect 249294 466634 249914 466718
rect 249294 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 249914 466634
rect 249294 430954 249914 466398
rect 249294 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 249914 430954
rect 249294 430634 249914 430718
rect 249294 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 249914 430634
rect 249294 394954 249914 430398
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 249294 358954 249914 394398
rect 249294 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 249914 358954
rect 249294 358634 249914 358718
rect 249294 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 249914 358634
rect 249294 322954 249914 358398
rect 249294 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 249914 322954
rect 249294 322634 249914 322718
rect 249294 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 249914 322634
rect 249294 286954 249914 322398
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 252507 296852 252573 296853
rect 252507 296788 252508 296852
rect 252572 296788 252573 296852
rect 252507 296787 252573 296788
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 214954 249914 250398
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 248643 214572 248709 214573
rect 248643 214508 248644 214572
rect 248708 214508 248709 214572
rect 248643 214507 248709 214508
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 178000 245414 209898
rect 248646 175810 248706 214507
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 178000 249914 178398
rect 249379 177580 249445 177581
rect 249379 177516 249380 177580
rect 249444 177516 249445 177580
rect 249379 177515 249445 177516
rect 248646 175750 249258 175810
rect 227874 151954 228194 151986
rect 227874 151718 227916 151954
rect 228152 151718 228194 151954
rect 227874 151634 228194 151718
rect 227874 151398 227916 151634
rect 228152 151398 228194 151634
rect 227874 151366 228194 151398
rect 237805 151954 238125 151986
rect 237805 151718 237847 151954
rect 238083 151718 238125 151954
rect 237805 151634 238125 151718
rect 237805 151398 237847 151634
rect 238083 151398 238125 151634
rect 237805 151366 238125 151398
rect 222910 147454 223230 147486
rect 222910 147218 222952 147454
rect 223188 147218 223230 147454
rect 222910 147134 223230 147218
rect 222910 146898 222952 147134
rect 223188 146898 223230 147134
rect 222910 146866 223230 146898
rect 232840 147454 233160 147486
rect 232840 147218 232882 147454
rect 233118 147218 233160 147454
rect 232840 147134 233160 147218
rect 232840 146898 232882 147134
rect 233118 146898 233160 147134
rect 232840 146866 233160 146898
rect 242771 147454 243091 147486
rect 242771 147218 242813 147454
rect 243049 147218 243091 147454
rect 242771 147134 243091 147218
rect 242771 146898 242813 147134
rect 243049 146898 243091 147134
rect 242771 146866 243091 146898
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 249198 139501 249258 175750
rect 249382 174317 249442 177515
rect 249747 176084 249813 176085
rect 249747 176020 249748 176084
rect 249812 176020 249813 176084
rect 249747 176019 249813 176020
rect 249379 174316 249445 174317
rect 249379 174252 249380 174316
rect 249444 174252 249445 174316
rect 249379 174251 249445 174252
rect 249750 173773 249810 176019
rect 249747 173772 249813 173773
rect 249747 173708 249748 173772
rect 249812 173708 249813 173772
rect 249747 173707 249813 173708
rect 251955 155276 252021 155277
rect 251955 155212 251956 155276
rect 252020 155212 252021 155276
rect 251955 155211 252021 155212
rect 249195 139500 249261 139501
rect 249195 139436 249196 139500
rect 249260 139436 249261 139500
rect 249195 139435 249261 139436
rect 251771 138684 251837 138685
rect 251771 138620 251772 138684
rect 251836 138620 251837 138684
rect 251771 138619 251837 138620
rect 227874 115954 228194 115986
rect 227874 115718 227916 115954
rect 228152 115718 228194 115954
rect 227874 115634 228194 115718
rect 227874 115398 227916 115634
rect 228152 115398 228194 115634
rect 227874 115366 228194 115398
rect 237805 115954 238125 115986
rect 237805 115718 237847 115954
rect 238083 115718 238125 115954
rect 237805 115634 238125 115718
rect 237805 115398 237847 115634
rect 238083 115398 238125 115634
rect 237805 115366 238125 115398
rect 222910 111454 223230 111486
rect 222910 111218 222952 111454
rect 223188 111218 223230 111454
rect 222910 111134 223230 111218
rect 222910 110898 222952 111134
rect 223188 110898 223230 111134
rect 222910 110866 223230 110898
rect 232840 111454 233160 111486
rect 232840 111218 232882 111454
rect 233118 111218 233160 111454
rect 232840 111134 233160 111218
rect 232840 110898 232882 111134
rect 233118 110898 233160 111134
rect 232840 110866 233160 110898
rect 242771 111454 243091 111486
rect 242771 111218 242813 111454
rect 243049 111218 243091 111454
rect 242771 111134 243091 111218
rect 242771 110898 242813 111134
rect 243049 110898 243091 111134
rect 242771 110866 243091 110898
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 251774 105093 251834 138619
rect 251958 133789 252018 155211
rect 252510 152693 252570 296787
rect 253794 291454 254414 326898
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 258294 367954 258914 403398
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 258294 331954 258914 367398
rect 258294 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 258914 331954
rect 258294 331634 258914 331718
rect 258294 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 258914 331634
rect 258294 295954 258914 331398
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 256739 295492 256805 295493
rect 256739 295428 256740 295492
rect 256804 295428 256805 295492
rect 256739 295427 256805 295428
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 252507 152692 252573 152693
rect 252507 152628 252508 152692
rect 252572 152628 252573 152692
rect 252507 152627 252573 152628
rect 253794 147454 254414 182898
rect 255267 180028 255333 180029
rect 255267 179964 255268 180028
rect 255332 179964 255333 180028
rect 255267 179963 255333 179964
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 251955 133788 252021 133789
rect 251955 133724 251956 133788
rect 252020 133724 252021 133788
rect 251955 133723 252021 133724
rect 253794 111454 254414 146898
rect 255270 140453 255330 179963
rect 255267 140452 255333 140453
rect 255267 140388 255268 140452
rect 255332 140388 255333 140452
rect 255267 140387 255333 140388
rect 256742 137597 256802 295427
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 223954 258914 259398
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 372454 263414 407898
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 336454 263414 371898
rect 262794 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 263414 336454
rect 262794 336134 263414 336218
rect 262794 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 263414 336134
rect 262794 300454 263414 335898
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 376954 267914 412398
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 340954 267914 376398
rect 267294 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 267914 340954
rect 267294 340634 267914 340718
rect 267294 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 267914 340634
rect 267294 304954 267914 340398
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 265019 299572 265085 299573
rect 265019 299508 265020 299572
rect 265084 299508 265085 299572
rect 265019 299507 265085 299508
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 260971 243540 261037 243541
rect 260971 243476 260972 243540
rect 261036 243476 261037 243540
rect 260971 243475 261037 243476
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 259499 188324 259565 188325
rect 259499 188260 259500 188324
rect 259564 188260 259565 188324
rect 259499 188259 259565 188260
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 256923 184380 256989 184381
rect 256923 184316 256924 184380
rect 256988 184316 256989 184380
rect 256923 184315 256989 184316
rect 256926 150245 256986 184315
rect 257843 180164 257909 180165
rect 257843 180100 257844 180164
rect 257908 180100 257909 180164
rect 257843 180099 257909 180100
rect 257846 152965 257906 180099
rect 257843 152964 257909 152965
rect 257843 152900 257844 152964
rect 257908 152900 257909 152964
rect 257843 152899 257909 152900
rect 258294 151954 258914 187398
rect 259502 156365 259562 188259
rect 260051 176764 260117 176765
rect 260051 176700 260052 176764
rect 260116 176700 260117 176764
rect 260051 176699 260117 176700
rect 259499 156364 259565 156365
rect 259499 156300 259500 156364
rect 259564 156300 259565 156364
rect 259499 156299 259565 156300
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 256923 150244 256989 150245
rect 256923 150180 256924 150244
rect 256988 150180 256989 150244
rect 256923 150179 256989 150180
rect 256739 137596 256805 137597
rect 256739 137532 256740 137596
rect 256804 137532 256805 137596
rect 256739 137531 256805 137532
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 251771 105092 251837 105093
rect 251771 105028 251772 105092
rect 251836 105028 251837 105092
rect 251771 105027 251837 105028
rect 214419 104956 214485 104957
rect 214419 104892 214420 104956
rect 214484 104892 214485 104956
rect 214419 104891 214485 104892
rect 214422 93805 214482 104891
rect 214419 93804 214485 93805
rect 214419 93740 214420 93804
rect 214484 93740 214485 93804
rect 214419 93739 214485 93740
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 75454 218414 94000
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 79954 222914 94000
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 84454 227414 94000
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 88954 231914 94000
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 93454 236414 94000
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 61954 240914 94000
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 66454 245414 94000
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 70954 249914 94000
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 260054 97069 260114 176699
rect 260974 142357 261034 243475
rect 262794 228454 263414 263898
rect 262794 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 263414 228454
rect 262794 228134 263414 228218
rect 262794 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 263414 228134
rect 262794 192454 263414 227898
rect 263731 208996 263797 208997
rect 263731 208932 263732 208996
rect 263796 208932 263797 208996
rect 263731 208931 263797 208932
rect 263547 193900 263613 193901
rect 263547 193836 263548 193900
rect 263612 193836 263613 193900
rect 263547 193835 263613 193836
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262259 184244 262325 184245
rect 262259 184180 262260 184244
rect 262324 184180 262325 184244
rect 262259 184179 262325 184180
rect 260971 142356 261037 142357
rect 260971 142292 260972 142356
rect 261036 142292 261037 142356
rect 260971 142291 261037 142292
rect 262262 141813 262322 184179
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262259 141812 262325 141813
rect 262259 141748 262260 141812
rect 262324 141748 262325 141812
rect 262259 141747 262325 141748
rect 262794 120454 263414 155898
rect 263550 138141 263610 193835
rect 263734 163437 263794 208931
rect 263731 163436 263797 163437
rect 263731 163372 263732 163436
rect 263796 163372 263797 163436
rect 263731 163371 263797 163372
rect 265022 142493 265082 299507
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 232954 267914 268398
rect 267294 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 267914 232954
rect 267294 232634 267914 232718
rect 267294 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 267914 232634
rect 265203 207636 265269 207637
rect 265203 207572 265204 207636
rect 265268 207572 265269 207636
rect 265203 207571 265269 207572
rect 265206 162077 265266 207571
rect 267294 196954 267914 232398
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 265203 162076 265269 162077
rect 265203 162012 265204 162076
rect 265268 162012 265269 162076
rect 265203 162011 265269 162012
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 265019 142492 265085 142493
rect 265019 142428 265020 142492
rect 265084 142428 265085 142492
rect 265019 142427 265085 142428
rect 263547 138140 263613 138141
rect 263547 138076 263548 138140
rect 263612 138076 263613 138140
rect 263547 138075 263613 138076
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 260051 97068 260117 97069
rect 260051 97004 260052 97068
rect 260116 97004 260117 97068
rect 260051 97003 260117 97004
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 529954 276914 565398
rect 276294 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 276914 529954
rect 276294 529634 276914 529718
rect 276294 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 276914 529634
rect 276294 493954 276914 529398
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 349954 276914 385398
rect 276294 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 276914 349954
rect 276294 349634 276914 349718
rect 276294 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 276914 349634
rect 276294 313954 276914 349398
rect 276294 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 276914 313954
rect 276294 313634 276914 313718
rect 276294 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 276914 313634
rect 276294 277954 276914 313398
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 241954 276914 277398
rect 276294 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 276914 241954
rect 276294 241634 276914 241718
rect 276294 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 276914 241634
rect 276294 205954 276914 241398
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 534454 281414 569898
rect 280794 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 281414 534454
rect 280794 534134 281414 534218
rect 280794 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 281414 534134
rect 280794 498454 281414 533898
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 462454 281414 497898
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 354454 281414 389898
rect 280794 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 281414 354454
rect 280794 354134 281414 354218
rect 280794 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 281414 354134
rect 280794 318454 281414 353898
rect 280794 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 281414 318454
rect 280794 318134 281414 318218
rect 280794 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 281414 318134
rect 280794 282454 281414 317898
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 246454 281414 281898
rect 280794 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 281414 246454
rect 280794 246134 281414 246218
rect 280794 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 281414 246134
rect 280794 210454 281414 245898
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 322954 285914 358398
rect 285294 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 285914 322954
rect 285294 322634 285914 322718
rect 285294 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 285914 322634
rect 285294 286954 285914 322398
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 214954 285914 250398
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294294 331954 294914 367398
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 223954 294914 259398
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 552454 299414 587898
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 298794 516454 299414 551898
rect 298794 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 299414 516454
rect 298794 516134 299414 516218
rect 298794 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 299414 516134
rect 298794 480454 299414 515898
rect 298794 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 299414 480454
rect 298794 480134 299414 480218
rect 298794 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 299414 480134
rect 298794 444454 299414 479898
rect 298794 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 299414 444454
rect 298794 444134 299414 444218
rect 298794 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 299414 444134
rect 298794 408454 299414 443898
rect 298794 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 299414 408454
rect 298794 408134 299414 408218
rect 298794 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 299414 408134
rect 298794 372454 299414 407898
rect 298794 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 299414 372454
rect 298794 372134 299414 372218
rect 298794 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 299414 372134
rect 298794 336454 299414 371898
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 298794 300454 299414 335898
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 228454 299414 263898
rect 298794 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 299414 228454
rect 298794 228134 299414 228218
rect 298794 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 299414 228134
rect 298794 192454 299414 227898
rect 298794 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 299414 192454
rect 298794 192134 299414 192218
rect 298794 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 299414 192134
rect 298794 156454 299414 191898
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 556954 303914 592398
rect 303294 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 303914 556954
rect 303294 556634 303914 556718
rect 303294 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 303914 556634
rect 303294 520954 303914 556398
rect 303294 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 303914 520954
rect 303294 520634 303914 520718
rect 303294 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 303914 520634
rect 303294 484954 303914 520398
rect 303294 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 303914 484954
rect 303294 484634 303914 484718
rect 303294 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 303914 484634
rect 303294 448954 303914 484398
rect 303294 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 303914 448954
rect 303294 448634 303914 448718
rect 303294 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 303914 448634
rect 303294 412954 303914 448398
rect 303294 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 303914 412954
rect 303294 412634 303914 412718
rect 303294 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 303914 412634
rect 303294 376954 303914 412398
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 303294 340954 303914 376398
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 303294 304954 303914 340398
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 232954 303914 268398
rect 303294 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 303914 232954
rect 303294 232634 303914 232718
rect 303294 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 303914 232634
rect 303294 196954 303914 232398
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 178000 308414 200898
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 529954 312914 565398
rect 312294 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 312914 529954
rect 312294 529634 312914 529718
rect 312294 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 312914 529634
rect 312294 493954 312914 529398
rect 312294 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 312914 493954
rect 312294 493634 312914 493718
rect 312294 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 312914 493634
rect 312294 457954 312914 493398
rect 312294 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 312914 457954
rect 312294 457634 312914 457718
rect 312294 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 312914 457634
rect 312294 421954 312914 457398
rect 312294 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 312914 421954
rect 312294 421634 312914 421718
rect 312294 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 312914 421634
rect 312294 385954 312914 421398
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 313954 312914 349398
rect 312294 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 312914 313954
rect 312294 313634 312914 313718
rect 312294 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 312914 313634
rect 312294 277954 312914 313398
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 241954 312914 277398
rect 312294 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 312914 241954
rect 312294 241634 312914 241718
rect 312294 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 312914 241634
rect 312294 205954 312914 241398
rect 312294 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 312914 205954
rect 312294 205634 312914 205718
rect 312294 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 312914 205634
rect 312294 178000 312914 205398
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 534454 317414 569898
rect 316794 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 317414 534454
rect 316794 534134 317414 534218
rect 316794 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 317414 534134
rect 316794 498454 317414 533898
rect 316794 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 317414 498454
rect 316794 498134 317414 498218
rect 316794 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 317414 498134
rect 316794 462454 317414 497898
rect 316794 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 317414 462454
rect 316794 462134 317414 462218
rect 316794 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 317414 462134
rect 316794 426454 317414 461898
rect 316794 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 317414 426454
rect 316794 426134 317414 426218
rect 316794 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 317414 426134
rect 316794 390454 317414 425898
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 318454 317414 353898
rect 316794 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 317414 318454
rect 316794 318134 317414 318218
rect 316794 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 317414 318134
rect 316794 282454 317414 317898
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 246454 317414 281898
rect 316794 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 317414 246454
rect 316794 246134 317414 246218
rect 316794 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 317414 246134
rect 316794 210454 317414 245898
rect 316794 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 317414 210454
rect 316794 210134 317414 210218
rect 316794 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 317414 210134
rect 316794 178000 317414 209898
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 538954 321914 574398
rect 321294 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 321914 538954
rect 321294 538634 321914 538718
rect 321294 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 321914 538634
rect 321294 502954 321914 538398
rect 321294 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 321914 502954
rect 321294 502634 321914 502718
rect 321294 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 321914 502634
rect 321294 466954 321914 502398
rect 321294 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 321914 466954
rect 321294 466634 321914 466718
rect 321294 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 321914 466634
rect 321294 430954 321914 466398
rect 321294 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 321914 430954
rect 321294 430634 321914 430718
rect 321294 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 321914 430634
rect 321294 394954 321914 430398
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 322954 321914 358398
rect 321294 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 321914 322954
rect 321294 322634 321914 322718
rect 321294 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 321914 322634
rect 321294 286954 321914 322398
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 214954 321914 250398
rect 321294 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 321914 214954
rect 321294 214634 321914 214718
rect 321294 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 321914 214634
rect 320219 186964 320285 186965
rect 320219 186900 320220 186964
rect 320284 186900 320285 186964
rect 320219 186899 320285 186900
rect 306971 175676 307037 175677
rect 306971 175612 306972 175676
rect 307036 175612 307037 175676
rect 306971 175611 307037 175612
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 301451 130660 301517 130661
rect 301451 130596 301452 130660
rect 301516 130596 301517 130660
rect 301451 130595 301517 130596
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 297219 115292 297285 115293
rect 297219 115228 297220 115292
rect 297284 115228 297285 115292
rect 297219 115227 297285 115228
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 297222 69597 297282 115227
rect 298794 84454 299414 119898
rect 299979 99652 300045 99653
rect 299979 99588 299980 99652
rect 300044 99588 300045 99652
rect 299979 99587 300045 99588
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 297219 69596 297285 69597
rect 297219 69532 297220 69596
rect 297284 69532 297285 69596
rect 297219 69531 297285 69532
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 299982 22677 300042 99587
rect 301454 75173 301514 130595
rect 303294 124954 303914 160398
rect 306974 144125 307034 175611
rect 320222 170370 320282 186899
rect 321294 178954 321914 214398
rect 321294 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 321914 178954
rect 321294 178634 321914 178718
rect 321294 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 321914 178634
rect 321294 178000 321914 178398
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 511954 330914 547398
rect 330294 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 330914 511954
rect 330294 511634 330914 511718
rect 330294 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 330914 511634
rect 330294 475954 330914 511398
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 330294 439954 330914 475398
rect 330294 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 330914 439954
rect 330294 439634 330914 439718
rect 330294 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 330914 439634
rect 330294 403954 330914 439398
rect 330294 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 330914 403954
rect 330294 403634 330914 403718
rect 330294 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 330914 403634
rect 330294 367954 330914 403398
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 331954 330914 367398
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 552454 335414 587898
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 516454 335414 551898
rect 334794 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 335414 516454
rect 334794 516134 335414 516218
rect 334794 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 335414 516134
rect 334794 480454 335414 515898
rect 334794 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 335414 480454
rect 334794 480134 335414 480218
rect 334794 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 335414 480134
rect 334794 444454 335414 479898
rect 334794 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 335414 444454
rect 334794 444134 335414 444218
rect 334794 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 335414 444134
rect 334794 408454 335414 443898
rect 334794 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 335414 408454
rect 334794 408134 335414 408218
rect 334794 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 335414 408134
rect 334794 372454 335414 407898
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 334794 336454 335414 371898
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 331259 302292 331325 302293
rect 331259 302228 331260 302292
rect 331324 302228 331325 302292
rect 331259 302227 331325 302228
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 329787 224228 329853 224229
rect 329787 224164 329788 224228
rect 329852 224164 329853 224228
rect 329787 224163 329853 224164
rect 328499 221508 328565 221509
rect 328499 221444 328500 221508
rect 328564 221444 328565 221508
rect 328499 221443 328565 221444
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 327027 204916 327093 204917
rect 327027 204852 327028 204916
rect 327092 204852 327093 204916
rect 327027 204851 327093 204852
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 321323 176764 321389 176765
rect 321323 176700 321324 176764
rect 321388 176700 321389 176764
rect 321323 176699 321389 176700
rect 321326 171053 321386 176699
rect 321507 176220 321573 176221
rect 321507 176156 321508 176220
rect 321572 176156 321573 176220
rect 321507 176155 321573 176156
rect 321510 174453 321570 176155
rect 321507 174452 321573 174453
rect 321507 174388 321508 174452
rect 321572 174388 321573 174452
rect 321507 174387 321573 174388
rect 321323 171052 321389 171053
rect 321323 170988 321324 171052
rect 321388 170988 321389 171052
rect 321323 170987 321389 170988
rect 321323 170372 321389 170373
rect 321323 170370 321324 170372
rect 320222 170310 321324 170370
rect 321323 170308 321324 170310
rect 321388 170308 321389 170372
rect 321323 170307 321389 170308
rect 314208 151954 314528 151986
rect 314208 151718 314250 151954
rect 314486 151718 314528 151954
rect 314208 151634 314528 151718
rect 314208 151398 314250 151634
rect 314486 151398 314528 151634
rect 314208 151366 314528 151398
rect 317472 151954 317792 151986
rect 317472 151718 317514 151954
rect 317750 151718 317792 151954
rect 317472 151634 317792 151718
rect 317472 151398 317514 151634
rect 317750 151398 317792 151634
rect 317472 151366 317792 151398
rect 312576 147454 312896 147486
rect 312576 147218 312618 147454
rect 312854 147218 312896 147454
rect 312576 147134 312896 147218
rect 312576 146898 312618 147134
rect 312854 146898 312896 147134
rect 312576 146866 312896 146898
rect 315840 147454 316160 147486
rect 315840 147218 315882 147454
rect 316118 147218 316160 147454
rect 315840 147134 316160 147218
rect 315840 146898 315882 147134
rect 316118 146898 316160 147134
rect 315840 146866 316160 146898
rect 319104 147454 319424 147486
rect 319104 147218 319146 147454
rect 319382 147218 319424 147454
rect 319104 147134 319424 147218
rect 319104 146898 319146 147134
rect 319382 146898 319424 147134
rect 319104 146866 319424 146898
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 306971 144124 307037 144125
rect 306971 144060 306972 144124
rect 307036 144060 307037 144124
rect 306971 144059 307037 144060
rect 307707 143852 307773 143853
rect 307707 143788 307708 143852
rect 307772 143788 307773 143852
rect 307707 143787 307773 143788
rect 307710 142765 307770 143787
rect 307707 142764 307773 142765
rect 307707 142700 307708 142764
rect 307772 142700 307773 142764
rect 307707 142699 307773 142700
rect 306419 142492 306485 142493
rect 306419 142428 306420 142492
rect 306484 142428 306485 142492
rect 306419 142427 306485 142428
rect 306422 141405 306482 142427
rect 306419 141404 306485 141405
rect 306419 141340 306420 141404
rect 306484 141340 306485 141404
rect 306419 141339 306485 141340
rect 307707 140860 307773 140861
rect 307707 140796 307708 140860
rect 307772 140796 307773 140860
rect 307707 140795 307773 140796
rect 307710 133109 307770 140795
rect 307707 133108 307773 133109
rect 307707 133044 307708 133108
rect 307772 133044 307773 133108
rect 307707 133043 307773 133044
rect 306971 132700 307037 132701
rect 306971 132636 306972 132700
rect 307036 132636 307037 132700
rect 306971 132635 307037 132636
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 302739 96660 302805 96661
rect 302739 96596 302740 96660
rect 302804 96596 302805 96660
rect 302739 96595 302805 96596
rect 301451 75172 301517 75173
rect 301451 75108 301452 75172
rect 301516 75108 301517 75172
rect 301451 75107 301517 75108
rect 302742 61437 302802 96595
rect 303294 88954 303914 124398
rect 304211 118284 304277 118285
rect 304211 118220 304212 118284
rect 304276 118220 304277 118284
rect 304211 118219 304277 118220
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 302739 61436 302805 61437
rect 302739 61372 302740 61436
rect 302804 61372 302805 61436
rect 302739 61371 302805 61372
rect 303294 52954 303914 88398
rect 304214 64157 304274 118219
rect 305499 112708 305565 112709
rect 305499 112644 305500 112708
rect 305564 112644 305565 112708
rect 305499 112643 305565 112644
rect 304211 64156 304277 64157
rect 304211 64092 304212 64156
rect 304276 64092 304277 64156
rect 304211 64091 304277 64092
rect 305502 57221 305562 112643
rect 305683 101284 305749 101285
rect 305683 101220 305684 101284
rect 305748 101220 305749 101284
rect 305683 101219 305749 101220
rect 305686 65517 305746 101219
rect 305683 65516 305749 65517
rect 305683 65452 305684 65516
rect 305748 65452 305749 65516
rect 305683 65451 305749 65452
rect 305499 57220 305565 57221
rect 305499 57156 305500 57220
rect 305564 57156 305565 57220
rect 305499 57155 305565 57156
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 299979 22676 300045 22677
rect 299979 22612 299980 22676
rect 300044 22612 300045 22676
rect 299979 22611 300045 22612
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 16954 303914 52398
rect 306974 43485 307034 132635
rect 314208 115954 314528 115986
rect 314208 115718 314250 115954
rect 314486 115718 314528 115954
rect 314208 115634 314528 115718
rect 314208 115398 314250 115634
rect 314486 115398 314528 115634
rect 314208 115366 314528 115398
rect 317472 115954 317792 115986
rect 317472 115718 317514 115954
rect 317750 115718 317792 115954
rect 317472 115634 317792 115718
rect 317472 115398 317514 115634
rect 317750 115398 317792 115634
rect 317472 115366 317792 115398
rect 307155 114068 307221 114069
rect 307155 114004 307156 114068
rect 307220 114004 307221 114068
rect 307155 114003 307221 114004
rect 307158 46205 307218 114003
rect 312576 111454 312896 111486
rect 312576 111218 312618 111454
rect 312854 111218 312896 111454
rect 312576 111134 312896 111218
rect 312576 110898 312618 111134
rect 312854 110898 312896 111134
rect 312576 110866 312896 110898
rect 315840 111454 316160 111486
rect 315840 111218 315882 111454
rect 316118 111218 316160 111454
rect 315840 111134 316160 111218
rect 315840 110898 315882 111134
rect 316118 110898 316160 111134
rect 315840 110866 316160 110898
rect 319104 111454 319424 111486
rect 319104 111218 319146 111454
rect 319382 111218 319424 111454
rect 319104 111134 319424 111218
rect 319104 110898 319146 111134
rect 319382 110898 319424 111134
rect 319104 110866 319424 110898
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 324267 104820 324333 104821
rect 324267 104756 324268 104820
rect 324332 104756 324333 104820
rect 324267 104755 324333 104756
rect 324270 95981 324330 104755
rect 324267 95980 324333 95981
rect 324267 95916 324268 95980
rect 324332 95916 324333 95980
rect 324267 95915 324333 95916
rect 307794 93454 308414 94000
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307155 46204 307221 46205
rect 307155 46140 307156 46204
rect 307220 46140 307221 46204
rect 307155 46139 307221 46140
rect 306971 43484 307037 43485
rect 306971 43420 306972 43484
rect 307036 43420 307037 43484
rect 306971 43419 307037 43420
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 61954 312914 94000
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 66454 317414 94000
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 70954 321914 94000
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 75454 326414 110898
rect 327030 104005 327090 204851
rect 327211 189684 327277 189685
rect 327211 189620 327212 189684
rect 327276 189620 327277 189684
rect 327211 189619 327277 189620
rect 327214 129437 327274 189619
rect 327211 129436 327277 129437
rect 327211 129372 327212 129436
rect 327276 129372 327277 129436
rect 327211 129371 327277 129372
rect 328502 106453 328562 221443
rect 329790 127125 329850 224163
rect 330294 223954 330914 259398
rect 330294 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 330914 223954
rect 330294 223634 330914 223718
rect 330294 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 330914 223634
rect 330294 187954 330914 223398
rect 330294 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 330914 187954
rect 330294 187634 330914 187718
rect 330294 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 330914 187634
rect 330294 151954 330914 187398
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 329787 127124 329853 127125
rect 329787 127060 329788 127124
rect 329852 127060 329853 127124
rect 329787 127059 329853 127060
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 328499 106452 328565 106453
rect 328499 106388 328500 106452
rect 328564 106388 328565 106452
rect 328499 106387 328565 106388
rect 327027 104004 327093 104005
rect 327027 103940 327028 104004
rect 327092 103940 327093 104004
rect 327027 103939 327093 103940
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 79954 330914 115398
rect 331262 98701 331322 302227
rect 334794 300454 335414 335898
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 556954 339914 592398
rect 339294 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 339914 556954
rect 339294 556634 339914 556718
rect 339294 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 339914 556634
rect 339294 520954 339914 556398
rect 339294 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 339914 520954
rect 339294 520634 339914 520718
rect 339294 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 339914 520634
rect 339294 484954 339914 520398
rect 339294 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 339914 484954
rect 339294 484634 339914 484718
rect 339294 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 339914 484634
rect 339294 448954 339914 484398
rect 339294 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 339914 448954
rect 339294 448634 339914 448718
rect 339294 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 339914 448634
rect 339294 412954 339914 448398
rect 339294 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 339914 412954
rect 339294 412634 339914 412718
rect 339294 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 339914 412634
rect 339294 376954 339914 412398
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 339294 340954 339914 376398
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 304954 339914 340398
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 335675 291956 335741 291957
rect 335675 291892 335676 291956
rect 335740 291892 335741 291956
rect 335675 291891 335741 291892
rect 335678 277410 335738 291891
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 332547 232524 332613 232525
rect 332547 232460 332548 232524
rect 332612 232460 332613 232524
rect 332547 232459 332613 232460
rect 331443 177308 331509 177309
rect 331443 177244 331444 177308
rect 331508 177244 331509 177308
rect 331443 177243 331509 177244
rect 331446 142765 331506 177243
rect 331443 142764 331509 142765
rect 331443 142700 331444 142764
rect 331508 142700 331509 142764
rect 331443 142699 331509 142700
rect 332550 101013 332610 232459
rect 334794 228454 335414 263898
rect 334794 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 335414 228454
rect 334794 228134 335414 228218
rect 334794 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 335414 228134
rect 334794 192454 335414 227898
rect 334794 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 335414 192454
rect 334794 192134 335414 192218
rect 334794 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 335414 192134
rect 334019 181388 334085 181389
rect 334019 181324 334020 181388
rect 334084 181324 334085 181388
rect 334019 181323 334085 181324
rect 332731 178804 332797 178805
rect 332731 178740 332732 178804
rect 332796 178740 332797 178804
rect 332731 178739 332797 178740
rect 332734 109581 332794 178739
rect 332731 109580 332797 109581
rect 332731 109516 332732 109580
rect 332796 109516 332797 109580
rect 332731 109515 332797 109516
rect 334022 102373 334082 181323
rect 334794 156454 335414 191898
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334019 102372 334085 102373
rect 334019 102308 334020 102372
rect 334084 102308 334085 102372
rect 334019 102307 334085 102308
rect 332547 101012 332613 101013
rect 332547 100948 332548 101012
rect 332612 100948 332613 101012
rect 332547 100947 332613 100948
rect 331259 98700 331325 98701
rect 331259 98636 331260 98700
rect 331324 98636 331325 98700
rect 331259 98635 331325 98636
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 84454 335414 119898
rect 335494 277350 335738 277410
rect 335494 109170 335554 277350
rect 339294 268954 339914 304398
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 340827 295356 340893 295357
rect 340827 295292 340828 295356
rect 340892 295292 340893 295356
rect 340827 295291 340893 295292
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 337331 259588 337397 259589
rect 337331 259524 337332 259588
rect 337396 259524 337397 259588
rect 337331 259523 337397 259524
rect 335675 206276 335741 206277
rect 335675 206212 335676 206276
rect 335740 206212 335741 206276
rect 335675 206211 335741 206212
rect 335678 142221 335738 206211
rect 336779 178668 336845 178669
rect 336779 178604 336780 178668
rect 336844 178604 336845 178668
rect 336779 178603 336845 178604
rect 335675 142220 335741 142221
rect 335675 142156 335676 142220
rect 335740 142156 335741 142220
rect 335675 142155 335741 142156
rect 336782 110533 336842 178603
rect 337334 165749 337394 259523
rect 339294 232954 339914 268398
rect 339294 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 339914 232954
rect 339294 232634 339914 232718
rect 339294 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 339914 232634
rect 338251 197980 338317 197981
rect 338251 197916 338252 197980
rect 338316 197916 338317 197980
rect 338251 197915 338317 197916
rect 337331 165748 337397 165749
rect 337331 165684 337332 165748
rect 337396 165684 337397 165748
rect 337331 165683 337397 165684
rect 338254 114613 338314 197915
rect 339294 196954 339914 232398
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 339294 160954 339914 196398
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 339294 124954 339914 160398
rect 340830 134197 340890 295291
rect 343794 273454 344414 308898
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 529954 348914 565398
rect 348294 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 348914 529954
rect 348294 529634 348914 529718
rect 348294 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 348914 529634
rect 348294 493954 348914 529398
rect 348294 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 348914 493954
rect 348294 493634 348914 493718
rect 348294 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 348914 493634
rect 348294 457954 348914 493398
rect 348294 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 348914 457954
rect 348294 457634 348914 457718
rect 348294 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 348914 457634
rect 348294 421954 348914 457398
rect 348294 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 348914 421954
rect 348294 421634 348914 421718
rect 348294 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 348914 421634
rect 348294 385954 348914 421398
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 313954 348914 349398
rect 348294 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 348914 313954
rect 348294 313634 348914 313718
rect 348294 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 348914 313634
rect 346163 291276 346229 291277
rect 346163 291212 346164 291276
rect 346228 291212 346229 291276
rect 346163 291211 346229 291212
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 342299 196620 342365 196621
rect 342299 196556 342300 196620
rect 342364 196556 342365 196620
rect 342299 196555 342365 196556
rect 340827 134196 340893 134197
rect 340827 134132 340828 134196
rect 340892 134132 340893 134196
rect 340827 134131 340893 134132
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 338251 114612 338317 114613
rect 338251 114548 338252 114612
rect 338316 114548 338317 114612
rect 338251 114547 338317 114548
rect 336779 110532 336845 110533
rect 336779 110468 336780 110532
rect 336844 110468 336845 110532
rect 336779 110467 336845 110468
rect 335675 109172 335741 109173
rect 335675 109170 335676 109172
rect 335494 109110 335676 109170
rect 335675 109108 335676 109110
rect 335740 109108 335741 109172
rect 335675 109107 335741 109108
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 88954 339914 124398
rect 342302 106317 342362 196555
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 346166 138141 346226 291211
rect 348294 277954 348914 313398
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 241954 348914 277398
rect 348294 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 348914 241954
rect 348294 241634 348914 241718
rect 348294 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 348914 241634
rect 348294 205954 348914 241398
rect 348294 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 348914 205954
rect 348294 205634 348914 205718
rect 348294 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 348914 205634
rect 348294 169954 348914 205398
rect 348294 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 348914 169954
rect 348294 169634 348914 169718
rect 348294 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 348914 169634
rect 346163 138140 346229 138141
rect 346163 138076 346164 138140
rect 346228 138076 346229 138140
rect 346163 138075 346229 138076
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 342299 106316 342365 106317
rect 342299 106252 342300 106316
rect 342364 106252 342365 106316
rect 342299 106251 342365 106252
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 133954 348914 169398
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 534454 353414 569898
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 352794 498454 353414 533898
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 426454 353414 461898
rect 352794 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 353414 426454
rect 352794 426134 353414 426218
rect 352794 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 353414 426134
rect 352794 390454 353414 425898
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 210454 353414 245898
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 138454 353414 173898
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 538954 357914 574398
rect 357294 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 357914 538954
rect 357294 538634 357914 538718
rect 357294 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 357914 538634
rect 357294 502954 357914 538398
rect 357294 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 357914 502954
rect 357294 502634 357914 502718
rect 357294 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 357914 502634
rect 357294 466954 357914 502398
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 430954 357914 466398
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 357294 430634 357914 430718
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 214954 357914 250398
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 241954 384914 277398
rect 384294 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 384914 241954
rect 384294 241634 384914 241718
rect 384294 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 384914 241634
rect 384294 205954 384914 241398
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 210454 389414 245898
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 214954 393914 250398
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 580211 246260 580277 246261
rect 580211 246196 580212 246260
rect 580276 246196 580277 246260
rect 580211 246195 580277 246196
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 580214 72997 580274 246195
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 580211 72996 580277 72997
rect 580211 72932 580212 72996
rect 580276 72932 580277 72996
rect 580211 72931 580277 72932
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< obsm4 >>
rect 68800 174494 96960 174600
rect 97020 174494 98320 174600
rect 98380 174494 99408 174600
rect 99468 174494 100768 174600
rect 100828 174494 101992 174600
rect 102052 174494 103352 174600
rect 103412 174494 104576 174600
rect 104636 174494 105664 174600
rect 105724 174494 107024 174600
rect 107084 174494 108112 174600
rect 108172 174494 109472 174600
rect 109532 174494 110696 174600
rect 110756 174494 112056 174600
rect 112116 174494 113144 174600
rect 113204 174494 114368 174600
rect 114428 174494 115728 174600
rect 115788 174494 116952 174600
rect 117012 174494 118312 174600
rect 118372 174494 119400 174600
rect 119460 174494 120760 174600
rect 120820 174494 121848 174600
rect 121908 174494 123072 174600
rect 123132 174494 124432 174600
rect 124492 174494 125656 174600
rect 125716 174494 127016 174600
rect 127076 174494 128104 174600
rect 128164 174494 129464 174600
rect 129524 174494 130688 174600
rect 130748 174494 132048 174600
rect 132108 174494 133136 174600
rect 133196 174494 134360 174600
rect 134420 174494 135720 174600
rect 135780 174494 148232 174600
rect 148292 174494 158840 174600
rect 158900 174494 164756 174600
rect 68800 151986 164756 174494
rect 68800 151366 69072 151986
rect 69420 151366 164136 151986
rect 164484 151366 164756 151986
rect 68800 147486 164756 151366
rect 68800 146866 69752 147486
rect 70100 146866 163456 147486
rect 163804 146866 164756 147486
rect 68800 115986 164756 146866
rect 68800 115366 69072 115986
rect 69420 115366 164136 115986
rect 164484 115366 164756 115986
rect 68800 111486 164756 115366
rect 68800 110866 69752 111486
rect 70100 110866 163456 111486
rect 163804 110866 164756 111486
rect 68800 95200 164756 110866
rect 68800 95100 74656 95200
rect 74716 95100 84312 95200
rect 84372 95100 85536 95200
rect 85596 95100 86624 95200
rect 86684 95100 87984 95200
rect 88044 95100 88936 95200
rect 88996 95100 90160 95200
rect 90220 95100 91384 95200
rect 91444 95100 92472 95200
rect 92532 95100 93832 95200
rect 93892 95100 94920 95200
rect 94980 95100 96008 95200
rect 96068 95100 96688 95200
rect 96748 95100 97096 95200
rect 97156 95100 98048 95200
rect 98108 95100 98456 95200
rect 98516 95100 99136 95200
rect 99196 95100 99544 95200
rect 99604 95100 100632 95200
rect 100692 95100 100768 95200
rect 100828 95100 101856 95200
rect 101916 95100 101992 95200
rect 102052 95100 102944 95200
rect 103004 95100 103216 95200
rect 103276 95100 104304 95200
rect 104364 95100 104440 95200
rect 104500 95100 105392 95200
rect 105452 95100 105664 95200
rect 105724 95100 106480 95200
rect 106540 95100 106616 95200
rect 106676 95100 107704 95200
rect 107764 95100 108112 95200
rect 108172 95100 109064 95200
rect 109124 95100 109472 95200
rect 109532 95100 110152 95200
rect 110212 95100 110696 95200
rect 110756 95100 111240 95200
rect 111300 95100 111920 95200
rect 111980 95100 112328 95200
rect 112388 95100 113144 95200
rect 113204 95100 113688 95200
rect 113748 95100 114368 95200
rect 114428 95100 114776 95200
rect 114836 95100 115456 95200
rect 115516 95100 115864 95200
rect 115924 95100 116680 95200
rect 116740 95100 117088 95200
rect 117148 95100 117904 95200
rect 117964 95100 118176 95200
rect 118236 95100 119400 95200
rect 119460 95100 119536 95200
rect 119596 95100 120216 95200
rect 120276 95100 120624 95200
rect 120684 95100 121712 95200
rect 121772 95100 121984 95200
rect 122044 95100 122800 95200
rect 122860 95100 123208 95200
rect 123268 95100 124024 95200
rect 124084 95100 124432 95200
rect 124492 95100 125384 95200
rect 125444 95100 125656 95200
rect 125716 95100 126472 95200
rect 126532 95100 126608 95200
rect 126668 95100 128104 95200
rect 128164 95100 129328 95200
rect 129388 95100 130688 95200
rect 130748 95100 131912 95200
rect 131972 95100 133136 95200
rect 133196 95100 134360 95200
rect 134420 95100 135584 95200
rect 135644 95100 151496 95200
rect 151556 95100 151632 95200
rect 151692 95100 151768 95200
rect 151828 95100 151904 95200
rect 151964 95100 164756 95200
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 89610 259718 89846 259954
rect 89610 259398 89846 259634
rect 74250 255218 74486 255454
rect 74250 254898 74486 255134
rect 104970 255218 105206 255454
rect 104970 254898 105206 255134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 118826 228218 119062 228454
rect 119146 228218 119382 228454
rect 118826 227898 119062 228134
rect 119146 227898 119382 228134
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 123326 232718 123562 232954
rect 123646 232718 123882 232954
rect 123326 232398 123562 232634
rect 123646 232398 123882 232634
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 132326 241718 132562 241954
rect 132646 241718 132882 241954
rect 132326 241398 132562 241634
rect 132646 241398 132882 241634
rect 132326 205718 132562 205954
rect 132646 205718 132882 205954
rect 132326 205398 132562 205634
rect 132646 205398 132882 205634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 136826 246218 137062 246454
rect 137146 246218 137382 246454
rect 136826 245898 137062 246134
rect 137146 245898 137382 246134
rect 136826 210218 137062 210454
rect 137146 210218 137382 210454
rect 136826 209898 137062 210134
rect 137146 209898 137382 210134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 141326 214718 141562 214954
rect 141646 214718 141882 214954
rect 141326 214398 141562 214634
rect 141646 214398 141882 214634
rect 141326 178718 141562 178954
rect 141646 178718 141882 178954
rect 141326 178398 141562 178634
rect 141646 178398 141882 178634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 150326 223718 150562 223954
rect 150646 223718 150882 223954
rect 150326 223398 150562 223634
rect 150646 223398 150882 223634
rect 150326 187718 150562 187954
rect 150646 187718 150882 187954
rect 150326 187398 150562 187634
rect 150646 187398 150882 187634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 154826 228218 155062 228454
rect 155146 228218 155382 228454
rect 154826 227898 155062 228134
rect 155146 227898 155382 228134
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 159326 232718 159562 232954
rect 159646 232718 159882 232954
rect 159326 232398 159562 232634
rect 159646 232398 159882 232634
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 168326 241718 168562 241954
rect 168646 241718 168882 241954
rect 168326 241398 168562 241634
rect 168646 241398 168882 241634
rect 168326 205718 168562 205954
rect 168646 205718 168882 205954
rect 168326 205398 168562 205634
rect 168646 205398 168882 205634
rect 168326 169718 168562 169954
rect 168646 169718 168882 169954
rect 168326 169398 168562 169634
rect 168646 169398 168882 169634
rect 69128 151718 69364 151954
rect 69128 151398 69364 151634
rect 164192 151718 164428 151954
rect 164192 151398 164428 151634
rect 69808 147218 70044 147454
rect 69808 146898 70044 147134
rect 163512 147218 163748 147454
rect 163512 146898 163748 147134
rect 69128 115718 69364 115954
rect 69128 115398 69364 115634
rect 164192 115718 164428 115954
rect 164192 115398 164428 115634
rect 69808 111218 70044 111454
rect 69808 110898 70044 111134
rect 163512 111218 163748 111454
rect 163512 110898 163748 111134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 84218 119062 84454
rect 119146 84218 119382 84454
rect 118826 83898 119062 84134
rect 119146 83898 119382 84134
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 88718 123562 88954
rect 123646 88718 123882 88954
rect 123326 88398 123562 88634
rect 123646 88398 123882 88634
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 79718 150562 79954
rect 150646 79718 150882 79954
rect 150326 79398 150562 79634
rect 150646 79398 150882 79634
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 154826 84218 155062 84454
rect 155146 84218 155382 84454
rect 154826 83898 155062 84134
rect 155146 83898 155382 84134
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 159326 88718 159562 88954
rect 159646 88718 159882 88954
rect 159326 88398 159562 88634
rect 159646 88398 159882 88634
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 172826 246218 173062 246454
rect 173146 246218 173382 246454
rect 172826 245898 173062 246134
rect 173146 245898 173382 246134
rect 172826 210218 173062 210454
rect 173146 210218 173382 210454
rect 172826 209898 173062 210134
rect 173146 209898 173382 210134
rect 172826 174218 173062 174454
rect 173146 174218 173382 174454
rect 172826 173898 173062 174134
rect 173146 173898 173382 174134
rect 172826 138218 173062 138454
rect 173146 138218 173382 138454
rect 172826 137898 173062 138134
rect 173146 137898 173382 138134
rect 168326 133718 168562 133954
rect 168646 133718 168882 133954
rect 168326 133398 168562 133634
rect 168646 133398 168882 133634
rect 168326 97718 168562 97954
rect 168646 97718 168882 97954
rect 168326 97398 168562 97634
rect 168646 97398 168882 97634
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 172826 102218 173062 102454
rect 173146 102218 173382 102454
rect 172826 101898 173062 102134
rect 173146 101898 173382 102134
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 177326 214718 177562 214954
rect 177646 214718 177882 214954
rect 177326 214398 177562 214634
rect 177646 214398 177882 214634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 177326 106718 177562 106954
rect 177646 106718 177882 106954
rect 177326 106398 177562 106634
rect 177646 106398 177882 106634
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 186326 259718 186562 259954
rect 186646 259718 186882 259954
rect 186326 259398 186562 259634
rect 186646 259398 186882 259634
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 186326 115718 186562 115954
rect 186646 115718 186882 115954
rect 186326 115398 186562 115634
rect 186646 115398 186882 115634
rect 186326 79718 186562 79954
rect 186646 79718 186882 79954
rect 186326 79398 186562 79634
rect 186646 79398 186882 79634
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 190826 228218 191062 228454
rect 191146 228218 191382 228454
rect 190826 227898 191062 228134
rect 191146 227898 191382 228134
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 190826 120218 191062 120454
rect 191146 120218 191382 120454
rect 190826 119898 191062 120134
rect 191146 119898 191382 120134
rect 190826 84218 191062 84454
rect 191146 84218 191382 84454
rect 190826 83898 191062 84134
rect 191146 83898 191382 84134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 195326 232718 195562 232954
rect 195646 232718 195882 232954
rect 195326 232398 195562 232634
rect 195646 232398 195882 232634
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 204326 241718 204562 241954
rect 204646 241718 204882 241954
rect 204326 241398 204562 241634
rect 204646 241398 204882 241634
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 208826 246218 209062 246454
rect 209146 246218 209382 246454
rect 208826 245898 209062 246134
rect 209146 245898 209382 246134
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 222326 547718 222562 547954
rect 222646 547718 222882 547954
rect 222326 547398 222562 547634
rect 222646 547398 222882 547634
rect 222326 511718 222562 511954
rect 222646 511718 222882 511954
rect 222326 511398 222562 511634
rect 222646 511398 222882 511634
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 226826 552218 227062 552454
rect 227146 552218 227382 552454
rect 226826 551898 227062 552134
rect 227146 551898 227382 552134
rect 226826 516218 227062 516454
rect 227146 516218 227382 516454
rect 226826 515898 227062 516134
rect 227146 515898 227382 516134
rect 226826 480218 227062 480454
rect 227146 480218 227382 480454
rect 226826 479898 227062 480134
rect 227146 479898 227382 480134
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 226826 228218 227062 228454
rect 227146 228218 227382 228454
rect 226826 227898 227062 228134
rect 227146 227898 227382 228134
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 231326 556718 231562 556954
rect 231646 556718 231882 556954
rect 231326 556398 231562 556634
rect 231646 556398 231882 556634
rect 231326 520718 231562 520954
rect 231646 520718 231882 520954
rect 231326 520398 231562 520634
rect 231646 520398 231882 520634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 231326 412718 231562 412954
rect 231646 412718 231882 412954
rect 231326 412398 231562 412634
rect 231646 412398 231882 412634
rect 231326 376718 231562 376954
rect 231646 376718 231882 376954
rect 231326 376398 231562 376634
rect 231646 376398 231882 376634
rect 231326 340718 231562 340954
rect 231646 340718 231882 340954
rect 231326 340398 231562 340634
rect 231646 340398 231882 340634
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 231326 232718 231562 232954
rect 231646 232718 231882 232954
rect 231326 232398 231562 232634
rect 231646 232398 231882 232634
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 240326 529718 240562 529954
rect 240646 529718 240882 529954
rect 240326 529398 240562 529634
rect 240646 529398 240882 529634
rect 240326 493718 240562 493954
rect 240646 493718 240882 493954
rect 240326 493398 240562 493634
rect 240646 493398 240882 493634
rect 240326 457718 240562 457954
rect 240646 457718 240882 457954
rect 240326 457398 240562 457634
rect 240646 457398 240882 457634
rect 240326 421718 240562 421954
rect 240646 421718 240882 421954
rect 240326 421398 240562 421634
rect 240646 421398 240882 421634
rect 240326 385718 240562 385954
rect 240646 385718 240882 385954
rect 240326 385398 240562 385634
rect 240646 385398 240882 385634
rect 240326 349718 240562 349954
rect 240646 349718 240882 349954
rect 240326 349398 240562 349634
rect 240646 349398 240882 349634
rect 240326 313718 240562 313954
rect 240646 313718 240882 313954
rect 240326 313398 240562 313634
rect 240646 313398 240882 313634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 240326 241718 240562 241954
rect 240646 241718 240882 241954
rect 240326 241398 240562 241634
rect 240646 241398 240882 241634
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 244826 534218 245062 534454
rect 245146 534218 245382 534454
rect 244826 533898 245062 534134
rect 245146 533898 245382 534134
rect 244826 498218 245062 498454
rect 245146 498218 245382 498454
rect 244826 497898 245062 498134
rect 245146 497898 245382 498134
rect 244826 462218 245062 462454
rect 245146 462218 245382 462454
rect 244826 461898 245062 462134
rect 245146 461898 245382 462134
rect 244826 426218 245062 426454
rect 245146 426218 245382 426454
rect 244826 425898 245062 426134
rect 245146 425898 245382 426134
rect 244826 390218 245062 390454
rect 245146 390218 245382 390454
rect 244826 389898 245062 390134
rect 245146 389898 245382 390134
rect 244826 354218 245062 354454
rect 245146 354218 245382 354454
rect 244826 353898 245062 354134
rect 245146 353898 245382 354134
rect 244826 318218 245062 318454
rect 245146 318218 245382 318454
rect 244826 317898 245062 318134
rect 245146 317898 245382 318134
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 244826 246218 245062 246454
rect 245146 246218 245382 246454
rect 244826 245898 245062 246134
rect 245146 245898 245382 246134
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 249326 538718 249562 538954
rect 249646 538718 249882 538954
rect 249326 538398 249562 538634
rect 249646 538398 249882 538634
rect 249326 502718 249562 502954
rect 249646 502718 249882 502954
rect 249326 502398 249562 502634
rect 249646 502398 249882 502634
rect 249326 466718 249562 466954
rect 249646 466718 249882 466954
rect 249326 466398 249562 466634
rect 249646 466398 249882 466634
rect 249326 430718 249562 430954
rect 249646 430718 249882 430954
rect 249326 430398 249562 430634
rect 249646 430398 249882 430634
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 249326 358718 249562 358954
rect 249646 358718 249882 358954
rect 249326 358398 249562 358634
rect 249646 358398 249882 358634
rect 249326 322718 249562 322954
rect 249646 322718 249882 322954
rect 249326 322398 249562 322634
rect 249646 322398 249882 322634
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 227916 151718 228152 151954
rect 227916 151398 228152 151634
rect 237847 151718 238083 151954
rect 237847 151398 238083 151634
rect 222952 147218 223188 147454
rect 222952 146898 223188 147134
rect 232882 147218 233118 147454
rect 232882 146898 233118 147134
rect 242813 147218 243049 147454
rect 242813 146898 243049 147134
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 227916 115718 228152 115954
rect 227916 115398 228152 115634
rect 237847 115718 238083 115954
rect 237847 115398 238083 115634
rect 222952 111218 223188 111454
rect 222952 110898 223188 111134
rect 232882 111218 233118 111454
rect 232882 110898 233118 111134
rect 242813 111218 243049 111454
rect 242813 110898 243049 111134
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 258326 331718 258562 331954
rect 258646 331718 258882 331954
rect 258326 331398 258562 331634
rect 258646 331398 258882 331634
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 262826 336218 263062 336454
rect 263146 336218 263382 336454
rect 262826 335898 263062 336134
rect 263146 335898 263382 336134
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 267326 340718 267562 340954
rect 267646 340718 267882 340954
rect 267326 340398 267562 340634
rect 267646 340398 267882 340634
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 262826 228218 263062 228454
rect 263146 228218 263382 228454
rect 262826 227898 263062 228134
rect 263146 227898 263382 228134
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 267326 232718 267562 232954
rect 267646 232718 267882 232954
rect 267326 232398 267562 232634
rect 267646 232398 267882 232634
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 276326 529718 276562 529954
rect 276646 529718 276882 529954
rect 276326 529398 276562 529634
rect 276646 529398 276882 529634
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 276326 349718 276562 349954
rect 276646 349718 276882 349954
rect 276326 349398 276562 349634
rect 276646 349398 276882 349634
rect 276326 313718 276562 313954
rect 276646 313718 276882 313954
rect 276326 313398 276562 313634
rect 276646 313398 276882 313634
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 276326 241718 276562 241954
rect 276646 241718 276882 241954
rect 276326 241398 276562 241634
rect 276646 241398 276882 241634
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 280826 534218 281062 534454
rect 281146 534218 281382 534454
rect 280826 533898 281062 534134
rect 281146 533898 281382 534134
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 280826 354218 281062 354454
rect 281146 354218 281382 354454
rect 280826 353898 281062 354134
rect 281146 353898 281382 354134
rect 280826 318218 281062 318454
rect 281146 318218 281382 318454
rect 280826 317898 281062 318134
rect 281146 317898 281382 318134
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 280826 246218 281062 246454
rect 281146 246218 281382 246454
rect 280826 245898 281062 246134
rect 281146 245898 281382 246134
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 285326 322718 285562 322954
rect 285646 322718 285882 322954
rect 285326 322398 285562 322634
rect 285646 322398 285882 322634
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 298826 516218 299062 516454
rect 299146 516218 299382 516454
rect 298826 515898 299062 516134
rect 299146 515898 299382 516134
rect 298826 480218 299062 480454
rect 299146 480218 299382 480454
rect 298826 479898 299062 480134
rect 299146 479898 299382 480134
rect 298826 444218 299062 444454
rect 299146 444218 299382 444454
rect 298826 443898 299062 444134
rect 299146 443898 299382 444134
rect 298826 408218 299062 408454
rect 299146 408218 299382 408454
rect 298826 407898 299062 408134
rect 299146 407898 299382 408134
rect 298826 372218 299062 372454
rect 299146 372218 299382 372454
rect 298826 371898 299062 372134
rect 299146 371898 299382 372134
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 298826 228218 299062 228454
rect 299146 228218 299382 228454
rect 298826 227898 299062 228134
rect 299146 227898 299382 228134
rect 298826 192218 299062 192454
rect 299146 192218 299382 192454
rect 298826 191898 299062 192134
rect 299146 191898 299382 192134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 303326 556718 303562 556954
rect 303646 556718 303882 556954
rect 303326 556398 303562 556634
rect 303646 556398 303882 556634
rect 303326 520718 303562 520954
rect 303646 520718 303882 520954
rect 303326 520398 303562 520634
rect 303646 520398 303882 520634
rect 303326 484718 303562 484954
rect 303646 484718 303882 484954
rect 303326 484398 303562 484634
rect 303646 484398 303882 484634
rect 303326 448718 303562 448954
rect 303646 448718 303882 448954
rect 303326 448398 303562 448634
rect 303646 448398 303882 448634
rect 303326 412718 303562 412954
rect 303646 412718 303882 412954
rect 303326 412398 303562 412634
rect 303646 412398 303882 412634
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 303326 232718 303562 232954
rect 303646 232718 303882 232954
rect 303326 232398 303562 232634
rect 303646 232398 303882 232634
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 312326 529718 312562 529954
rect 312646 529718 312882 529954
rect 312326 529398 312562 529634
rect 312646 529398 312882 529634
rect 312326 493718 312562 493954
rect 312646 493718 312882 493954
rect 312326 493398 312562 493634
rect 312646 493398 312882 493634
rect 312326 457718 312562 457954
rect 312646 457718 312882 457954
rect 312326 457398 312562 457634
rect 312646 457398 312882 457634
rect 312326 421718 312562 421954
rect 312646 421718 312882 421954
rect 312326 421398 312562 421634
rect 312646 421398 312882 421634
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 312326 313718 312562 313954
rect 312646 313718 312882 313954
rect 312326 313398 312562 313634
rect 312646 313398 312882 313634
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 312326 241718 312562 241954
rect 312646 241718 312882 241954
rect 312326 241398 312562 241634
rect 312646 241398 312882 241634
rect 312326 205718 312562 205954
rect 312646 205718 312882 205954
rect 312326 205398 312562 205634
rect 312646 205398 312882 205634
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 316826 534218 317062 534454
rect 317146 534218 317382 534454
rect 316826 533898 317062 534134
rect 317146 533898 317382 534134
rect 316826 498218 317062 498454
rect 317146 498218 317382 498454
rect 316826 497898 317062 498134
rect 317146 497898 317382 498134
rect 316826 462218 317062 462454
rect 317146 462218 317382 462454
rect 316826 461898 317062 462134
rect 317146 461898 317382 462134
rect 316826 426218 317062 426454
rect 317146 426218 317382 426454
rect 316826 425898 317062 426134
rect 317146 425898 317382 426134
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 316826 318218 317062 318454
rect 317146 318218 317382 318454
rect 316826 317898 317062 318134
rect 317146 317898 317382 318134
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 316826 246218 317062 246454
rect 317146 246218 317382 246454
rect 316826 245898 317062 246134
rect 317146 245898 317382 246134
rect 316826 210218 317062 210454
rect 317146 210218 317382 210454
rect 316826 209898 317062 210134
rect 317146 209898 317382 210134
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 321326 538718 321562 538954
rect 321646 538718 321882 538954
rect 321326 538398 321562 538634
rect 321646 538398 321882 538634
rect 321326 502718 321562 502954
rect 321646 502718 321882 502954
rect 321326 502398 321562 502634
rect 321646 502398 321882 502634
rect 321326 466718 321562 466954
rect 321646 466718 321882 466954
rect 321326 466398 321562 466634
rect 321646 466398 321882 466634
rect 321326 430718 321562 430954
rect 321646 430718 321882 430954
rect 321326 430398 321562 430634
rect 321646 430398 321882 430634
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 321326 322718 321562 322954
rect 321646 322718 321882 322954
rect 321326 322398 321562 322634
rect 321646 322398 321882 322634
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 321326 214718 321562 214954
rect 321646 214718 321882 214954
rect 321326 214398 321562 214634
rect 321646 214398 321882 214634
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 321326 178718 321562 178954
rect 321646 178718 321882 178954
rect 321326 178398 321562 178634
rect 321646 178398 321882 178634
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 330326 511718 330562 511954
rect 330646 511718 330882 511954
rect 330326 511398 330562 511634
rect 330646 511398 330882 511634
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 330326 439718 330562 439954
rect 330646 439718 330882 439954
rect 330326 439398 330562 439634
rect 330646 439398 330882 439634
rect 330326 403718 330562 403954
rect 330646 403718 330882 403954
rect 330326 403398 330562 403634
rect 330646 403398 330882 403634
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 334826 516218 335062 516454
rect 335146 516218 335382 516454
rect 334826 515898 335062 516134
rect 335146 515898 335382 516134
rect 334826 480218 335062 480454
rect 335146 480218 335382 480454
rect 334826 479898 335062 480134
rect 335146 479898 335382 480134
rect 334826 444218 335062 444454
rect 335146 444218 335382 444454
rect 334826 443898 335062 444134
rect 335146 443898 335382 444134
rect 334826 408218 335062 408454
rect 335146 408218 335382 408454
rect 334826 407898 335062 408134
rect 335146 407898 335382 408134
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 314250 151718 314486 151954
rect 314250 151398 314486 151634
rect 317514 151718 317750 151954
rect 317514 151398 317750 151634
rect 312618 147218 312854 147454
rect 312618 146898 312854 147134
rect 315882 147218 316118 147454
rect 315882 146898 316118 147134
rect 319146 147218 319382 147454
rect 319146 146898 319382 147134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 314250 115718 314486 115954
rect 314250 115398 314486 115634
rect 317514 115718 317750 115954
rect 317514 115398 317750 115634
rect 312618 111218 312854 111454
rect 312618 110898 312854 111134
rect 315882 111218 316118 111454
rect 315882 110898 316118 111134
rect 319146 111218 319382 111454
rect 319146 110898 319382 111134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 330326 223718 330562 223954
rect 330646 223718 330882 223954
rect 330326 223398 330562 223634
rect 330646 223398 330882 223634
rect 330326 187718 330562 187954
rect 330646 187718 330882 187954
rect 330326 187398 330562 187634
rect 330646 187398 330882 187634
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 339326 556718 339562 556954
rect 339646 556718 339882 556954
rect 339326 556398 339562 556634
rect 339646 556398 339882 556634
rect 339326 520718 339562 520954
rect 339646 520718 339882 520954
rect 339326 520398 339562 520634
rect 339646 520398 339882 520634
rect 339326 484718 339562 484954
rect 339646 484718 339882 484954
rect 339326 484398 339562 484634
rect 339646 484398 339882 484634
rect 339326 448718 339562 448954
rect 339646 448718 339882 448954
rect 339326 448398 339562 448634
rect 339646 448398 339882 448634
rect 339326 412718 339562 412954
rect 339646 412718 339882 412954
rect 339326 412398 339562 412634
rect 339646 412398 339882 412634
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 334826 228218 335062 228454
rect 335146 228218 335382 228454
rect 334826 227898 335062 228134
rect 335146 227898 335382 228134
rect 334826 192218 335062 192454
rect 335146 192218 335382 192454
rect 334826 191898 335062 192134
rect 335146 191898 335382 192134
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 339326 232718 339562 232954
rect 339646 232718 339882 232954
rect 339326 232398 339562 232634
rect 339646 232398 339882 232634
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 348326 529718 348562 529954
rect 348646 529718 348882 529954
rect 348326 529398 348562 529634
rect 348646 529398 348882 529634
rect 348326 493718 348562 493954
rect 348646 493718 348882 493954
rect 348326 493398 348562 493634
rect 348646 493398 348882 493634
rect 348326 457718 348562 457954
rect 348646 457718 348882 457954
rect 348326 457398 348562 457634
rect 348646 457398 348882 457634
rect 348326 421718 348562 421954
rect 348646 421718 348882 421954
rect 348326 421398 348562 421634
rect 348646 421398 348882 421634
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 348326 313718 348562 313954
rect 348646 313718 348882 313954
rect 348326 313398 348562 313634
rect 348646 313398 348882 313634
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 348326 241718 348562 241954
rect 348646 241718 348882 241954
rect 348326 241398 348562 241634
rect 348646 241398 348882 241634
rect 348326 205718 348562 205954
rect 348646 205718 348882 205954
rect 348326 205398 348562 205634
rect 348646 205398 348882 205634
rect 348326 169718 348562 169954
rect 348646 169718 348882 169954
rect 348326 169398 348562 169634
rect 348646 169398 348882 169634
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 352826 426218 353062 426454
rect 353146 426218 353382 426454
rect 352826 425898 353062 426134
rect 353146 425898 353382 426134
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 357326 538718 357562 538954
rect 357646 538718 357882 538954
rect 357326 538398 357562 538634
rect 357646 538398 357882 538634
rect 357326 502718 357562 502954
rect 357646 502718 357882 502954
rect 357326 502398 357562 502634
rect 357646 502398 357882 502634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 384326 241718 384562 241954
rect 384646 241718 384882 241954
rect 384326 241398 384562 241634
rect 384646 241398 384882 241634
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 89610 259954
rect 89846 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 89610 259634
rect 89846 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 74250 255454
rect 74486 255218 104970 255454
rect 105206 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 74250 255134
rect 74486 254898 104970 255134
rect 105206 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 69128 151954
rect 69364 151718 164192 151954
rect 164428 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 227916 151954
rect 228152 151718 237847 151954
rect 238083 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 314250 151954
rect 314486 151718 317514 151954
rect 317750 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 69128 151634
rect 69364 151398 164192 151634
rect 164428 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 227916 151634
rect 228152 151398 237847 151634
rect 238083 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 314250 151634
rect 314486 151398 317514 151634
rect 317750 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 69808 147454
rect 70044 147218 163512 147454
rect 163748 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 222952 147454
rect 223188 147218 232882 147454
rect 233118 147218 242813 147454
rect 243049 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 312618 147454
rect 312854 147218 315882 147454
rect 316118 147218 319146 147454
rect 319382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 69808 147134
rect 70044 146898 163512 147134
rect 163748 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 222952 147134
rect 223188 146898 232882 147134
rect 233118 146898 242813 147134
rect 243049 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 312618 147134
rect 312854 146898 315882 147134
rect 316118 146898 319146 147134
rect 319382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 69128 115954
rect 69364 115718 164192 115954
rect 164428 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 227916 115954
rect 228152 115718 237847 115954
rect 238083 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 314250 115954
rect 314486 115718 317514 115954
rect 317750 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 69128 115634
rect 69364 115398 164192 115634
rect 164428 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 227916 115634
rect 228152 115398 237847 115634
rect 238083 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 314250 115634
rect 314486 115398 317514 115634
rect 317750 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 69808 111454
rect 70044 111218 163512 111454
rect 163748 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 222952 111454
rect 223188 111218 232882 111454
rect 233118 111218 242813 111454
rect 243049 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 312618 111454
rect 312854 111218 315882 111454
rect 316118 111218 319146 111454
rect 319382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 69808 111134
rect 70044 110898 163512 111134
rect 163748 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 222952 111134
rect 223188 110898 232882 111134
rect 233118 110898 242813 111134
rect 243049 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 312618 111134
rect 312854 110898 315882 111134
rect 316118 110898 319146 111134
rect 319382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use sky130_sram_1kbyte_1rw1r_32x256_8  openram_1kB
timestamp 0
transform 1 0 68800 0 1 95100
box 0 0 95956 79500
use wb_bridge_2way  wb_bridge_2way
timestamp 0
transform 1 0 310000 0 1 96000
box 0 144 12000 80000
use wb_openram_wrapper  wb_openram_wrapper
timestamp 0
transform 1 0 217000 0 1 96000
box 0 144 32000 79688
use wrapped_function_generator  wrapped_function_generator_0
timestamp 0
transform 1 0 70000 0 1 240000
box 0 0 50000 52000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 93100 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 176600 74414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 294000 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 93100 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 176600 110414 238000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 294000 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 93100 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 176600 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 94000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 178000 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 93100 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 176600 83414 238000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 294000 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 93100 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 176600 119414 238000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 294000 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 93100 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 176600 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 94000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 178000 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 93100 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 176600 92414 238000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 294000 92414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 93100 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 176600 128414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 93100 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 176600 164414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 94000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 178000 236414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 94000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 178000 308414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 -7654 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 -7654 101414 93100 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 294000 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 93100 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 176600 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 -7654 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 -7654 245414 94000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 178000 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 -7654 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 -7654 317414 94000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 178000 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 -7654 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 -7654 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 93100 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 294000 96914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 93100 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 176600 132914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 94000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 178000 240914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 94000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 178000 312914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 93100 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 176600 69914 238000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 294000 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 93100 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 176600 105914 238000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 294000 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 93100 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 176600 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 94000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 178000 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 94000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 178000 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 93100 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 176600 78914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 294000 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 93100 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 176600 114914 238000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 294000 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 93100 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 176600 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 94000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 178000 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 93100 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 176600 87914 238000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 294000 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 93100 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 176600 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 93100 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 176600 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 94000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 178000 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
