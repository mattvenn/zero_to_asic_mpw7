VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_etpu
  CLASS BLOCK ;
  FOREIGN wrapped_etpu ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 900.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.170 896.000 3.730 900.000 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 271.740 900.000 272.940 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.490 0.000 667.050 4.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.690 0.000 699.250 4.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.030 0.000 206.590 4.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 135.740 900.000 136.940 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 101.740 900.000 102.940 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.610 0.000 332.170 4.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.340 4.000 133.540 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 455.340 900.000 456.540 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 336.340 900.000 337.540 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.670 0.000 728.230 4.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.750 896.000 290.310 900.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 20.140 900.000 21.340 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 655.940 900.000 657.140 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.750 896.000 129.310 900.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.310 896.000 766.870 900.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.540 4.000 619.740 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.490 896.000 828.050 900.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.430 896.000 431.990 900.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.590 0.000 683.150 4.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.340 4.000 116.540 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.990 0.000 586.550 4.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.050 896.000 177.610 900.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.370 896.000 35.930 900.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.450 896.000 242.010 900.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 366.940 4.000 368.140 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 33.740 900.000 34.940 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.290 0.000 473.850 4.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 302.340 900.000 303.540 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 819.140 4.000 820.340 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 604.940 900.000 606.140 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.870 0.000 760.430 4.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.540 4.000 738.740 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.410 0.000 299.970 4.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.010 0.000 396.570 4.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.770 0.000 744.330 4.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.340 4.000 184.540 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.340 4.000 82.540 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.090 0.000 602.650 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.610 896.000 654.170 900.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.070 0.000 792.630 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.810 896.000 686.370 900.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 536.940 900.000 538.140 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 723.940 900.000 725.140 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 523.340 900.000 524.540 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 298.940 4.000 300.140 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.310 0.000 444.870 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.390 896.000 811.950 900.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.340 4.000 167.540 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 50.740 900.000 51.940 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.340 4.000 14.540 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.110 0.000 251.670 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 822.540 900.000 823.740 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.110 896.000 734.670 900.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.230 0.000 77.790 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.310 0.000 283.870 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 506.340 900.000 507.540 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.890 0.000 570.450 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.940 4.000 283.140 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.330 896.000 415.890 900.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.540 4.000 670.740 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.450 896.000 81.010 900.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.790 896.000 876.350 900.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.930 896.000 512.490 900.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 774.940 900.000 776.140 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 788.540 900.000 789.740 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 451.940 4.000 453.140 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.210 896.000 750.770 900.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 570.940 900.000 572.140 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.950 896.000 161.510 900.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 254.740 900.000 255.940 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 751.140 4.000 752.340 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.550 896.000 97.110 900.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 839.540 900.000 840.740 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 438.340 900.000 439.540 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 383.940 4.000 385.140 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 853.140 4.000 854.340 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.340 4.000 31.540 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.390 0.000 489.950 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 400.940 4.000 402.140 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.010 896.000 557.570 900.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.890 896.000 892.450 900.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.540 4.000 602.740 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.330 0.000 93.890 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.830 896.000 335.390 900.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 203.740 900.000 204.940 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.410 896.000 782.970 900.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.340 4.000 48.540 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 332.940 4.000 334.140 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.970 0.000 776.530 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.690 896.000 860.250 900.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.310 896.000 605.870 900.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 553.940 900.000 555.140 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.540 4.000 687.740 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.670 0.000 889.230 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 387.340 900.000 388.540 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.130 896.000 544.690 900.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.710 896.000 670.270 900.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 285.340 900.000 286.540 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.340 4.000 65.540 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.210 896.000 589.770 900.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.350 896.000 225.910 900.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.030 896.000 367.590 900.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.830 896.000 496.390 900.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.570 0.000 873.130 4.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.340 4.000 201.540 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 67.740 900.000 68.940 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.630 0.000 142.190 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.540 4.000 500.740 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.730 896.000 480.290 900.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 404.340 900.000 405.540 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 169.740 900.000 170.940 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 870.140 4.000 871.340 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 757.940 900.000 759.140 ;
    END
  END io_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 886.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 886.960 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.850 896.000 306.410 900.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 873.540 900.000 874.740 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.540 4.000 653.740 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 587.940 900.000 589.140 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 740.940 900.000 742.140 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.540 4.000 534.740 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.030 0.000 45.590 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.710 0.000 348.270 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 220.740 900.000 221.940 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.630 896.000 464.190 900.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.110 0.000 412.670 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 152.740 900.000 153.940 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.470 0.000 857.030 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 802.140 4.000 803.340 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.540 4.000 585.740 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 489.340 900.000 490.540 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.540 4.000 721.740 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 315.940 4.000 317.140 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.270 0.000 824.830 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.650 896.000 274.210 900.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.810 0.000 364.370 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 434.940 4.000 436.140 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.540 4.000 568.740 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 264.940 4.000 266.140 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.550 896.000 258.110 900.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.210 0.000 267.770 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.650 896.000 113.210 900.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 84.740 900.000 85.940 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.690 0.000 538.250 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 706.940 900.000 708.140 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.340 4.000 99.540 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.130 0.000 222.690 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.150 896.000 193.710 900.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.570 0.000 712.130 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.540 4.000 551.740 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.010 896.000 718.570 900.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.270 896.000 19.830 900.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.250 896.000 209.810 900.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.930 896.000 351.490 900.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.730 896.000 319.290 900.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.930 0.000 29.490 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.730 0.000 158.290 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.940 4.000 249.140 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.210 0.000 428.770 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 856.540 900.000 857.740 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.470 896.000 52.030 900.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.530 896.000 448.090 900.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.430 0.000 109.990 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 319.340 900.000 320.540 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 672.940 900.000 674.140 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 417.940 4.000 419.140 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 472.340 900.000 473.540 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 785.140 4.000 786.340 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.340 4.000 150.540 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 805.540 900.000 806.740 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.030 896.000 528.590 900.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.010 0.000 235.570 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 353.340 900.000 354.540 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.290 0.000 634.850 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 118.740 900.000 119.940 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 836.140 4.000 837.340 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.170 0.000 808.730 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.530 0.000 126.090 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.910 0.000 380.470 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 237.740 900.000 238.940 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 890.540 900.000 891.740 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.340 4.000 235.540 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.370 0.000 840.930 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.940 4.000 351.140 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 370.340 900.000 371.540 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.830 0.000 13.390 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 689.940 900.000 691.140 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.590 896.000 844.150 900.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 3.140 900.000 4.340 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.290 896.000 795.850 900.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 485.940 4.000 487.140 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.540 4.000 517.740 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.790 0.000 554.350 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -0.050 0.000 0.510 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.390 0.000 650.950 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.540 4.000 636.740 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.570 896.000 68.130 900.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.230 896.000 399.790 900.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 468.940 4.000 470.140 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.830 0.000 174.390 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.130 0.000 61.690 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.110 896.000 573.670 900.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.130 896.000 383.690 900.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.410 0.000 460.970 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.910 896.000 702.470 900.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 186.740 900.000 187.940 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.540 4.000 704.740 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 638.940 900.000 640.140 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.930 0.000 190.490 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.510 0.000 316.070 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.490 0.000 506.050 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 621.940 900.000 623.140 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.590 0.000 522.150 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.510 896.000 638.070 900.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.410 896.000 621.970 900.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 887.140 4.000 888.340 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.850 896.000 145.410 900.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.190 0.000 618.750 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.340 4.000 218.540 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 768.140 4.000 769.340 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 421.340 900.000 422.540 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 894.240 886.805 ;
      LAYER met1 ;
        RECT 0.070 6.500 894.240 886.960 ;
      LAYER met2 ;
        RECT 0.100 895.720 2.890 897.330 ;
        RECT 4.010 895.720 18.990 897.330 ;
        RECT 20.110 895.720 35.090 897.330 ;
        RECT 36.210 895.720 51.190 897.330 ;
        RECT 52.310 895.720 67.290 897.330 ;
        RECT 68.410 895.720 80.170 897.330 ;
        RECT 81.290 895.720 96.270 897.330 ;
        RECT 97.390 895.720 112.370 897.330 ;
        RECT 113.490 895.720 128.470 897.330 ;
        RECT 129.590 895.720 144.570 897.330 ;
        RECT 145.690 895.720 160.670 897.330 ;
        RECT 161.790 895.720 176.770 897.330 ;
        RECT 177.890 895.720 192.870 897.330 ;
        RECT 193.990 895.720 208.970 897.330 ;
        RECT 210.090 895.720 225.070 897.330 ;
        RECT 226.190 895.720 241.170 897.330 ;
        RECT 242.290 895.720 257.270 897.330 ;
        RECT 258.390 895.720 273.370 897.330 ;
        RECT 274.490 895.720 289.470 897.330 ;
        RECT 290.590 895.720 305.570 897.330 ;
        RECT 306.690 895.720 318.450 897.330 ;
        RECT 319.570 895.720 334.550 897.330 ;
        RECT 335.670 895.720 350.650 897.330 ;
        RECT 351.770 895.720 366.750 897.330 ;
        RECT 367.870 895.720 382.850 897.330 ;
        RECT 383.970 895.720 398.950 897.330 ;
        RECT 400.070 895.720 415.050 897.330 ;
        RECT 416.170 895.720 431.150 897.330 ;
        RECT 432.270 895.720 447.250 897.330 ;
        RECT 448.370 895.720 463.350 897.330 ;
        RECT 464.470 895.720 479.450 897.330 ;
        RECT 480.570 895.720 495.550 897.330 ;
        RECT 496.670 895.720 511.650 897.330 ;
        RECT 512.770 895.720 527.750 897.330 ;
        RECT 528.870 895.720 543.850 897.330 ;
        RECT 544.970 895.720 556.730 897.330 ;
        RECT 557.850 895.720 572.830 897.330 ;
        RECT 573.950 895.720 588.930 897.330 ;
        RECT 590.050 895.720 605.030 897.330 ;
        RECT 606.150 895.720 621.130 897.330 ;
        RECT 622.250 895.720 637.230 897.330 ;
        RECT 638.350 895.720 653.330 897.330 ;
        RECT 654.450 895.720 669.430 897.330 ;
        RECT 670.550 895.720 685.530 897.330 ;
        RECT 686.650 895.720 701.630 897.330 ;
        RECT 702.750 895.720 717.730 897.330 ;
        RECT 718.850 895.720 733.830 897.330 ;
        RECT 734.950 895.720 749.930 897.330 ;
        RECT 751.050 895.720 766.030 897.330 ;
        RECT 767.150 895.720 782.130 897.330 ;
        RECT 783.250 895.720 795.010 897.330 ;
        RECT 796.130 895.720 811.110 897.330 ;
        RECT 812.230 895.720 827.210 897.330 ;
        RECT 828.330 895.720 843.310 897.330 ;
        RECT 844.430 895.720 859.410 897.330 ;
        RECT 860.530 895.720 875.510 897.330 ;
        RECT 876.630 895.720 891.610 897.330 ;
        RECT 0.100 4.280 892.300 895.720 ;
        RECT 0.790 3.555 12.550 4.280 ;
        RECT 13.670 3.555 28.650 4.280 ;
        RECT 29.770 3.555 44.750 4.280 ;
        RECT 45.870 3.555 60.850 4.280 ;
        RECT 61.970 3.555 76.950 4.280 ;
        RECT 78.070 3.555 93.050 4.280 ;
        RECT 94.170 3.555 109.150 4.280 ;
        RECT 110.270 3.555 125.250 4.280 ;
        RECT 126.370 3.555 141.350 4.280 ;
        RECT 142.470 3.555 157.450 4.280 ;
        RECT 158.570 3.555 173.550 4.280 ;
        RECT 174.670 3.555 189.650 4.280 ;
        RECT 190.770 3.555 205.750 4.280 ;
        RECT 206.870 3.555 221.850 4.280 ;
        RECT 222.970 3.555 234.730 4.280 ;
        RECT 235.850 3.555 250.830 4.280 ;
        RECT 251.950 3.555 266.930 4.280 ;
        RECT 268.050 3.555 283.030 4.280 ;
        RECT 284.150 3.555 299.130 4.280 ;
        RECT 300.250 3.555 315.230 4.280 ;
        RECT 316.350 3.555 331.330 4.280 ;
        RECT 332.450 3.555 347.430 4.280 ;
        RECT 348.550 3.555 363.530 4.280 ;
        RECT 364.650 3.555 379.630 4.280 ;
        RECT 380.750 3.555 395.730 4.280 ;
        RECT 396.850 3.555 411.830 4.280 ;
        RECT 412.950 3.555 427.930 4.280 ;
        RECT 429.050 3.555 444.030 4.280 ;
        RECT 445.150 3.555 460.130 4.280 ;
        RECT 461.250 3.555 473.010 4.280 ;
        RECT 474.130 3.555 489.110 4.280 ;
        RECT 490.230 3.555 505.210 4.280 ;
        RECT 506.330 3.555 521.310 4.280 ;
        RECT 522.430 3.555 537.410 4.280 ;
        RECT 538.530 3.555 553.510 4.280 ;
        RECT 554.630 3.555 569.610 4.280 ;
        RECT 570.730 3.555 585.710 4.280 ;
        RECT 586.830 3.555 601.810 4.280 ;
        RECT 602.930 3.555 617.910 4.280 ;
        RECT 619.030 3.555 634.010 4.280 ;
        RECT 635.130 3.555 650.110 4.280 ;
        RECT 651.230 3.555 666.210 4.280 ;
        RECT 667.330 3.555 682.310 4.280 ;
        RECT 683.430 3.555 698.410 4.280 ;
        RECT 699.530 3.555 711.290 4.280 ;
        RECT 712.410 3.555 727.390 4.280 ;
        RECT 728.510 3.555 743.490 4.280 ;
        RECT 744.610 3.555 759.590 4.280 ;
        RECT 760.710 3.555 775.690 4.280 ;
        RECT 776.810 3.555 791.790 4.280 ;
        RECT 792.910 3.555 807.890 4.280 ;
        RECT 809.010 3.555 823.990 4.280 ;
        RECT 825.110 3.555 840.090 4.280 ;
        RECT 841.210 3.555 856.190 4.280 ;
        RECT 857.310 3.555 872.290 4.280 ;
        RECT 873.410 3.555 888.390 4.280 ;
        RECT 889.510 3.555 892.300 4.280 ;
      LAYER met3 ;
        RECT 4.000 890.140 895.600 891.305 ;
        RECT 4.000 888.740 896.000 890.140 ;
        RECT 4.400 886.740 896.000 888.740 ;
        RECT 4.000 875.140 896.000 886.740 ;
        RECT 4.000 873.140 895.600 875.140 ;
        RECT 4.000 871.740 896.000 873.140 ;
        RECT 4.400 869.740 896.000 871.740 ;
        RECT 4.000 858.140 896.000 869.740 ;
        RECT 4.000 856.140 895.600 858.140 ;
        RECT 4.000 854.740 896.000 856.140 ;
        RECT 4.400 852.740 896.000 854.740 ;
        RECT 4.000 841.140 896.000 852.740 ;
        RECT 4.000 839.140 895.600 841.140 ;
        RECT 4.000 837.740 896.000 839.140 ;
        RECT 4.400 835.740 896.000 837.740 ;
        RECT 4.000 824.140 896.000 835.740 ;
        RECT 4.000 822.140 895.600 824.140 ;
        RECT 4.000 820.740 896.000 822.140 ;
        RECT 4.400 818.740 896.000 820.740 ;
        RECT 4.000 807.140 896.000 818.740 ;
        RECT 4.000 805.140 895.600 807.140 ;
        RECT 4.000 803.740 896.000 805.140 ;
        RECT 4.400 801.740 896.000 803.740 ;
        RECT 4.000 790.140 896.000 801.740 ;
        RECT 4.000 788.140 895.600 790.140 ;
        RECT 4.000 786.740 896.000 788.140 ;
        RECT 4.400 784.740 896.000 786.740 ;
        RECT 4.000 776.540 896.000 784.740 ;
        RECT 4.000 774.540 895.600 776.540 ;
        RECT 4.000 769.740 896.000 774.540 ;
        RECT 4.400 767.740 896.000 769.740 ;
        RECT 4.000 759.540 896.000 767.740 ;
        RECT 4.000 757.540 895.600 759.540 ;
        RECT 4.000 752.740 896.000 757.540 ;
        RECT 4.400 750.740 896.000 752.740 ;
        RECT 4.000 742.540 896.000 750.740 ;
        RECT 4.000 740.540 895.600 742.540 ;
        RECT 4.000 739.140 896.000 740.540 ;
        RECT 4.400 737.140 896.000 739.140 ;
        RECT 4.000 725.540 896.000 737.140 ;
        RECT 4.000 723.540 895.600 725.540 ;
        RECT 4.000 722.140 896.000 723.540 ;
        RECT 4.400 720.140 896.000 722.140 ;
        RECT 4.000 708.540 896.000 720.140 ;
        RECT 4.000 706.540 895.600 708.540 ;
        RECT 4.000 705.140 896.000 706.540 ;
        RECT 4.400 703.140 896.000 705.140 ;
        RECT 4.000 691.540 896.000 703.140 ;
        RECT 4.000 689.540 895.600 691.540 ;
        RECT 4.000 688.140 896.000 689.540 ;
        RECT 4.400 686.140 896.000 688.140 ;
        RECT 4.000 674.540 896.000 686.140 ;
        RECT 4.000 672.540 895.600 674.540 ;
        RECT 4.000 671.140 896.000 672.540 ;
        RECT 4.400 669.140 896.000 671.140 ;
        RECT 4.000 657.540 896.000 669.140 ;
        RECT 4.000 655.540 895.600 657.540 ;
        RECT 4.000 654.140 896.000 655.540 ;
        RECT 4.400 652.140 896.000 654.140 ;
        RECT 4.000 640.540 896.000 652.140 ;
        RECT 4.000 638.540 895.600 640.540 ;
        RECT 4.000 637.140 896.000 638.540 ;
        RECT 4.400 635.140 896.000 637.140 ;
        RECT 4.000 623.540 896.000 635.140 ;
        RECT 4.000 621.540 895.600 623.540 ;
        RECT 4.000 620.140 896.000 621.540 ;
        RECT 4.400 618.140 896.000 620.140 ;
        RECT 4.000 606.540 896.000 618.140 ;
        RECT 4.000 604.540 895.600 606.540 ;
        RECT 4.000 603.140 896.000 604.540 ;
        RECT 4.400 601.140 896.000 603.140 ;
        RECT 4.000 589.540 896.000 601.140 ;
        RECT 4.000 587.540 895.600 589.540 ;
        RECT 4.000 586.140 896.000 587.540 ;
        RECT 4.400 584.140 896.000 586.140 ;
        RECT 4.000 572.540 896.000 584.140 ;
        RECT 4.000 570.540 895.600 572.540 ;
        RECT 4.000 569.140 896.000 570.540 ;
        RECT 4.400 567.140 896.000 569.140 ;
        RECT 4.000 555.540 896.000 567.140 ;
        RECT 4.000 553.540 895.600 555.540 ;
        RECT 4.000 552.140 896.000 553.540 ;
        RECT 4.400 550.140 896.000 552.140 ;
        RECT 4.000 538.540 896.000 550.140 ;
        RECT 4.000 536.540 895.600 538.540 ;
        RECT 4.000 535.140 896.000 536.540 ;
        RECT 4.400 533.140 896.000 535.140 ;
        RECT 4.000 524.940 896.000 533.140 ;
        RECT 4.000 522.940 895.600 524.940 ;
        RECT 4.000 518.140 896.000 522.940 ;
        RECT 4.400 516.140 896.000 518.140 ;
        RECT 4.000 507.940 896.000 516.140 ;
        RECT 4.000 505.940 895.600 507.940 ;
        RECT 4.000 501.140 896.000 505.940 ;
        RECT 4.400 499.140 896.000 501.140 ;
        RECT 4.000 490.940 896.000 499.140 ;
        RECT 4.000 488.940 895.600 490.940 ;
        RECT 4.000 487.540 896.000 488.940 ;
        RECT 4.400 485.540 896.000 487.540 ;
        RECT 4.000 473.940 896.000 485.540 ;
        RECT 4.000 471.940 895.600 473.940 ;
        RECT 4.000 470.540 896.000 471.940 ;
        RECT 4.400 468.540 896.000 470.540 ;
        RECT 4.000 456.940 896.000 468.540 ;
        RECT 4.000 454.940 895.600 456.940 ;
        RECT 4.000 453.540 896.000 454.940 ;
        RECT 4.400 451.540 896.000 453.540 ;
        RECT 4.000 439.940 896.000 451.540 ;
        RECT 4.000 437.940 895.600 439.940 ;
        RECT 4.000 436.540 896.000 437.940 ;
        RECT 4.400 434.540 896.000 436.540 ;
        RECT 4.000 422.940 896.000 434.540 ;
        RECT 4.000 420.940 895.600 422.940 ;
        RECT 4.000 419.540 896.000 420.940 ;
        RECT 4.400 417.540 896.000 419.540 ;
        RECT 4.000 405.940 896.000 417.540 ;
        RECT 4.000 403.940 895.600 405.940 ;
        RECT 4.000 402.540 896.000 403.940 ;
        RECT 4.400 400.540 896.000 402.540 ;
        RECT 4.000 388.940 896.000 400.540 ;
        RECT 4.000 386.940 895.600 388.940 ;
        RECT 4.000 385.540 896.000 386.940 ;
        RECT 4.400 383.540 896.000 385.540 ;
        RECT 4.000 371.940 896.000 383.540 ;
        RECT 4.000 369.940 895.600 371.940 ;
        RECT 4.000 368.540 896.000 369.940 ;
        RECT 4.400 366.540 896.000 368.540 ;
        RECT 4.000 354.940 896.000 366.540 ;
        RECT 4.000 352.940 895.600 354.940 ;
        RECT 4.000 351.540 896.000 352.940 ;
        RECT 4.400 349.540 896.000 351.540 ;
        RECT 4.000 337.940 896.000 349.540 ;
        RECT 4.000 335.940 895.600 337.940 ;
        RECT 4.000 334.540 896.000 335.940 ;
        RECT 4.400 332.540 896.000 334.540 ;
        RECT 4.000 320.940 896.000 332.540 ;
        RECT 4.000 318.940 895.600 320.940 ;
        RECT 4.000 317.540 896.000 318.940 ;
        RECT 4.400 315.540 896.000 317.540 ;
        RECT 4.000 303.940 896.000 315.540 ;
        RECT 4.000 301.940 895.600 303.940 ;
        RECT 4.000 300.540 896.000 301.940 ;
        RECT 4.400 298.540 896.000 300.540 ;
        RECT 4.000 286.940 896.000 298.540 ;
        RECT 4.000 284.940 895.600 286.940 ;
        RECT 4.000 283.540 896.000 284.940 ;
        RECT 4.400 281.540 896.000 283.540 ;
        RECT 4.000 273.340 896.000 281.540 ;
        RECT 4.000 271.340 895.600 273.340 ;
        RECT 4.000 266.540 896.000 271.340 ;
        RECT 4.400 264.540 896.000 266.540 ;
        RECT 4.000 256.340 896.000 264.540 ;
        RECT 4.000 254.340 895.600 256.340 ;
        RECT 4.000 249.540 896.000 254.340 ;
        RECT 4.400 247.540 896.000 249.540 ;
        RECT 4.000 239.340 896.000 247.540 ;
        RECT 4.000 237.340 895.600 239.340 ;
        RECT 4.000 235.940 896.000 237.340 ;
        RECT 4.400 233.940 896.000 235.940 ;
        RECT 4.000 222.340 896.000 233.940 ;
        RECT 4.000 220.340 895.600 222.340 ;
        RECT 4.000 218.940 896.000 220.340 ;
        RECT 4.400 216.940 896.000 218.940 ;
        RECT 4.000 205.340 896.000 216.940 ;
        RECT 4.000 203.340 895.600 205.340 ;
        RECT 4.000 201.940 896.000 203.340 ;
        RECT 4.400 199.940 896.000 201.940 ;
        RECT 4.000 188.340 896.000 199.940 ;
        RECT 4.000 186.340 895.600 188.340 ;
        RECT 4.000 184.940 896.000 186.340 ;
        RECT 4.400 182.940 896.000 184.940 ;
        RECT 4.000 171.340 896.000 182.940 ;
        RECT 4.000 169.340 895.600 171.340 ;
        RECT 4.000 167.940 896.000 169.340 ;
        RECT 4.400 165.940 896.000 167.940 ;
        RECT 4.000 154.340 896.000 165.940 ;
        RECT 4.000 152.340 895.600 154.340 ;
        RECT 4.000 150.940 896.000 152.340 ;
        RECT 4.400 148.940 896.000 150.940 ;
        RECT 4.000 137.340 896.000 148.940 ;
        RECT 4.000 135.340 895.600 137.340 ;
        RECT 4.000 133.940 896.000 135.340 ;
        RECT 4.400 131.940 896.000 133.940 ;
        RECT 4.000 120.340 896.000 131.940 ;
        RECT 4.000 118.340 895.600 120.340 ;
        RECT 4.000 116.940 896.000 118.340 ;
        RECT 4.400 114.940 896.000 116.940 ;
        RECT 4.000 103.340 896.000 114.940 ;
        RECT 4.000 101.340 895.600 103.340 ;
        RECT 4.000 99.940 896.000 101.340 ;
        RECT 4.400 97.940 896.000 99.940 ;
        RECT 4.000 86.340 896.000 97.940 ;
        RECT 4.000 84.340 895.600 86.340 ;
        RECT 4.000 82.940 896.000 84.340 ;
        RECT 4.400 80.940 896.000 82.940 ;
        RECT 4.000 69.340 896.000 80.940 ;
        RECT 4.000 67.340 895.600 69.340 ;
        RECT 4.000 65.940 896.000 67.340 ;
        RECT 4.400 63.940 896.000 65.940 ;
        RECT 4.000 52.340 896.000 63.940 ;
        RECT 4.000 50.340 895.600 52.340 ;
        RECT 4.000 48.940 896.000 50.340 ;
        RECT 4.400 46.940 896.000 48.940 ;
        RECT 4.000 35.340 896.000 46.940 ;
        RECT 4.000 33.340 895.600 35.340 ;
        RECT 4.000 31.940 896.000 33.340 ;
        RECT 4.400 29.940 896.000 31.940 ;
        RECT 4.000 21.740 896.000 29.940 ;
        RECT 4.000 19.740 895.600 21.740 ;
        RECT 4.000 14.940 896.000 19.740 ;
        RECT 4.400 12.940 896.000 14.940 ;
        RECT 4.000 4.740 896.000 12.940 ;
        RECT 4.000 3.575 895.600 4.740 ;
      LAYER met4 ;
        RECT 254.215 11.735 327.840 752.585 ;
        RECT 330.240 11.735 404.640 752.585 ;
        RECT 407.040 11.735 481.440 752.585 ;
        RECT 483.840 11.735 558.240 752.585 ;
        RECT 560.640 11.735 635.040 752.585 ;
        RECT 637.440 11.735 711.840 752.585 ;
        RECT 714.240 11.735 766.985 752.585 ;
  END
END wrapped_etpu
END LIBRARY

